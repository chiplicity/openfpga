magic
tech EFS8A
magscale 1 2
timestamp 1604431093
<< locali >>
rect 9137 27999 9171 28169
rect 12081 21539 12115 21641
rect 3433 14807 3467 15113
rect 5273 9367 5307 9605
<< viali >>
rect 5457 36873 5491 36907
rect 5273 36669 5307 36703
rect 5917 36533 5951 36567
rect 5641 36329 5675 36363
rect 9873 36329 9907 36363
rect 5457 36193 5491 36227
rect 9689 36193 9723 36227
rect 1593 35785 1627 35819
rect 3157 35785 3191 35819
rect 4261 35785 4295 35819
rect 5825 35785 5859 35819
rect 8125 35785 8159 35819
rect 9597 35785 9631 35819
rect 7021 35717 7055 35751
rect 9873 35717 9907 35751
rect 5457 35649 5491 35683
rect 1409 35581 1443 35615
rect 2973 35581 3007 35615
rect 3525 35581 3559 35615
rect 4077 35581 4111 35615
rect 5641 35581 5675 35615
rect 6837 35581 6871 35615
rect 7941 35581 7975 35615
rect 9689 35581 9723 35615
rect 1869 35445 1903 35479
rect 4629 35445 4663 35479
rect 6285 35445 6319 35479
rect 7481 35445 7515 35479
rect 8585 35445 8619 35479
rect 10333 35445 10367 35479
rect 1593 35241 1627 35275
rect 2697 35241 2731 35275
rect 4721 35241 4755 35275
rect 5825 35241 5859 35275
rect 7573 35241 7607 35275
rect 12541 35241 12575 35275
rect 1409 35105 1443 35139
rect 2513 35105 2547 35139
rect 4537 35105 4571 35139
rect 5641 35105 5675 35139
rect 7389 35105 7423 35139
rect 8493 35105 8527 35139
rect 9945 35105 9979 35139
rect 9689 35037 9723 35071
rect 8677 34969 8711 35003
rect 7941 34901 7975 34935
rect 9505 34901 9539 34935
rect 11069 34901 11103 34935
rect 1593 34697 1627 34731
rect 12173 34697 12207 34731
rect 5733 34629 5767 34663
rect 13001 34561 13035 34595
rect 1409 34493 1443 34527
rect 2053 34493 2087 34527
rect 2513 34493 2547 34527
rect 3341 34493 3375 34527
rect 3433 34493 3467 34527
rect 7389 34493 7423 34527
rect 7656 34493 7690 34527
rect 9321 34493 9355 34527
rect 9873 34493 9907 34527
rect 12909 34493 12943 34527
rect 3678 34425 3712 34459
rect 6653 34425 6687 34459
rect 10140 34425 10174 34459
rect 4813 34357 4847 34391
rect 7205 34357 7239 34391
rect 8769 34357 8803 34391
rect 9781 34357 9815 34391
rect 11253 34357 11287 34391
rect 11897 34357 11931 34391
rect 12449 34357 12483 34391
rect 12817 34357 12851 34391
rect 1961 34153 1995 34187
rect 3065 34153 3099 34187
rect 5365 34153 5399 34187
rect 9505 34153 9539 34187
rect 9965 34153 9999 34187
rect 1685 34085 1719 34119
rect 10701 34085 10735 34119
rect 11713 34085 11747 34119
rect 12142 34085 12176 34119
rect 1777 34017 1811 34051
rect 2881 34017 2915 34051
rect 4077 34017 4111 34051
rect 5181 34017 5215 34051
rect 6552 34017 6586 34051
rect 10793 34017 10827 34051
rect 11345 34017 11379 34051
rect 6285 33949 6319 33983
rect 10977 33949 11011 33983
rect 11897 33949 11931 33983
rect 4261 33881 4295 33915
rect 3525 33813 3559 33847
rect 4721 33813 4755 33847
rect 7665 33813 7699 33847
rect 10333 33813 10367 33847
rect 13277 33813 13311 33847
rect 1593 33609 1627 33643
rect 9045 33609 9079 33643
rect 10701 33609 10735 33643
rect 13829 33541 13863 33575
rect 2329 33473 2363 33507
rect 10241 33473 10275 33507
rect 11345 33473 11379 33507
rect 12909 33473 12943 33507
rect 13093 33473 13127 33507
rect 13461 33473 13495 33507
rect 1409 33405 1443 33439
rect 1961 33405 1995 33439
rect 4261 33405 4295 33439
rect 6377 33405 6411 33439
rect 7573 33405 7607 33439
rect 7665 33405 7699 33439
rect 10517 33405 10551 33439
rect 11069 33405 11103 33439
rect 11897 33405 11931 33439
rect 4506 33337 4540 33371
rect 7932 33337 7966 33371
rect 9873 33337 9907 33371
rect 11161 33337 11195 33371
rect 12817 33337 12851 33371
rect 14197 33337 14231 33371
rect 2973 33269 3007 33303
rect 3709 33269 3743 33303
rect 4169 33269 4203 33303
rect 5641 33269 5675 33303
rect 7021 33269 7055 33303
rect 12449 33269 12483 33303
rect 1593 33065 1627 33099
rect 4261 33065 4295 33099
rect 5917 33065 5951 33099
rect 7113 33065 7147 33099
rect 7573 33065 7607 33099
rect 10793 33065 10827 33099
rect 11253 33065 11287 33099
rect 12357 33065 12391 33099
rect 12817 33065 12851 33099
rect 7481 32997 7515 33031
rect 1409 32929 1443 32963
rect 11161 32929 11195 32963
rect 12725 32929 12759 32963
rect 6009 32861 6043 32895
rect 6193 32861 6227 32895
rect 7665 32861 7699 32895
rect 9689 32861 9723 32895
rect 11437 32861 11471 32895
rect 12909 32861 12943 32895
rect 9137 32793 9171 32827
rect 5181 32725 5215 32759
rect 5549 32725 5583 32759
rect 7021 32725 7055 32759
rect 8217 32725 8251 32759
rect 9413 32725 9447 32759
rect 10425 32725 10459 32759
rect 11989 32725 12023 32759
rect 7205 32521 7239 32555
rect 8585 32521 8619 32555
rect 8861 32521 8895 32555
rect 10241 32521 10275 32555
rect 10793 32521 10827 32555
rect 12909 32521 12943 32555
rect 1685 32453 1719 32487
rect 5181 32453 5215 32487
rect 7481 32453 7515 32487
rect 4353 32385 4387 32419
rect 5733 32385 5767 32419
rect 8125 32385 8159 32419
rect 9505 32385 9539 32419
rect 9597 32385 9631 32419
rect 11253 32385 11287 32419
rect 11437 32385 11471 32419
rect 12265 32385 12299 32419
rect 12449 32385 12483 32419
rect 4721 32317 4755 32351
rect 5549 32317 5583 32351
rect 7941 32317 7975 32351
rect 9413 32317 9447 32351
rect 5089 32249 5123 32283
rect 6561 32249 6595 32283
rect 7849 32249 7883 32283
rect 5641 32181 5675 32215
rect 6193 32181 6227 32215
rect 9045 32181 9079 32215
rect 10701 32181 10735 32215
rect 11161 32181 11195 32215
rect 11897 32181 11931 32215
rect 6009 31977 6043 32011
rect 6469 31977 6503 32011
rect 6837 31977 6871 32011
rect 7389 31977 7423 32011
rect 10057 31977 10091 32011
rect 10149 31977 10183 32011
rect 10517 31977 10551 32011
rect 11529 31977 11563 32011
rect 12449 31977 12483 32011
rect 7205 31909 7239 31943
rect 4077 31841 4111 31875
rect 4344 31841 4378 31875
rect 7757 31841 7791 31875
rect 11253 31841 11287 31875
rect 7849 31773 7883 31807
rect 8033 31773 8067 31807
rect 10609 31773 10643 31807
rect 10793 31773 10827 31807
rect 3065 31637 3099 31671
rect 5457 31637 5491 31671
rect 9137 31637 9171 31671
rect 4077 31433 4111 31467
rect 8125 31433 8159 31467
rect 9137 31433 9171 31467
rect 10885 31433 10919 31467
rect 13737 31433 13771 31467
rect 7481 31365 7515 31399
rect 2881 31297 2915 31331
rect 3617 31297 3651 31331
rect 5089 31297 5123 31331
rect 9689 31297 9723 31331
rect 4445 31229 4479 31263
rect 4997 31229 5031 31263
rect 9505 31229 9539 31263
rect 13553 31229 13587 31263
rect 14013 31229 14047 31263
rect 2513 31161 2547 31195
rect 3341 31161 3375 31195
rect 4905 31161 4939 31195
rect 5549 31161 5583 31195
rect 2973 31093 3007 31127
rect 3433 31093 3467 31127
rect 4537 31093 4571 31127
rect 7757 31093 7791 31127
rect 9045 31093 9079 31127
rect 9597 31093 9631 31127
rect 10149 31093 10183 31127
rect 10609 31093 10643 31127
rect 2421 30889 2455 30923
rect 2789 30889 2823 30923
rect 5549 30889 5583 30923
rect 6745 30889 6779 30923
rect 7481 30889 7515 30923
rect 7941 30889 7975 30923
rect 8309 30889 8343 30923
rect 9689 30889 9723 30923
rect 12909 30889 12943 30923
rect 2881 30821 2915 30855
rect 9229 30821 9263 30855
rect 11774 30821 11808 30855
rect 4445 30753 4479 30787
rect 10057 30753 10091 30787
rect 10149 30753 10183 30787
rect 2973 30685 3007 30719
rect 3801 30685 3835 30719
rect 4537 30685 4571 30719
rect 4721 30685 4755 30719
rect 6837 30685 6871 30719
rect 6929 30685 6963 30719
rect 8401 30685 8435 30719
rect 8493 30685 8527 30719
rect 10241 30685 10275 30719
rect 11529 30685 11563 30719
rect 3525 30617 3559 30651
rect 4077 30617 4111 30651
rect 5089 30617 5123 30651
rect 5825 30549 5859 30583
rect 6377 30549 6411 30583
rect 2145 30345 2179 30379
rect 4169 30345 4203 30379
rect 6193 30345 6227 30379
rect 10977 30345 11011 30379
rect 11897 30345 11931 30379
rect 8033 30277 8067 30311
rect 3341 30209 3375 30243
rect 3433 30209 3467 30243
rect 5641 30209 5675 30243
rect 5825 30209 5859 30243
rect 7297 30209 7331 30243
rect 7481 30209 7515 30243
rect 8769 30209 8803 30243
rect 10241 30209 10275 30243
rect 3249 30141 3283 30175
rect 6653 30141 6687 30175
rect 5549 30073 5583 30107
rect 9505 30073 9539 30107
rect 10057 30073 10091 30107
rect 11529 30073 11563 30107
rect 2513 30005 2547 30039
rect 2881 30005 2915 30039
rect 4537 30005 4571 30039
rect 4997 30005 5031 30039
rect 5181 30005 5215 30039
rect 6837 30005 6871 30039
rect 7205 30005 7239 30039
rect 8309 30005 8343 30039
rect 9045 30005 9079 30039
rect 9597 30005 9631 30039
rect 9965 30005 9999 30039
rect 10701 30005 10735 30039
rect 1593 29801 1627 29835
rect 3249 29801 3283 29835
rect 4353 29801 4387 29835
rect 6929 29801 6963 29835
rect 7573 29801 7607 29835
rect 7205 29733 7239 29767
rect 1409 29665 1443 29699
rect 2973 29665 3007 29699
rect 5172 29665 5206 29699
rect 8125 29665 8159 29699
rect 10508 29665 10542 29699
rect 4905 29597 4939 29631
rect 8217 29597 8251 29631
rect 8401 29597 8435 29631
rect 10241 29597 10275 29631
rect 2513 29461 2547 29495
rect 6285 29461 6319 29495
rect 7757 29461 7791 29495
rect 8861 29461 8895 29495
rect 9873 29461 9907 29495
rect 11621 29461 11655 29495
rect 1593 29257 1627 29291
rect 1961 29257 1995 29291
rect 4997 29257 5031 29291
rect 8125 29257 8159 29291
rect 9689 29257 9723 29291
rect 2329 29189 2363 29223
rect 5089 29189 5123 29223
rect 6101 29189 6135 29223
rect 10793 29189 10827 29223
rect 11805 29189 11839 29223
rect 4077 29121 4111 29155
rect 5549 29121 5583 29155
rect 5641 29121 5675 29155
rect 11253 29121 11287 29155
rect 11437 29121 11471 29155
rect 1409 29053 1443 29087
rect 4629 29053 4663 29087
rect 8309 29053 8343 29087
rect 11161 29053 11195 29087
rect 5457 28985 5491 29019
rect 7757 28985 7791 29019
rect 8576 28985 8610 29019
rect 10241 28985 10275 29019
rect 10609 28985 10643 29019
rect 7481 28917 7515 28951
rect 3065 28713 3099 28747
rect 4537 28713 4571 28747
rect 7665 28713 7699 28747
rect 8677 28713 8711 28747
rect 9413 28713 9447 28747
rect 10885 28713 10919 28747
rect 6530 28645 6564 28679
rect 11244 28645 11278 28679
rect 4905 28577 4939 28611
rect 6285 28577 6319 28611
rect 8401 28577 8435 28611
rect 10977 28577 11011 28611
rect 4997 28509 5031 28543
rect 5089 28509 5123 28543
rect 5641 28441 5675 28475
rect 10333 28441 10367 28475
rect 5917 28373 5951 28407
rect 12357 28373 12391 28407
rect 2881 28169 2915 28203
rect 3065 28169 3099 28203
rect 4997 28169 5031 28203
rect 5273 28169 5307 28203
rect 6009 28169 6043 28203
rect 6377 28169 6411 28203
rect 9137 28169 9171 28203
rect 9229 28169 9263 28203
rect 9413 28169 9447 28203
rect 11069 28169 11103 28203
rect 11437 28169 11471 28203
rect 3617 28033 3651 28067
rect 8493 28033 8527 28067
rect 8861 28033 8895 28067
rect 9965 28033 9999 28067
rect 3433 27965 3467 27999
rect 7389 27965 7423 27999
rect 8217 27965 8251 27999
rect 9137 27965 9171 27999
rect 9873 27965 9907 27999
rect 2605 27897 2639 27931
rect 3525 27897 3559 27931
rect 4629 27897 4663 27931
rect 7757 27897 7791 27931
rect 9781 27897 9815 27931
rect 7849 27829 7883 27863
rect 8309 27829 8343 27863
rect 2421 27625 2455 27659
rect 5457 27625 5491 27659
rect 7573 27625 7607 27659
rect 8033 27625 8067 27659
rect 10885 27625 10919 27659
rect 2881 27557 2915 27591
rect 7941 27557 7975 27591
rect 9505 27557 9539 27591
rect 11805 27557 11839 27591
rect 12142 27557 12176 27591
rect 2789 27489 2823 27523
rect 4344 27489 4378 27523
rect 10057 27489 10091 27523
rect 11897 27489 11931 27523
rect 3065 27421 3099 27455
rect 4077 27421 4111 27455
rect 8125 27421 8159 27455
rect 10149 27421 10183 27455
rect 10333 27421 10367 27455
rect 9137 27353 9171 27387
rect 9689 27353 9723 27387
rect 6929 27285 6963 27319
rect 13277 27285 13311 27319
rect 1777 27081 1811 27115
rect 3985 27081 4019 27115
rect 4905 27081 4939 27115
rect 8217 27081 8251 27115
rect 10241 27081 10275 27115
rect 2145 27013 2179 27047
rect 2513 27013 2547 27047
rect 4629 27013 4663 27047
rect 6285 27013 6319 27047
rect 7941 27013 7975 27047
rect 13461 27013 13495 27047
rect 7297 26945 7331 26979
rect 7481 26945 7515 26979
rect 8769 26945 8803 26979
rect 9689 26945 9723 26979
rect 9873 26945 9907 26979
rect 11345 26945 11379 26979
rect 13001 26945 13035 26979
rect 2605 26877 2639 26911
rect 9597 26877 9631 26911
rect 12909 26877 12943 26911
rect 2872 26809 2906 26843
rect 6653 26809 6687 26843
rect 11253 26809 11287 26843
rect 12265 26809 12299 26843
rect 12817 26809 12851 26843
rect 6837 26741 6871 26775
rect 7205 26741 7239 26775
rect 9045 26741 9079 26775
rect 9229 26741 9263 26775
rect 10609 26741 10643 26775
rect 10793 26741 10827 26775
rect 11161 26741 11195 26775
rect 11805 26741 11839 26775
rect 12449 26741 12483 26775
rect 2697 26537 2731 26571
rect 2973 26537 3007 26571
rect 5825 26537 5859 26571
rect 6377 26537 6411 26571
rect 7941 26537 7975 26571
rect 9965 26537 9999 26571
rect 10885 26537 10919 26571
rect 12357 26537 12391 26571
rect 10517 26469 10551 26503
rect 11244 26469 11278 26503
rect 13001 26469 13035 26503
rect 5457 26401 5491 26435
rect 6285 26401 6319 26435
rect 6469 26333 6503 26367
rect 7021 26333 7055 26367
rect 7481 26333 7515 26367
rect 10977 26333 11011 26367
rect 5917 26265 5951 26299
rect 9321 26265 9355 26299
rect 4629 26197 4663 26231
rect 8677 26197 8711 26231
rect 1593 25993 1627 26027
rect 6193 25993 6227 26027
rect 6837 25993 6871 26027
rect 10057 25993 10091 26027
rect 11161 25993 11195 26027
rect 11529 25993 11563 26027
rect 8585 25925 8619 25959
rect 10149 25925 10183 25959
rect 5089 25857 5123 25891
rect 7389 25857 7423 25891
rect 8493 25857 8527 25891
rect 9229 25857 9263 25891
rect 10609 25857 10643 25891
rect 10701 25857 10735 25891
rect 1409 25789 1443 25823
rect 4905 25789 4939 25823
rect 7205 25789 7239 25823
rect 8953 25789 8987 25823
rect 10517 25789 10551 25823
rect 9045 25721 9079 25755
rect 9689 25721 9723 25755
rect 1961 25653 1995 25687
rect 4077 25653 4111 25687
rect 4353 25653 4387 25687
rect 4537 25653 4571 25687
rect 4997 25653 5031 25687
rect 5917 25653 5951 25687
rect 6653 25653 6687 25687
rect 7297 25653 7331 25687
rect 2329 25449 2363 25483
rect 6561 25449 6595 25483
rect 8677 25449 8711 25483
rect 10241 25449 10275 25483
rect 2697 25381 2731 25415
rect 5448 25381 5482 25415
rect 2789 25245 2823 25279
rect 2973 25245 3007 25279
rect 4169 25245 4203 25279
rect 4629 25245 4663 25279
rect 5181 25245 5215 25279
rect 2237 25109 2271 25143
rect 7941 25109 7975 25143
rect 4077 24905 4111 24939
rect 6101 24905 6135 24939
rect 4537 24769 4571 24803
rect 5089 24769 5123 24803
rect 5181 24769 5215 24803
rect 2053 24701 2087 24735
rect 2145 24701 2179 24735
rect 2412 24701 2446 24735
rect 4997 24701 5031 24735
rect 5733 24701 5767 24735
rect 7757 24701 7791 24735
rect 7849 24701 7883 24735
rect 8105 24701 8139 24735
rect 1685 24565 1719 24599
rect 3525 24565 3559 24599
rect 4629 24565 4663 24599
rect 9229 24565 9263 24599
rect 2421 24361 2455 24395
rect 2789 24361 2823 24395
rect 4077 24361 4111 24395
rect 4537 24361 4571 24395
rect 7297 24361 7331 24395
rect 7849 24361 7883 24395
rect 9689 24361 9723 24395
rect 10149 24361 10183 24395
rect 7757 24293 7791 24327
rect 4445 24225 4479 24259
rect 10057 24225 10091 24259
rect 11345 24225 11379 24259
rect 11612 24225 11646 24259
rect 4629 24157 4663 24191
rect 8033 24157 8067 24191
rect 10241 24157 10275 24191
rect 6929 24021 6963 24055
rect 7389 24021 7423 24055
rect 8401 24021 8435 24055
rect 9229 24021 9263 24055
rect 12725 24021 12759 24055
rect 4169 23817 4203 23851
rect 4537 23817 4571 23851
rect 4813 23817 4847 23851
rect 7849 23817 7883 23851
rect 8585 23817 8619 23851
rect 10517 23817 10551 23851
rect 11437 23817 11471 23851
rect 8217 23749 8251 23783
rect 11069 23749 11103 23783
rect 7297 23681 7331 23715
rect 7389 23681 7423 23715
rect 6285 23613 6319 23647
rect 7205 23613 7239 23647
rect 9137 23613 9171 23647
rect 9404 23613 9438 23647
rect 6653 23545 6687 23579
rect 5825 23477 5859 23511
rect 6837 23477 6871 23511
rect 9045 23477 9079 23511
rect 11897 23477 11931 23511
rect 1593 23273 1627 23307
rect 5641 23273 5675 23307
rect 6193 23273 6227 23307
rect 7849 23273 7883 23307
rect 8217 23273 8251 23307
rect 11069 23273 11103 23307
rect 12633 23273 12667 23307
rect 4445 23205 4479 23239
rect 1409 23137 1443 23171
rect 4537 23137 4571 23171
rect 6101 23137 6135 23171
rect 7757 23137 7791 23171
rect 9956 23137 9990 23171
rect 12541 23137 12575 23171
rect 4629 23069 4663 23103
rect 6285 23069 6319 23103
rect 7113 23069 7147 23103
rect 8309 23069 8343 23103
rect 8401 23069 8435 23103
rect 9229 23069 9263 23103
rect 9689 23069 9723 23103
rect 12725 23069 12759 23103
rect 2789 22933 2823 22967
rect 4077 22933 4111 22967
rect 5733 22933 5767 22967
rect 12173 22933 12207 22967
rect 13185 22933 13219 22967
rect 2513 22729 2547 22763
rect 2697 22729 2731 22763
rect 4169 22729 4203 22763
rect 5641 22729 5675 22763
rect 6285 22729 6319 22763
rect 8033 22729 8067 22763
rect 8585 22729 8619 22763
rect 9965 22729 9999 22763
rect 11253 22729 11287 22763
rect 11897 22729 11931 22763
rect 1685 22661 1719 22695
rect 7021 22661 7055 22695
rect 8493 22661 8527 22695
rect 3157 22593 3191 22627
rect 3341 22593 3375 22627
rect 7481 22593 7515 22627
rect 7665 22593 7699 22627
rect 9137 22593 9171 22627
rect 10701 22593 10735 22627
rect 13093 22593 13127 22627
rect 13829 22593 13863 22627
rect 4261 22525 4295 22559
rect 6653 22525 6687 22559
rect 7389 22525 7423 22559
rect 9045 22525 9079 22559
rect 13461 22525 13495 22559
rect 3065 22457 3099 22491
rect 3801 22457 3835 22491
rect 4506 22457 4540 22491
rect 9689 22457 9723 22491
rect 10517 22457 10551 22491
rect 12265 22457 12299 22491
rect 12909 22457 12943 22491
rect 2237 22389 2271 22423
rect 8953 22389 8987 22423
rect 10149 22389 10183 22423
rect 10609 22389 10643 22423
rect 12449 22389 12483 22423
rect 12817 22389 12851 22423
rect 2421 22185 2455 22219
rect 2789 22185 2823 22219
rect 6193 22185 6227 22219
rect 7113 22185 7147 22219
rect 10057 22185 10091 22219
rect 11621 22185 11655 22219
rect 12817 22185 12851 22219
rect 2881 22117 2915 22151
rect 10793 22117 10827 22151
rect 1409 22049 1443 22083
rect 4629 22049 4663 22083
rect 5080 22049 5114 22083
rect 7665 22049 7699 22083
rect 7757 22049 7791 22083
rect 8953 22049 8987 22083
rect 11161 22049 11195 22083
rect 11713 22049 11747 22083
rect 3065 21981 3099 22015
rect 4353 21981 4387 22015
rect 4813 21981 4847 22015
rect 7941 21981 7975 22015
rect 10149 21981 10183 22015
rect 10333 21981 10367 22015
rect 11897 21981 11931 22015
rect 1593 21913 1627 21947
rect 7297 21913 7331 21947
rect 9505 21913 9539 21947
rect 11253 21913 11287 21947
rect 3893 21845 3927 21879
rect 8677 21845 8711 21879
rect 9689 21845 9723 21879
rect 12541 21845 12575 21879
rect 2145 21641 2179 21675
rect 4077 21641 4111 21675
rect 5181 21641 5215 21675
rect 6193 21641 6227 21675
rect 12081 21641 12115 21675
rect 12173 21641 12207 21675
rect 2513 21573 2547 21607
rect 9045 21573 9079 21607
rect 10149 21573 10183 21607
rect 12449 21573 12483 21607
rect 5825 21505 5859 21539
rect 9781 21505 9815 21539
rect 10793 21505 10827 21539
rect 11345 21505 11379 21539
rect 12081 21505 12115 21539
rect 13001 21505 13035 21539
rect 2697 21437 2731 21471
rect 6561 21437 6595 21471
rect 6837 21437 6871 21471
rect 7104 21437 7138 21471
rect 10517 21437 10551 21471
rect 1777 21369 1811 21403
rect 2964 21369 2998 21403
rect 5089 21369 5123 21403
rect 9413 21369 9447 21403
rect 12909 21369 12943 21403
rect 4721 21301 4755 21335
rect 5549 21301 5583 21335
rect 5641 21301 5675 21335
rect 8217 21301 8251 21335
rect 10609 21301 10643 21335
rect 11805 21301 11839 21335
rect 12817 21301 12851 21335
rect 2697 21097 2731 21131
rect 3065 21097 3099 21131
rect 4905 21097 4939 21131
rect 6745 21097 6779 21131
rect 7389 21097 7423 21131
rect 8861 21097 8895 21131
rect 9413 21097 9447 21131
rect 10517 21097 10551 21131
rect 11069 21097 11103 21131
rect 11161 21097 11195 21131
rect 12541 21097 12575 21131
rect 12909 21097 12943 21131
rect 5273 21029 5307 21063
rect 11621 21029 11655 21063
rect 5632 20961 5666 20995
rect 7665 20961 7699 20995
rect 8217 20961 8251 20995
rect 10241 20961 10275 20995
rect 11529 20961 11563 20995
rect 1685 20893 1719 20927
rect 5365 20893 5399 20927
rect 8309 20893 8343 20927
rect 8401 20893 8435 20927
rect 11805 20893 11839 20927
rect 7849 20757 7883 20791
rect 13185 20757 13219 20791
rect 5733 20553 5767 20587
rect 7297 20553 7331 20587
rect 8217 20553 8251 20587
rect 10425 20553 10459 20587
rect 11897 20553 11931 20587
rect 12449 20553 12483 20587
rect 11253 20485 11287 20519
rect 7389 20417 7423 20451
rect 13001 20417 13035 20451
rect 9045 20349 9079 20383
rect 12817 20349 12851 20383
rect 9312 20281 9346 20315
rect 12909 20281 12943 20315
rect 13461 20281 13495 20315
rect 5365 20213 5399 20247
rect 7849 20213 7883 20247
rect 8861 20213 8895 20247
rect 11529 20213 11563 20247
rect 7849 20009 7883 20043
rect 10057 20009 10091 20043
rect 10517 20009 10551 20043
rect 13001 20009 13035 20043
rect 11888 19941 11922 19975
rect 10425 19873 10459 19907
rect 11621 19873 11655 19907
rect 10701 19805 10735 19839
rect 9965 19737 9999 19771
rect 6929 19669 6963 19703
rect 8493 19669 8527 19703
rect 9137 19669 9171 19703
rect 11897 19465 11931 19499
rect 6653 19397 6687 19431
rect 7481 19329 7515 19363
rect 8953 19329 8987 19363
rect 11161 19329 11195 19363
rect 8309 19261 8343 19295
rect 10977 19261 11011 19295
rect 6285 19193 6319 19227
rect 7941 19193 7975 19227
rect 10149 19193 10183 19227
rect 10885 19193 10919 19227
rect 11529 19193 11563 19227
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 7297 19125 7331 19159
rect 8401 19125 8435 19159
rect 8769 19125 8803 19159
rect 8861 19125 8895 19159
rect 9781 19125 9815 19159
rect 10517 19125 10551 19159
rect 10057 18921 10091 18955
rect 10701 18921 10735 18955
rect 11161 18921 11195 18955
rect 11713 18921 11747 18955
rect 5181 18785 5215 18819
rect 5448 18785 5482 18819
rect 8217 18785 8251 18819
rect 8309 18717 8343 18751
rect 8401 18717 8435 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 6561 18581 6595 18615
rect 7849 18581 7883 18615
rect 9689 18581 9723 18615
rect 1593 18377 1627 18411
rect 7297 18377 7331 18411
rect 9505 18377 9539 18411
rect 10425 18377 10459 18411
rect 7665 18309 7699 18343
rect 1961 18241 1995 18275
rect 5641 18241 5675 18275
rect 1409 18173 1443 18207
rect 3617 18173 3651 18207
rect 8125 18173 8159 18207
rect 3884 18105 3918 18139
rect 5917 18105 5951 18139
rect 8392 18105 8426 18139
rect 3525 18037 3559 18071
rect 4997 18037 5031 18071
rect 8033 18037 8067 18071
rect 10057 18037 10091 18071
rect 10885 18037 10919 18071
rect 7389 17833 7423 17867
rect 10149 17833 10183 17867
rect 6254 17765 6288 17799
rect 12050 17765 12084 17799
rect 4353 17697 4387 17731
rect 4813 17697 4847 17731
rect 4905 17697 4939 17731
rect 10057 17697 10091 17731
rect 4997 17629 5031 17663
rect 6009 17629 6043 17663
rect 8493 17629 8527 17663
rect 10333 17629 10367 17663
rect 11805 17629 11839 17663
rect 3709 17561 3743 17595
rect 9689 17561 9723 17595
rect 4445 17493 4479 17527
rect 8125 17493 8159 17527
rect 9321 17493 9355 17527
rect 13185 17493 13219 17527
rect 6837 17289 6871 17323
rect 10609 17289 10643 17323
rect 11161 17289 11195 17323
rect 12173 17289 12207 17323
rect 5733 17221 5767 17255
rect 6101 17153 6135 17187
rect 7389 17153 7423 17187
rect 3525 17085 3559 17119
rect 3617 17085 3651 17119
rect 7849 17085 7883 17119
rect 9229 17085 9263 17119
rect 9496 17085 9530 17119
rect 3884 17017 3918 17051
rect 7297 17017 7331 17051
rect 9045 17017 9079 17051
rect 4997 16949 5031 16983
rect 6561 16949 6595 16983
rect 7205 16949 7239 16983
rect 11805 16949 11839 16983
rect 4905 16745 4939 16779
rect 5273 16745 5307 16779
rect 6469 16745 6503 16779
rect 7205 16745 7239 16779
rect 7665 16745 7699 16779
rect 9965 16745 9999 16779
rect 11897 16745 11931 16779
rect 5733 16677 5767 16711
rect 8861 16677 8895 16711
rect 5641 16609 5675 16643
rect 7573 16609 7607 16643
rect 9321 16609 9355 16643
rect 10517 16609 10551 16643
rect 10784 16609 10818 16643
rect 5825 16541 5859 16575
rect 7757 16541 7791 16575
rect 3709 16405 3743 16439
rect 4537 16405 4571 16439
rect 6837 16405 6871 16439
rect 10425 16405 10459 16439
rect 1593 16201 1627 16235
rect 7205 16201 7239 16235
rect 8309 16201 8343 16235
rect 8769 16201 8803 16235
rect 2329 16133 2363 16167
rect 3525 16133 3559 16167
rect 10333 16133 10367 16167
rect 1961 16065 1995 16099
rect 3433 16065 3467 16099
rect 4077 16065 4111 16099
rect 5549 16065 5583 16099
rect 7113 16065 7147 16099
rect 7757 16065 7791 16099
rect 9229 16065 9263 16099
rect 9321 16065 9355 16099
rect 10241 16065 10275 16099
rect 10885 16065 10919 16099
rect 1409 15997 1443 16031
rect 2421 15997 2455 16031
rect 3065 15997 3099 16031
rect 3893 15997 3927 16031
rect 8677 15997 8711 16031
rect 9137 15997 9171 16031
rect 6009 15929 6043 15963
rect 7573 15929 7607 15963
rect 9873 15929 9907 15963
rect 10701 15929 10735 15963
rect 2605 15861 2639 15895
rect 3985 15861 4019 15895
rect 4905 15861 4939 15895
rect 5273 15861 5307 15895
rect 6653 15861 6687 15895
rect 7665 15861 7699 15895
rect 10793 15861 10827 15895
rect 11437 15861 11471 15895
rect 3617 15657 3651 15691
rect 4077 15657 4111 15691
rect 6653 15657 6687 15691
rect 7113 15657 7147 15691
rect 7665 15657 7699 15691
rect 8861 15657 8895 15691
rect 10609 15657 10643 15691
rect 11805 15589 11839 15623
rect 12265 15589 12299 15623
rect 4445 15521 4479 15555
rect 7573 15521 7607 15555
rect 4537 15453 4571 15487
rect 4629 15453 4663 15487
rect 7757 15453 7791 15487
rect 9689 15453 9723 15487
rect 12357 15453 12391 15487
rect 12541 15453 12575 15487
rect 5181 15317 5215 15351
rect 7205 15317 7239 15351
rect 10977 15317 11011 15351
rect 11897 15317 11931 15351
rect 13001 15317 13035 15351
rect 3433 15113 3467 15147
rect 3617 15113 3651 15147
rect 7849 15113 7883 15147
rect 10793 15113 10827 15147
rect 12173 15113 12207 15147
rect 13461 15113 13495 15147
rect 3249 14841 3283 14875
rect 3985 15045 4019 15079
rect 6285 15045 6319 15079
rect 11805 15045 11839 15079
rect 5365 14977 5399 15011
rect 5917 14977 5951 15011
rect 7389 14977 7423 15011
rect 8585 14977 8619 15011
rect 9597 14977 9631 15011
rect 10701 14977 10735 15011
rect 11437 14977 11471 15011
rect 13001 14977 13035 15011
rect 4353 14909 4387 14943
rect 7297 14909 7331 14943
rect 8953 14909 8987 14943
rect 9505 14909 9539 14943
rect 11161 14909 11195 14943
rect 4629 14841 4663 14875
rect 5273 14841 5307 14875
rect 6653 14841 6687 14875
rect 9413 14841 9447 14875
rect 12817 14841 12851 14875
rect 3433 14773 3467 14807
rect 4813 14773 4847 14807
rect 5181 14773 5215 14807
rect 6837 14773 6871 14807
rect 7205 14773 7239 14807
rect 9045 14773 9079 14807
rect 10333 14773 10367 14807
rect 11253 14773 11287 14807
rect 12449 14773 12483 14807
rect 12909 14773 12943 14807
rect 4261 14569 4295 14603
rect 4721 14569 4755 14603
rect 6561 14569 6595 14603
rect 7297 14569 7331 14603
rect 7665 14569 7699 14603
rect 8033 14569 8067 14603
rect 9137 14569 9171 14603
rect 10241 14569 10275 14603
rect 11253 14569 11287 14603
rect 13185 14569 13219 14603
rect 6653 14501 6687 14535
rect 12072 14501 12106 14535
rect 4629 14433 4663 14467
rect 8401 14433 8435 14467
rect 10609 14433 10643 14467
rect 4813 14365 4847 14399
rect 6745 14365 6779 14399
rect 8493 14365 8527 14399
rect 8677 14365 8711 14399
rect 10149 14365 10183 14399
rect 10701 14365 10735 14399
rect 10885 14365 10919 14399
rect 11805 14365 11839 14399
rect 3065 14229 3099 14263
rect 6193 14229 6227 14263
rect 11713 14229 11747 14263
rect 5917 14025 5951 14059
rect 9229 14025 9263 14059
rect 10425 14025 10459 14059
rect 11529 14025 11563 14059
rect 12173 14025 12207 14059
rect 4353 13957 4387 13991
rect 6653 13957 6687 13991
rect 10333 13957 10367 13991
rect 7389 13889 7423 13923
rect 9965 13889 9999 13923
rect 11069 13889 11103 13923
rect 2881 13821 2915 13855
rect 2973 13821 3007 13855
rect 4997 13821 5031 13855
rect 5365 13821 5399 13855
rect 6285 13821 6319 13855
rect 7849 13821 7883 13855
rect 8116 13821 8150 13855
rect 10793 13821 10827 13855
rect 11805 13821 11839 13855
rect 3240 13753 3274 13787
rect 7757 13753 7791 13787
rect 12449 13753 12483 13787
rect 10885 13685 10919 13719
rect 1593 13481 1627 13515
rect 2421 13481 2455 13515
rect 4721 13481 4755 13515
rect 7941 13481 7975 13515
rect 8033 13481 8067 13515
rect 9045 13481 9079 13515
rect 9413 13481 9447 13515
rect 10149 13481 10183 13515
rect 11161 13481 11195 13515
rect 12081 13481 12115 13515
rect 2881 13413 2915 13447
rect 5172 13413 5206 13447
rect 7573 13413 7607 13447
rect 1409 13345 1443 13379
rect 2789 13345 2823 13379
rect 8401 13345 8435 13379
rect 10517 13345 10551 13379
rect 2973 13277 3007 13311
rect 4261 13277 4295 13311
rect 4905 13277 4939 13311
rect 8493 13277 8527 13311
rect 8585 13277 8619 13311
rect 10609 13277 10643 13311
rect 10701 13277 10735 13311
rect 12173 13277 12207 13311
rect 12357 13277 12391 13311
rect 10057 13209 10091 13243
rect 11713 13209 11747 13243
rect 6285 13141 6319 13175
rect 6929 13141 6963 13175
rect 1777 12937 1811 12971
rect 4629 12937 4663 12971
rect 6285 12937 6319 12971
rect 8033 12937 8067 12971
rect 8493 12937 8527 12971
rect 10517 12937 10551 12971
rect 11805 12937 11839 12971
rect 12633 12937 12667 12971
rect 6837 12869 6871 12903
rect 4261 12801 4295 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 7389 12801 7423 12835
rect 12081 12801 12115 12835
rect 2145 12733 2179 12767
rect 2237 12733 2271 12767
rect 5549 12733 5583 12767
rect 7205 12733 7239 12767
rect 9045 12733 9079 12767
rect 9137 12733 9171 12767
rect 2504 12665 2538 12699
rect 4997 12665 5031 12699
rect 6561 12665 6595 12699
rect 7297 12665 7331 12699
rect 9382 12665 9416 12699
rect 3617 12597 3651 12631
rect 5181 12597 5215 12631
rect 11161 12597 11195 12631
rect 1685 12393 1719 12427
rect 2605 12393 2639 12427
rect 5549 12393 5583 12427
rect 6929 12393 6963 12427
rect 8493 12393 8527 12427
rect 9229 12393 9263 12427
rect 10241 12393 10275 12427
rect 11897 12393 11931 12427
rect 5273 12325 5307 12359
rect 5917 12325 5951 12359
rect 7380 12325 7414 12359
rect 4905 12257 4939 12291
rect 7113 12257 7147 12291
rect 10784 12257 10818 12291
rect 6009 12189 6043 12223
rect 6193 12189 6227 12223
rect 10517 12189 10551 12223
rect 2329 12121 2363 12155
rect 3065 12053 3099 12087
rect 3709 11849 3743 11883
rect 4813 11849 4847 11883
rect 5917 11849 5951 11883
rect 10517 11849 10551 11883
rect 10885 11849 10919 11883
rect 4353 11781 4387 11815
rect 2237 11713 2271 11747
rect 2329 11713 2363 11747
rect 5365 11713 5399 11747
rect 6653 11713 6687 11747
rect 6837 11713 6871 11747
rect 5181 11645 5215 11679
rect 5273 11645 5307 11679
rect 6285 11645 6319 11679
rect 7093 11645 7127 11679
rect 2574 11577 2608 11611
rect 4721 11577 4755 11611
rect 8217 11509 8251 11543
rect 4813 11305 4847 11339
rect 5273 11305 5307 11339
rect 5917 11305 5951 11339
rect 6377 11305 6411 11339
rect 7941 11305 7975 11339
rect 5181 11237 5215 11271
rect 6193 11237 6227 11271
rect 7481 11237 7515 11271
rect 6745 11169 6779 11203
rect 5365 11101 5399 11135
rect 6837 11101 6871 11135
rect 7021 11101 7055 11135
rect 1869 10965 1903 10999
rect 2329 10965 2363 10999
rect 3433 10965 3467 10999
rect 12541 10965 12575 10999
rect 3249 10761 3283 10795
rect 4905 10761 4939 10795
rect 5549 10761 5583 10795
rect 6101 10761 6135 10795
rect 3341 10693 3375 10727
rect 5181 10693 5215 10727
rect 1685 10625 1719 10659
rect 2329 10625 2363 10659
rect 3801 10625 3835 10659
rect 3893 10625 3927 10659
rect 13001 10625 13035 10659
rect 2145 10557 2179 10591
rect 2881 10489 2915 10523
rect 3709 10489 3743 10523
rect 6469 10489 6503 10523
rect 12265 10489 12299 10523
rect 12817 10489 12851 10523
rect 1777 10421 1811 10455
rect 2237 10421 2271 10455
rect 4445 10421 4479 10455
rect 7021 10421 7055 10455
rect 7757 10421 7791 10455
rect 12449 10421 12483 10455
rect 12909 10421 12943 10455
rect 1869 10217 1903 10251
rect 2421 10217 2455 10251
rect 4353 10217 4387 10251
rect 8125 10217 8159 10251
rect 12541 10217 12575 10251
rect 2789 10149 2823 10183
rect 4721 10081 4755 10115
rect 8033 10081 8067 10115
rect 10425 10081 10459 10115
rect 10692 10081 10726 10115
rect 13277 10081 13311 10115
rect 13369 10081 13403 10115
rect 2329 10013 2363 10047
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 4813 10013 4847 10047
rect 4905 10013 4939 10047
rect 8217 10013 8251 10047
rect 13461 10013 13495 10047
rect 12909 9945 12943 9979
rect 7389 9877 7423 9911
rect 7665 9877 7699 9911
rect 8953 9877 8987 9911
rect 11805 9877 11839 9911
rect 2881 9673 2915 9707
rect 10793 9673 10827 9707
rect 12449 9673 12483 9707
rect 1593 9605 1627 9639
rect 4445 9605 4479 9639
rect 5273 9605 5307 9639
rect 5825 9605 5859 9639
rect 11897 9605 11931 9639
rect 2053 9537 2087 9571
rect 3525 9537 3559 9571
rect 5089 9537 5123 9571
rect 1409 9469 1443 9503
rect 2421 9469 2455 9503
rect 3985 9469 4019 9503
rect 4353 9469 4387 9503
rect 4813 9469 4847 9503
rect 3341 9401 3375 9435
rect 4905 9401 4939 9435
rect 7941 9537 7975 9571
rect 12265 9537 12299 9571
rect 13001 9537 13035 9571
rect 14197 9537 14231 9571
rect 7665 9469 7699 9503
rect 8769 9469 8803 9503
rect 8861 9469 8895 9503
rect 11345 9469 11379 9503
rect 12817 9469 12851 9503
rect 13829 9469 13863 9503
rect 5457 9401 5491 9435
rect 7205 9401 7239 9435
rect 8401 9401 8435 9435
rect 9128 9401 9162 9435
rect 11161 9401 11195 9435
rect 2789 9333 2823 9367
rect 3249 9333 3283 9367
rect 5273 9333 5307 9367
rect 6193 9333 6227 9367
rect 6653 9333 6687 9367
rect 7297 9333 7331 9367
rect 7757 9333 7791 9367
rect 10241 9333 10275 9367
rect 12909 9333 12943 9367
rect 13461 9333 13495 9367
rect 2421 9129 2455 9163
rect 5457 9129 5491 9163
rect 7021 9129 7055 9163
rect 8033 9129 8067 9163
rect 10609 9129 10643 9163
rect 13093 9129 13127 9163
rect 13645 9129 13679 9163
rect 1961 9061 1995 9095
rect 7757 9061 7791 9095
rect 11980 9061 12014 9095
rect 2329 8993 2363 9027
rect 2789 8993 2823 9027
rect 4077 8993 4111 9027
rect 4344 8993 4378 9027
rect 8401 8993 8435 9027
rect 10517 8993 10551 9027
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 8493 8925 8527 8959
rect 8585 8925 8619 8959
rect 10701 8925 10735 8959
rect 11713 8925 11747 8959
rect 10149 8789 10183 8823
rect 1685 8585 1719 8619
rect 2053 8585 2087 8619
rect 2513 8585 2547 8619
rect 3341 8585 3375 8619
rect 6285 8585 6319 8619
rect 9045 8585 9079 8619
rect 10977 8585 11011 8619
rect 11713 8585 11747 8619
rect 12173 8585 12207 8619
rect 12449 8585 12483 8619
rect 9597 8517 9631 8551
rect 10701 8517 10735 8551
rect 11437 8517 11471 8551
rect 3985 8449 4019 8483
rect 4905 8449 4939 8483
rect 10149 8449 10183 8483
rect 12909 8449 12943 8483
rect 13001 8449 13035 8483
rect 2881 8381 2915 8415
rect 7113 8381 7147 8415
rect 9965 8381 9999 8415
rect 12817 8381 12851 8415
rect 3709 8313 3743 8347
rect 4721 8313 4755 8347
rect 6653 8313 6687 8347
rect 7380 8313 7414 8347
rect 9413 8313 9447 8347
rect 10057 8313 10091 8347
rect 3249 8245 3283 8279
rect 3801 8245 3835 8279
rect 4445 8245 4479 8279
rect 8493 8245 8527 8279
rect 2513 8041 2547 8075
rect 7113 8041 7147 8075
rect 8033 8041 8067 8075
rect 9045 8041 9079 8075
rect 10333 8041 10367 8075
rect 10425 8041 10459 8075
rect 12449 8041 12483 8075
rect 12909 8041 12943 8075
rect 7573 7973 7607 8007
rect 5448 7905 5482 7939
rect 7941 7905 7975 7939
rect 8401 7905 8435 7939
rect 10793 7905 10827 7939
rect 3433 7837 3467 7871
rect 5181 7837 5215 7871
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 9413 7837 9447 7871
rect 9873 7837 9907 7871
rect 10885 7837 10919 7871
rect 10977 7837 11011 7871
rect 6561 7701 6595 7735
rect 5089 7497 5123 7531
rect 8125 7497 8159 7531
rect 8401 7497 8435 7531
rect 9321 7497 9355 7531
rect 10793 7497 10827 7531
rect 6653 7429 6687 7463
rect 9413 7429 9447 7463
rect 11161 7429 11195 7463
rect 4353 7361 4387 7395
rect 5825 7361 5859 7395
rect 7481 7361 7515 7395
rect 7665 7361 7699 7395
rect 10057 7361 10091 7395
rect 1409 7293 1443 7327
rect 5549 7293 5583 7327
rect 5641 7293 5675 7327
rect 7389 7293 7423 7327
rect 8769 7293 8803 7327
rect 4721 7225 4755 7259
rect 6285 7225 6319 7259
rect 9781 7225 9815 7259
rect 1593 7157 1627 7191
rect 1961 7157 1995 7191
rect 5181 7157 5215 7191
rect 7021 7157 7055 7191
rect 9873 7157 9907 7191
rect 10425 7157 10459 7191
rect 5181 6953 5215 6987
rect 7021 6953 7055 6987
rect 1409 6817 1443 6851
rect 2421 6817 2455 6851
rect 4905 6817 4939 6851
rect 5641 6817 5675 6851
rect 5908 6817 5942 6851
rect 8125 6817 8159 6851
rect 9505 6817 9539 6851
rect 12081 6817 12115 6851
rect 12348 6817 12382 6851
rect 2605 6681 2639 6715
rect 9045 6681 9079 6715
rect 1593 6613 1627 6647
rect 1869 6613 1903 6647
rect 2329 6613 2363 6647
rect 7849 6613 7883 6647
rect 8309 6613 8343 6647
rect 8677 6613 8711 6647
rect 10057 6613 10091 6647
rect 13461 6613 13495 6647
rect 3065 6409 3099 6443
rect 6193 6409 6227 6443
rect 6653 6409 6687 6443
rect 7113 6409 7147 6443
rect 12081 6409 12115 6443
rect 12633 6409 12667 6443
rect 10057 6341 10091 6375
rect 4353 6273 4387 6307
rect 5365 6273 5399 6307
rect 8861 6273 8895 6307
rect 10609 6273 10643 6307
rect 1685 6205 1719 6239
rect 5273 6205 5307 6239
rect 7205 6205 7239 6239
rect 8769 6205 8803 6239
rect 9873 6205 9907 6239
rect 10425 6205 10459 6239
rect 1930 6137 1964 6171
rect 4721 6137 4755 6171
rect 7849 6137 7883 6171
rect 8677 6137 8711 6171
rect 10517 6137 10551 6171
rect 4813 6069 4847 6103
rect 5181 6069 5215 6103
rect 5825 6069 5859 6103
rect 7389 6069 7423 6103
rect 8125 6069 8159 6103
rect 8309 6069 8343 6103
rect 9597 6069 9631 6103
rect 1961 5865 1995 5899
rect 2421 5865 2455 5899
rect 7297 5865 7331 5899
rect 8217 5865 8251 5899
rect 9321 5865 9355 5899
rect 9873 5865 9907 5899
rect 10517 5865 10551 5899
rect 11069 5865 11103 5899
rect 1409 5729 1443 5763
rect 2881 5729 2915 5763
rect 3893 5729 3927 5763
rect 4445 5729 4479 5763
rect 5917 5729 5951 5763
rect 6184 5729 6218 5763
rect 8401 5729 8435 5763
rect 10425 5729 10459 5763
rect 11621 5729 11655 5763
rect 11888 5729 11922 5763
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 5457 5661 5491 5695
rect 10609 5661 10643 5695
rect 3433 5593 3467 5627
rect 1593 5525 1627 5559
rect 3065 5525 3099 5559
rect 4077 5525 4111 5559
rect 5825 5525 5859 5559
rect 8585 5525 8619 5559
rect 8953 5525 8987 5559
rect 10057 5525 10091 5559
rect 13001 5525 13035 5559
rect 2329 5321 2363 5355
rect 2789 5321 2823 5355
rect 4261 5321 4295 5355
rect 6193 5321 6227 5355
rect 7481 5321 7515 5355
rect 10149 5321 10183 5355
rect 11621 5321 11655 5355
rect 2053 5253 2087 5287
rect 2881 5185 2915 5219
rect 5549 5185 5583 5219
rect 7941 5185 7975 5219
rect 10425 5185 10459 5219
rect 11161 5185 11195 5219
rect 11989 5185 12023 5219
rect 1409 5117 1443 5151
rect 5641 5117 5675 5151
rect 6837 5117 6871 5151
rect 8125 5117 8159 5151
rect 10977 5117 11011 5151
rect 3126 5049 3160 5083
rect 6653 5049 6687 5083
rect 8370 5049 8404 5083
rect 11069 5049 11103 5083
rect 1593 4981 1627 5015
rect 4905 4981 4939 5015
rect 5825 4981 5859 5015
rect 7021 4981 7055 5015
rect 9505 4981 9539 5015
rect 10609 4981 10643 5015
rect 12633 4981 12667 5015
rect 2421 4777 2455 4811
rect 2789 4777 2823 4811
rect 4629 4777 4663 4811
rect 5089 4777 5123 4811
rect 6193 4777 6227 4811
rect 6653 4777 6687 4811
rect 7757 4777 7791 4811
rect 8125 4777 8159 4811
rect 8861 4777 8895 4811
rect 9505 4777 9539 4811
rect 10149 4777 10183 4811
rect 10885 4777 10919 4811
rect 11805 4777 11839 4811
rect 12449 4777 12483 4811
rect 2881 4709 2915 4743
rect 3525 4709 3559 4743
rect 3893 4709 3927 4743
rect 5733 4709 5767 4743
rect 8217 4709 8251 4743
rect 11437 4709 11471 4743
rect 4997 4641 5031 4675
rect 6561 4641 6595 4675
rect 7573 4641 7607 4675
rect 10793 4641 10827 4675
rect 12357 4641 12391 4675
rect 1409 4573 1443 4607
rect 1961 4573 1995 4607
rect 2973 4573 3007 4607
rect 5273 4573 5307 4607
rect 6745 4573 6779 4607
rect 8309 4573 8343 4607
rect 10977 4573 11011 4607
rect 12541 4573 12575 4607
rect 4537 4505 4571 4539
rect 6101 4505 6135 4539
rect 11989 4505 12023 4539
rect 2329 4437 2363 4471
rect 7297 4437 7331 4471
rect 10425 4437 10459 4471
rect 13001 4437 13035 4471
rect 4169 4233 4203 4267
rect 5089 4233 5123 4267
rect 5457 4233 5491 4267
rect 6653 4233 6687 4267
rect 6837 4233 6871 4267
rect 2605 4097 2639 4131
rect 2789 4097 2823 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 8125 4097 8159 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 9413 4097 9447 4131
rect 10701 4097 10735 4131
rect 10885 4097 10919 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 1593 4029 1627 4063
rect 2237 4029 2271 4063
rect 5641 4029 5675 4063
rect 8769 4029 8803 4063
rect 10149 4029 10183 4063
rect 11621 4029 11655 4063
rect 11989 4029 12023 4063
rect 12817 4029 12851 4063
rect 13461 4029 13495 4063
rect 3056 3961 3090 3995
rect 6193 3961 6227 3995
rect 1777 3893 1811 3927
rect 4813 3893 4847 3927
rect 5825 3893 5859 3927
rect 7205 3893 7239 3927
rect 8401 3893 8435 3927
rect 10241 3893 10275 3927
rect 10609 3893 10643 3927
rect 11345 3893 11379 3927
rect 12449 3893 12483 3927
rect 1685 3689 1719 3723
rect 2789 3689 2823 3723
rect 3525 3689 3559 3723
rect 3893 3689 3927 3723
rect 4721 3689 4755 3723
rect 4905 3689 4939 3723
rect 5273 3689 5307 3723
rect 6285 3689 6319 3723
rect 6837 3689 6871 3723
rect 7481 3689 7515 3723
rect 8033 3689 8067 3723
rect 8401 3689 8435 3723
rect 9505 3689 9539 3723
rect 12357 3689 12391 3723
rect 13001 3689 13035 3723
rect 5365 3621 5399 3655
rect 6929 3621 6963 3655
rect 11244 3621 11278 3655
rect 1777 3553 1811 3587
rect 2329 3553 2363 3587
rect 2881 3553 2915 3587
rect 8493 3553 8527 3587
rect 9689 3553 9723 3587
rect 10977 3553 11011 3587
rect 4261 3485 4295 3519
rect 5457 3485 5491 3519
rect 7021 3485 7055 3519
rect 8677 3485 8711 3519
rect 13461 3485 13495 3519
rect 1961 3417 1995 3451
rect 6469 3417 6503 3451
rect 13277 3417 13311 3451
rect 3065 3349 3099 3383
rect 5917 3349 5951 3383
rect 7849 3349 7883 3383
rect 9045 3349 9079 3383
rect 9873 3349 9907 3383
rect 10333 3349 10367 3383
rect 10885 3349 10919 3383
rect 1961 3145 1995 3179
rect 2973 3145 3007 3179
rect 3709 3145 3743 3179
rect 4169 3145 4203 3179
rect 5641 3145 5675 3179
rect 6193 3145 6227 3179
rect 7113 3145 7147 3179
rect 8217 3145 8251 3179
rect 10057 3145 10091 3179
rect 10701 3145 10735 3179
rect 11069 3145 11103 3179
rect 11805 3145 11839 3179
rect 12173 3145 12207 3179
rect 12449 3145 12483 3179
rect 6653 3077 6687 3111
rect 4261 3009 4295 3043
rect 7757 3009 7791 3043
rect 12909 3009 12943 3043
rect 13001 3009 13035 3043
rect 2053 2941 2087 2975
rect 3157 2941 3191 2975
rect 7481 2941 7515 2975
rect 8677 2941 8711 2975
rect 8944 2941 8978 2975
rect 11161 2941 11195 2975
rect 4528 2873 4562 2907
rect 7573 2873 7607 2907
rect 2237 2805 2271 2839
rect 3341 2805 3375 2839
rect 8585 2805 8619 2839
rect 11345 2805 11379 2839
rect 12817 2805 12851 2839
rect 13461 2805 13495 2839
rect 1961 2601 1995 2635
rect 3525 2601 3559 2635
rect 4997 2601 5031 2635
rect 5641 2601 5675 2635
rect 6745 2601 6779 2635
rect 8125 2601 8159 2635
rect 8493 2601 8527 2635
rect 11713 2601 11747 2635
rect 12633 2601 12667 2635
rect 13001 2601 13035 2635
rect 13645 2601 13679 2635
rect 5733 2533 5767 2567
rect 6377 2533 6411 2567
rect 9229 2533 9263 2567
rect 10048 2533 10082 2567
rect 13093 2533 13127 2567
rect 1777 2465 1811 2499
rect 2881 2465 2915 2499
rect 3893 2465 3927 2499
rect 4077 2465 4111 2499
rect 6929 2465 6963 2499
rect 7481 2465 7515 2499
rect 9597 2465 9631 2499
rect 9781 2465 9815 2499
rect 12449 2465 12483 2499
rect 5825 2397 5859 2431
rect 8585 2397 8619 2431
rect 8769 2397 8803 2431
rect 13277 2397 13311 2431
rect 14013 2397 14047 2431
rect 2789 2329 2823 2363
rect 4261 2329 4295 2363
rect 8033 2329 8067 2363
rect 2421 2261 2455 2295
rect 3065 2261 3099 2295
rect 5273 2261 5307 2295
rect 7113 2261 7147 2295
rect 11161 2261 11195 2295
rect 14381 2261 14415 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 5350 36864 5356 36916
rect 5408 36904 5414 36916
rect 5445 36907 5503 36913
rect 5445 36904 5457 36907
rect 5408 36876 5457 36904
rect 5408 36864 5414 36876
rect 5445 36873 5457 36876
rect 5491 36873 5503 36907
rect 5445 36867 5503 36873
rect 5261 36703 5319 36709
rect 5261 36669 5273 36703
rect 5307 36700 5319 36703
rect 5307 36672 5948 36700
rect 5307 36669 5319 36672
rect 5261 36663 5319 36669
rect 5920 36576 5948 36672
rect 5902 36564 5908 36576
rect 5863 36536 5908 36564
rect 5902 36524 5908 36536
rect 5960 36524 5966 36576
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 5629 36363 5687 36369
rect 5629 36329 5641 36363
rect 5675 36360 5687 36363
rect 6178 36360 6184 36372
rect 5675 36332 6184 36360
rect 5675 36329 5687 36332
rect 5629 36323 5687 36329
rect 6178 36320 6184 36332
rect 6236 36320 6242 36372
rect 9858 36360 9864 36372
rect 9819 36332 9864 36360
rect 9858 36320 9864 36332
rect 9916 36320 9922 36372
rect 5442 36224 5448 36236
rect 5403 36196 5448 36224
rect 5442 36184 5448 36196
rect 5500 36184 5506 36236
rect 9674 36224 9680 36236
rect 9635 36196 9680 36224
rect 9674 36184 9680 36196
rect 9732 36184 9738 36236
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 1578 35816 1584 35828
rect 1539 35788 1584 35816
rect 1578 35776 1584 35788
rect 1636 35776 1642 35828
rect 3145 35819 3203 35825
rect 3145 35785 3157 35819
rect 3191 35816 3203 35819
rect 3326 35816 3332 35828
rect 3191 35788 3332 35816
rect 3191 35785 3203 35788
rect 3145 35779 3203 35785
rect 3326 35776 3332 35788
rect 3384 35776 3390 35828
rect 3970 35776 3976 35828
rect 4028 35816 4034 35828
rect 4249 35819 4307 35825
rect 4249 35816 4261 35819
rect 4028 35788 4261 35816
rect 4028 35776 4034 35788
rect 4249 35785 4261 35788
rect 4295 35785 4307 35819
rect 4249 35779 4307 35785
rect 5813 35819 5871 35825
rect 5813 35785 5825 35819
rect 5859 35816 5871 35819
rect 6638 35816 6644 35828
rect 5859 35788 6644 35816
rect 5859 35785 5871 35788
rect 5813 35779 5871 35785
rect 6638 35776 6644 35788
rect 6696 35776 6702 35828
rect 7374 35776 7380 35828
rect 7432 35816 7438 35828
rect 8113 35819 8171 35825
rect 8113 35816 8125 35819
rect 7432 35788 8125 35816
rect 7432 35776 7438 35788
rect 8113 35785 8125 35788
rect 8159 35785 8171 35819
rect 9582 35816 9588 35828
rect 9543 35788 9588 35816
rect 8113 35779 8171 35785
rect 9582 35776 9588 35788
rect 9640 35776 9646 35828
rect 5718 35708 5724 35760
rect 5776 35748 5782 35760
rect 7009 35751 7067 35757
rect 7009 35748 7021 35751
rect 5776 35720 7021 35748
rect 5776 35708 5782 35720
rect 7009 35717 7021 35720
rect 7055 35717 7067 35751
rect 9858 35748 9864 35760
rect 9819 35720 9864 35748
rect 7009 35711 7067 35717
rect 9858 35708 9864 35720
rect 9916 35708 9922 35760
rect 4430 35640 4436 35692
rect 4488 35680 4494 35692
rect 5442 35680 5448 35692
rect 4488 35652 5448 35680
rect 4488 35640 4494 35652
rect 5442 35640 5448 35652
rect 5500 35640 5506 35692
rect 1397 35615 1455 35621
rect 1397 35581 1409 35615
rect 1443 35612 1455 35615
rect 1443 35584 1900 35612
rect 1443 35581 1455 35584
rect 1397 35575 1455 35581
rect 1872 35488 1900 35584
rect 2774 35572 2780 35624
rect 2832 35612 2838 35624
rect 2961 35615 3019 35621
rect 2961 35612 2973 35615
rect 2832 35584 2973 35612
rect 2832 35572 2838 35584
rect 2961 35581 2973 35584
rect 3007 35612 3019 35615
rect 3513 35615 3571 35621
rect 3513 35612 3525 35615
rect 3007 35584 3525 35612
rect 3007 35581 3019 35584
rect 2961 35575 3019 35581
rect 3513 35581 3525 35584
rect 3559 35581 3571 35615
rect 3513 35575 3571 35581
rect 4065 35615 4123 35621
rect 4065 35581 4077 35615
rect 4111 35612 4123 35615
rect 5629 35615 5687 35621
rect 4111 35584 4660 35612
rect 4111 35581 4123 35584
rect 4065 35575 4123 35581
rect 4632 35488 4660 35584
rect 5629 35581 5641 35615
rect 5675 35612 5687 35615
rect 6825 35615 6883 35621
rect 5675 35584 6316 35612
rect 5675 35581 5687 35584
rect 5629 35575 5687 35581
rect 1854 35476 1860 35488
rect 1815 35448 1860 35476
rect 1854 35436 1860 35448
rect 1912 35436 1918 35488
rect 4614 35476 4620 35488
rect 4575 35448 4620 35476
rect 4614 35436 4620 35448
rect 4672 35436 4678 35488
rect 6288 35485 6316 35584
rect 6825 35581 6837 35615
rect 6871 35612 6883 35615
rect 7929 35615 7987 35621
rect 6871 35584 7512 35612
rect 6871 35581 6883 35584
rect 6825 35575 6883 35581
rect 6273 35479 6331 35485
rect 6273 35445 6285 35479
rect 6319 35476 6331 35479
rect 6730 35476 6736 35488
rect 6319 35448 6736 35476
rect 6319 35445 6331 35448
rect 6273 35439 6331 35445
rect 6730 35436 6736 35448
rect 6788 35436 6794 35488
rect 7484 35485 7512 35584
rect 7929 35581 7941 35615
rect 7975 35612 7987 35615
rect 9677 35615 9735 35621
rect 7975 35584 8616 35612
rect 7975 35581 7987 35584
rect 7929 35575 7987 35581
rect 7469 35479 7527 35485
rect 7469 35445 7481 35479
rect 7515 35476 7527 35479
rect 8110 35476 8116 35488
rect 7515 35448 8116 35476
rect 7515 35445 7527 35448
rect 7469 35439 7527 35445
rect 8110 35436 8116 35448
rect 8168 35436 8174 35488
rect 8588 35485 8616 35584
rect 9677 35581 9689 35615
rect 9723 35612 9735 35615
rect 9723 35584 10364 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 8573 35479 8631 35485
rect 8573 35445 8585 35479
rect 8619 35476 8631 35479
rect 8662 35476 8668 35488
rect 8619 35448 8668 35476
rect 8619 35445 8631 35448
rect 8573 35439 8631 35445
rect 8662 35436 8668 35448
rect 8720 35436 8726 35488
rect 10336 35485 10364 35584
rect 10321 35479 10379 35485
rect 10321 35445 10333 35479
rect 10367 35476 10379 35479
rect 10410 35476 10416 35488
rect 10367 35448 10416 35476
rect 10367 35445 10379 35448
rect 10321 35439 10379 35445
rect 10410 35436 10416 35448
rect 10468 35436 10474 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 934 35232 940 35284
rect 992 35272 998 35284
rect 1581 35275 1639 35281
rect 1581 35272 1593 35275
rect 992 35244 1593 35272
rect 992 35232 998 35244
rect 1581 35241 1593 35244
rect 1627 35241 1639 35275
rect 1581 35235 1639 35241
rect 2130 35232 2136 35284
rect 2188 35272 2194 35284
rect 2685 35275 2743 35281
rect 2685 35272 2697 35275
rect 2188 35244 2697 35272
rect 2188 35232 2194 35244
rect 2685 35241 2697 35244
rect 2731 35241 2743 35275
rect 4706 35272 4712 35284
rect 4667 35244 4712 35272
rect 2685 35235 2743 35241
rect 4706 35232 4712 35244
rect 4764 35232 4770 35284
rect 4982 35232 4988 35284
rect 5040 35272 5046 35284
rect 5813 35275 5871 35281
rect 5813 35272 5825 35275
rect 5040 35244 5825 35272
rect 5040 35232 5046 35244
rect 5813 35241 5825 35244
rect 5859 35241 5871 35275
rect 7558 35272 7564 35284
rect 7519 35244 7564 35272
rect 5813 35235 5871 35241
rect 7558 35232 7564 35244
rect 7616 35232 7622 35284
rect 12526 35272 12532 35284
rect 12487 35244 12532 35272
rect 12526 35232 12532 35244
rect 12584 35232 12590 35284
rect 1397 35139 1455 35145
rect 1397 35105 1409 35139
rect 1443 35136 1455 35139
rect 1670 35136 1676 35148
rect 1443 35108 1676 35136
rect 1443 35105 1455 35108
rect 1397 35099 1455 35105
rect 1670 35096 1676 35108
rect 1728 35096 1734 35148
rect 2498 35136 2504 35148
rect 2459 35108 2504 35136
rect 2498 35096 2504 35108
rect 2556 35096 2562 35148
rect 4525 35139 4583 35145
rect 4525 35105 4537 35139
rect 4571 35136 4583 35139
rect 4706 35136 4712 35148
rect 4571 35108 4712 35136
rect 4571 35105 4583 35108
rect 4525 35099 4583 35105
rect 4706 35096 4712 35108
rect 4764 35096 4770 35148
rect 5626 35136 5632 35148
rect 5587 35108 5632 35136
rect 5626 35096 5632 35108
rect 5684 35096 5690 35148
rect 7190 35096 7196 35148
rect 7248 35136 7254 35148
rect 7377 35139 7435 35145
rect 7377 35136 7389 35139
rect 7248 35108 7389 35136
rect 7248 35096 7254 35108
rect 7377 35105 7389 35108
rect 7423 35105 7435 35139
rect 8478 35136 8484 35148
rect 8439 35108 8484 35136
rect 7377 35099 7435 35105
rect 8478 35096 8484 35108
rect 8536 35096 8542 35148
rect 9490 35096 9496 35148
rect 9548 35136 9554 35148
rect 9933 35139 9991 35145
rect 9933 35136 9945 35139
rect 9548 35108 9945 35136
rect 9548 35096 9554 35108
rect 9933 35105 9945 35108
rect 9979 35105 9991 35139
rect 9933 35099 9991 35105
rect 9674 35028 9680 35080
rect 9732 35068 9738 35080
rect 9732 35040 9777 35068
rect 9732 35028 9738 35040
rect 6914 34960 6920 35012
rect 6972 35000 6978 35012
rect 8665 35003 8723 35009
rect 8665 35000 8677 35003
rect 6972 34972 8677 35000
rect 6972 34960 6978 34972
rect 8665 34969 8677 34972
rect 8711 34969 8723 35003
rect 8665 34963 8723 34969
rect 7650 34892 7656 34944
rect 7708 34932 7714 34944
rect 7929 34935 7987 34941
rect 7929 34932 7941 34935
rect 7708 34904 7941 34932
rect 7708 34892 7714 34904
rect 7929 34901 7941 34904
rect 7975 34901 7987 34935
rect 7929 34895 7987 34901
rect 9493 34935 9551 34941
rect 9493 34901 9505 34935
rect 9539 34932 9551 34935
rect 11057 34935 11115 34941
rect 11057 34932 11069 34935
rect 9539 34904 11069 34932
rect 9539 34901 9551 34904
rect 9493 34895 9551 34901
rect 11057 34901 11069 34904
rect 11103 34932 11115 34935
rect 11146 34932 11152 34944
rect 11103 34904 11152 34932
rect 11103 34901 11115 34904
rect 11057 34895 11115 34901
rect 11146 34892 11152 34904
rect 11204 34892 11210 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 198 34688 204 34740
rect 256 34728 262 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 256 34700 1593 34728
rect 256 34688 262 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 1581 34691 1639 34697
rect 12066 34688 12072 34740
rect 12124 34728 12130 34740
rect 12161 34731 12219 34737
rect 12161 34728 12173 34731
rect 12124 34700 12173 34728
rect 12124 34688 12130 34700
rect 12161 34697 12173 34700
rect 12207 34697 12219 34731
rect 12161 34691 12219 34697
rect 5626 34620 5632 34672
rect 5684 34660 5690 34672
rect 5721 34663 5779 34669
rect 5721 34660 5733 34663
rect 5684 34632 5733 34660
rect 5684 34620 5690 34632
rect 5721 34629 5733 34632
rect 5767 34660 5779 34663
rect 7374 34660 7380 34672
rect 5767 34632 7380 34660
rect 5767 34629 5779 34632
rect 5721 34623 5779 34629
rect 7374 34620 7380 34632
rect 7432 34620 7438 34672
rect 12250 34552 12256 34604
rect 12308 34592 12314 34604
rect 12989 34595 13047 34601
rect 12989 34592 13001 34595
rect 12308 34564 13001 34592
rect 12308 34552 12314 34564
rect 12989 34561 13001 34564
rect 13035 34561 13047 34595
rect 12989 34555 13047 34561
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 2038 34524 2044 34536
rect 1443 34496 2044 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2130 34484 2136 34536
rect 2188 34524 2194 34536
rect 2498 34524 2504 34536
rect 2188 34496 2504 34524
rect 2188 34484 2194 34496
rect 2498 34484 2504 34496
rect 2556 34484 2562 34536
rect 3329 34527 3387 34533
rect 3329 34493 3341 34527
rect 3375 34524 3387 34527
rect 3421 34527 3479 34533
rect 3421 34524 3433 34527
rect 3375 34496 3433 34524
rect 3375 34493 3387 34496
rect 3329 34487 3387 34493
rect 3421 34493 3433 34496
rect 3467 34524 3479 34527
rect 4062 34524 4068 34536
rect 3467 34496 4068 34524
rect 3467 34493 3479 34496
rect 3421 34487 3479 34493
rect 4062 34484 4068 34496
rect 4120 34484 4126 34536
rect 7650 34533 7656 34536
rect 7377 34527 7435 34533
rect 7377 34493 7389 34527
rect 7423 34493 7435 34527
rect 7644 34524 7656 34533
rect 7611 34496 7656 34524
rect 7377 34487 7435 34493
rect 7644 34487 7656 34496
rect 7708 34524 7714 34536
rect 8202 34524 8208 34536
rect 7708 34496 8208 34524
rect 3510 34416 3516 34468
rect 3568 34456 3574 34468
rect 3666 34459 3724 34465
rect 3666 34456 3678 34459
rect 3568 34428 3678 34456
rect 3568 34416 3574 34428
rect 3666 34425 3678 34428
rect 3712 34425 3724 34459
rect 3666 34419 3724 34425
rect 6641 34459 6699 34465
rect 6641 34425 6653 34459
rect 6687 34456 6699 34459
rect 7392 34456 7420 34487
rect 7650 34484 7656 34487
rect 7708 34484 7714 34496
rect 8202 34484 8208 34496
rect 8260 34484 8266 34536
rect 8478 34484 8484 34536
rect 8536 34524 8542 34536
rect 9309 34527 9367 34533
rect 9309 34524 9321 34527
rect 8536 34496 9321 34524
rect 8536 34484 8542 34496
rect 9309 34493 9321 34496
rect 9355 34493 9367 34527
rect 9309 34487 9367 34493
rect 9674 34484 9680 34536
rect 9732 34524 9738 34536
rect 9861 34527 9919 34533
rect 9861 34524 9873 34527
rect 9732 34496 9873 34524
rect 9732 34484 9738 34496
rect 9861 34493 9873 34496
rect 9907 34493 9919 34527
rect 9861 34487 9919 34493
rect 7742 34456 7748 34468
rect 6687 34428 7748 34456
rect 6687 34425 6699 34428
rect 6641 34419 6699 34425
rect 7742 34416 7748 34428
rect 7800 34416 7806 34468
rect 4798 34388 4804 34400
rect 4759 34360 4804 34388
rect 4798 34348 4804 34360
rect 4856 34348 4862 34400
rect 7190 34388 7196 34400
rect 7151 34360 7196 34388
rect 7190 34348 7196 34360
rect 7248 34348 7254 34400
rect 8570 34348 8576 34400
rect 8628 34388 8634 34400
rect 8757 34391 8815 34397
rect 8757 34388 8769 34391
rect 8628 34360 8769 34388
rect 8628 34348 8634 34360
rect 8757 34357 8769 34360
rect 8803 34388 8815 34391
rect 9490 34388 9496 34400
rect 8803 34360 9496 34388
rect 8803 34357 8815 34360
rect 8757 34351 8815 34357
rect 9490 34348 9496 34360
rect 9548 34348 9554 34400
rect 9769 34391 9827 34397
rect 9769 34357 9781 34391
rect 9815 34388 9827 34391
rect 9876 34388 9904 34487
rect 12066 34484 12072 34536
rect 12124 34524 12130 34536
rect 12124 34496 12296 34524
rect 12124 34484 12130 34496
rect 10128 34459 10186 34465
rect 10128 34425 10140 34459
rect 10174 34456 10186 34459
rect 11146 34456 11152 34468
rect 10174 34428 11152 34456
rect 10174 34425 10186 34428
rect 10128 34419 10186 34425
rect 11146 34416 11152 34428
rect 11204 34416 11210 34468
rect 12268 34456 12296 34496
rect 12526 34484 12532 34536
rect 12584 34524 12590 34536
rect 12897 34527 12955 34533
rect 12897 34524 12909 34527
rect 12584 34496 12909 34524
rect 12584 34484 12590 34496
rect 12897 34493 12909 34496
rect 12943 34493 12955 34527
rect 12897 34487 12955 34493
rect 12268 34428 12848 34456
rect 12820 34400 12848 34428
rect 9950 34388 9956 34400
rect 9815 34360 9956 34388
rect 9815 34357 9827 34360
rect 9769 34351 9827 34357
rect 9950 34348 9956 34360
rect 10008 34348 10014 34400
rect 11241 34391 11299 34397
rect 11241 34357 11253 34391
rect 11287 34388 11299 34391
rect 11885 34391 11943 34397
rect 11885 34388 11897 34391
rect 11287 34360 11897 34388
rect 11287 34357 11299 34360
rect 11241 34351 11299 34357
rect 11885 34357 11897 34360
rect 11931 34388 11943 34391
rect 12066 34388 12072 34400
rect 11931 34360 12072 34388
rect 11931 34357 11943 34360
rect 11885 34351 11943 34357
rect 12066 34348 12072 34360
rect 12124 34388 12130 34400
rect 12250 34388 12256 34400
rect 12124 34360 12256 34388
rect 12124 34348 12130 34360
rect 12250 34348 12256 34360
rect 12308 34348 12314 34400
rect 12434 34348 12440 34400
rect 12492 34388 12498 34400
rect 12802 34388 12808 34400
rect 12492 34360 12537 34388
rect 12763 34360 12808 34388
rect 12492 34348 12498 34360
rect 12802 34348 12808 34360
rect 12860 34348 12866 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1394 34144 1400 34196
rect 1452 34184 1458 34196
rect 1949 34187 2007 34193
rect 1949 34184 1961 34187
rect 1452 34156 1961 34184
rect 1452 34144 1458 34156
rect 1949 34153 1961 34156
rect 1995 34153 2007 34187
rect 1949 34147 2007 34153
rect 2958 34144 2964 34196
rect 3016 34184 3022 34196
rect 3053 34187 3111 34193
rect 3053 34184 3065 34187
rect 3016 34156 3065 34184
rect 3016 34144 3022 34156
rect 3053 34153 3065 34156
rect 3099 34153 3111 34187
rect 3053 34147 3111 34153
rect 4154 34144 4160 34196
rect 4212 34184 4218 34196
rect 5353 34187 5411 34193
rect 5353 34184 5365 34187
rect 4212 34156 5365 34184
rect 4212 34144 4218 34156
rect 5353 34153 5365 34156
rect 5399 34153 5411 34187
rect 9490 34184 9496 34196
rect 9451 34156 9496 34184
rect 5353 34147 5411 34153
rect 9490 34144 9496 34156
rect 9548 34144 9554 34196
rect 9950 34184 9956 34196
rect 9863 34156 9956 34184
rect 9950 34144 9956 34156
rect 10008 34184 10014 34196
rect 11238 34184 11244 34196
rect 10008 34156 11244 34184
rect 10008 34144 10014 34156
rect 11238 34144 11244 34156
rect 11296 34144 11302 34196
rect 1670 34116 1676 34128
rect 1631 34088 1676 34116
rect 1670 34076 1676 34088
rect 1728 34076 1734 34128
rect 10689 34119 10747 34125
rect 10689 34085 10701 34119
rect 10735 34116 10747 34119
rect 10870 34116 10876 34128
rect 10735 34088 10876 34116
rect 10735 34085 10747 34088
rect 10689 34079 10747 34085
rect 10870 34076 10876 34088
rect 10928 34116 10934 34128
rect 11701 34119 11759 34125
rect 11701 34116 11713 34119
rect 10928 34088 11713 34116
rect 10928 34076 10934 34088
rect 11701 34085 11713 34088
rect 11747 34085 11759 34119
rect 11701 34079 11759 34085
rect 12066 34076 12072 34128
rect 12124 34125 12130 34128
rect 12124 34119 12188 34125
rect 12124 34085 12142 34119
rect 12176 34085 12188 34119
rect 12124 34079 12188 34085
rect 12124 34076 12130 34079
rect 1765 34051 1823 34057
rect 1765 34017 1777 34051
rect 1811 34048 1823 34051
rect 1946 34048 1952 34060
rect 1811 34020 1952 34048
rect 1811 34017 1823 34020
rect 1765 34011 1823 34017
rect 1946 34008 1952 34020
rect 2004 34008 2010 34060
rect 2869 34051 2927 34057
rect 2869 34017 2881 34051
rect 2915 34048 2927 34051
rect 3142 34048 3148 34060
rect 2915 34020 3148 34048
rect 2915 34017 2927 34020
rect 2869 34011 2927 34017
rect 3142 34008 3148 34020
rect 3200 34008 3206 34060
rect 4065 34051 4123 34057
rect 4065 34017 4077 34051
rect 4111 34048 4123 34051
rect 4154 34048 4160 34060
rect 4111 34020 4160 34048
rect 4111 34017 4123 34020
rect 4065 34011 4123 34017
rect 4154 34008 4160 34020
rect 4212 34008 4218 34060
rect 4982 34008 4988 34060
rect 5040 34048 5046 34060
rect 5169 34051 5227 34057
rect 5169 34048 5181 34051
rect 5040 34020 5181 34048
rect 5040 34008 5046 34020
rect 5169 34017 5181 34020
rect 5215 34017 5227 34051
rect 5169 34011 5227 34017
rect 6540 34051 6598 34057
rect 6540 34017 6552 34051
rect 6586 34048 6598 34051
rect 7006 34048 7012 34060
rect 6586 34020 7012 34048
rect 6586 34017 6598 34020
rect 6540 34011 6598 34017
rect 7006 34008 7012 34020
rect 7064 34008 7070 34060
rect 10778 34008 10784 34060
rect 10836 34048 10842 34060
rect 11333 34051 11391 34057
rect 11333 34048 11345 34051
rect 10836 34020 11345 34048
rect 10836 34008 10842 34020
rect 11333 34017 11345 34020
rect 11379 34017 11391 34051
rect 11333 34011 11391 34017
rect 6270 33980 6276 33992
rect 6231 33952 6276 33980
rect 6270 33940 6276 33952
rect 6328 33940 6334 33992
rect 10962 33980 10968 33992
rect 10923 33952 10968 33980
rect 10962 33940 10968 33952
rect 11020 33940 11026 33992
rect 11882 33980 11888 33992
rect 11843 33952 11888 33980
rect 11882 33940 11888 33952
rect 11940 33940 11946 33992
rect 4246 33912 4252 33924
rect 4207 33884 4252 33912
rect 4246 33872 4252 33884
rect 4304 33872 4310 33924
rect 10980 33912 11008 33940
rect 10980 33884 11744 33912
rect 3510 33844 3516 33856
rect 3471 33816 3516 33844
rect 3510 33804 3516 33816
rect 3568 33804 3574 33856
rect 4706 33844 4712 33856
rect 4667 33816 4712 33844
rect 4706 33804 4712 33816
rect 4764 33804 4770 33856
rect 7650 33844 7656 33856
rect 7611 33816 7656 33844
rect 7650 33804 7656 33816
rect 7708 33804 7714 33856
rect 10321 33847 10379 33853
rect 10321 33813 10333 33847
rect 10367 33844 10379 33847
rect 11054 33844 11060 33856
rect 10367 33816 11060 33844
rect 10367 33813 10379 33816
rect 10321 33807 10379 33813
rect 11054 33804 11060 33816
rect 11112 33804 11118 33856
rect 11716 33844 11744 33884
rect 13078 33844 13084 33856
rect 11716 33816 13084 33844
rect 13078 33804 13084 33816
rect 13136 33844 13142 33856
rect 13265 33847 13323 33853
rect 13265 33844 13277 33847
rect 13136 33816 13277 33844
rect 13136 33804 13142 33816
rect 13265 33813 13277 33816
rect 13311 33813 13323 33847
rect 13265 33807 13323 33813
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1486 33600 1492 33652
rect 1544 33640 1550 33652
rect 1581 33643 1639 33649
rect 1581 33640 1593 33643
rect 1544 33612 1593 33640
rect 1544 33600 1550 33612
rect 1581 33609 1593 33612
rect 1627 33609 1639 33643
rect 1581 33603 1639 33609
rect 8294 33600 8300 33652
rect 8352 33640 8358 33652
rect 8846 33640 8852 33652
rect 8352 33612 8852 33640
rect 8352 33600 8358 33612
rect 8846 33600 8852 33612
rect 8904 33640 8910 33652
rect 9033 33643 9091 33649
rect 9033 33640 9045 33643
rect 8904 33612 9045 33640
rect 8904 33600 8910 33612
rect 9033 33609 9045 33612
rect 9079 33609 9091 33643
rect 9033 33603 9091 33609
rect 10689 33643 10747 33649
rect 10689 33609 10701 33643
rect 10735 33640 10747 33643
rect 10778 33640 10784 33652
rect 10735 33612 10784 33640
rect 10735 33609 10747 33612
rect 10689 33603 10747 33609
rect 10778 33600 10784 33612
rect 10836 33600 10842 33652
rect 13817 33575 13875 33581
rect 13817 33572 13829 33575
rect 12912 33544 13829 33572
rect 2314 33504 2320 33516
rect 1412 33476 2320 33504
rect 1412 33445 1440 33476
rect 2314 33464 2320 33476
rect 2372 33464 2378 33516
rect 10229 33507 10287 33513
rect 10229 33473 10241 33507
rect 10275 33504 10287 33507
rect 11333 33507 11391 33513
rect 11333 33504 11345 33507
rect 10275 33476 11345 33504
rect 10275 33473 10287 33476
rect 10229 33467 10287 33473
rect 11333 33473 11345 33476
rect 11379 33504 11391 33507
rect 12066 33504 12072 33516
rect 11379 33476 12072 33504
rect 11379 33473 11391 33476
rect 11333 33467 11391 33473
rect 12066 33464 12072 33476
rect 12124 33464 12130 33516
rect 12434 33464 12440 33516
rect 12492 33504 12498 33516
rect 12912 33513 12940 33544
rect 13817 33541 13829 33544
rect 13863 33541 13875 33575
rect 13817 33535 13875 33541
rect 12897 33507 12955 33513
rect 12897 33504 12909 33507
rect 12492 33476 12909 33504
rect 12492 33464 12498 33476
rect 12897 33473 12909 33476
rect 12943 33473 12955 33507
rect 13078 33504 13084 33516
rect 13039 33476 13084 33504
rect 12897 33467 12955 33473
rect 13078 33464 13084 33476
rect 13136 33504 13142 33516
rect 13449 33507 13507 33513
rect 13449 33504 13461 33507
rect 13136 33476 13461 33504
rect 13136 33464 13142 33476
rect 13449 33473 13461 33476
rect 13495 33473 13507 33507
rect 13449 33467 13507 33473
rect 1397 33439 1455 33445
rect 1397 33405 1409 33439
rect 1443 33405 1455 33439
rect 1946 33436 1952 33448
rect 1907 33408 1952 33436
rect 1397 33399 1455 33405
rect 1946 33396 1952 33408
rect 2004 33396 2010 33448
rect 4062 33396 4068 33448
rect 4120 33436 4126 33448
rect 4246 33436 4252 33448
rect 4120 33408 4252 33436
rect 4120 33396 4126 33408
rect 4246 33396 4252 33408
rect 4304 33436 4310 33448
rect 6270 33436 6276 33448
rect 4304 33408 6276 33436
rect 4304 33396 4310 33408
rect 6270 33396 6276 33408
rect 6328 33436 6334 33448
rect 6365 33439 6423 33445
rect 6365 33436 6377 33439
rect 6328 33408 6377 33436
rect 6328 33396 6334 33408
rect 6365 33405 6377 33408
rect 6411 33436 6423 33439
rect 7561 33439 7619 33445
rect 7561 33436 7573 33439
rect 6411 33408 7573 33436
rect 6411 33405 6423 33408
rect 6365 33399 6423 33405
rect 7561 33405 7573 33408
rect 7607 33436 7619 33439
rect 7653 33439 7711 33445
rect 7653 33436 7665 33439
rect 7607 33408 7665 33436
rect 7607 33405 7619 33408
rect 7561 33399 7619 33405
rect 7653 33405 7665 33408
rect 7699 33436 7711 33439
rect 7742 33436 7748 33448
rect 7699 33408 7748 33436
rect 7699 33405 7711 33408
rect 7653 33399 7711 33405
rect 7742 33396 7748 33408
rect 7800 33396 7806 33448
rect 10134 33396 10140 33448
rect 10192 33436 10198 33448
rect 10505 33439 10563 33445
rect 10505 33436 10517 33439
rect 10192 33408 10517 33436
rect 10192 33396 10198 33408
rect 10505 33405 10517 33408
rect 10551 33436 10563 33439
rect 11057 33439 11115 33445
rect 11057 33436 11069 33439
rect 10551 33408 11069 33436
rect 10551 33405 10563 33408
rect 10505 33399 10563 33405
rect 11057 33405 11069 33408
rect 11103 33405 11115 33439
rect 11057 33399 11115 33405
rect 11238 33396 11244 33448
rect 11296 33436 11302 33448
rect 11882 33436 11888 33448
rect 11296 33408 11888 33436
rect 11296 33396 11302 33408
rect 11882 33396 11888 33408
rect 11940 33396 11946 33448
rect 4494 33371 4552 33377
rect 4494 33368 4506 33371
rect 3712 33340 4506 33368
rect 2961 33303 3019 33309
rect 2961 33269 2973 33303
rect 3007 33300 3019 33303
rect 3142 33300 3148 33312
rect 3007 33272 3148 33300
rect 3007 33269 3019 33272
rect 2961 33263 3019 33269
rect 3142 33260 3148 33272
rect 3200 33260 3206 33312
rect 3418 33260 3424 33312
rect 3476 33300 3482 33312
rect 3712 33309 3740 33340
rect 4494 33337 4506 33340
rect 4540 33368 4552 33371
rect 4798 33368 4804 33380
rect 4540 33340 4804 33368
rect 4540 33337 4552 33340
rect 4494 33331 4552 33337
rect 4798 33328 4804 33340
rect 4856 33328 4862 33380
rect 7920 33371 7978 33377
rect 7920 33337 7932 33371
rect 7966 33368 7978 33371
rect 8202 33368 8208 33380
rect 7966 33340 8208 33368
rect 7966 33337 7978 33340
rect 7920 33331 7978 33337
rect 8202 33328 8208 33340
rect 8260 33328 8266 33380
rect 9861 33371 9919 33377
rect 9861 33337 9873 33371
rect 9907 33368 9919 33371
rect 10226 33368 10232 33380
rect 9907 33340 10232 33368
rect 9907 33337 9919 33340
rect 9861 33331 9919 33337
rect 10226 33328 10232 33340
rect 10284 33368 10290 33380
rect 11149 33371 11207 33377
rect 11149 33368 11161 33371
rect 10284 33340 11161 33368
rect 10284 33328 10290 33340
rect 11149 33337 11161 33340
rect 11195 33337 11207 33371
rect 11149 33331 11207 33337
rect 12342 33328 12348 33380
rect 12400 33368 12406 33380
rect 12805 33371 12863 33377
rect 12805 33368 12817 33371
rect 12400 33340 12817 33368
rect 12400 33328 12406 33340
rect 12805 33337 12817 33340
rect 12851 33368 12863 33371
rect 14185 33371 14243 33377
rect 14185 33368 14197 33371
rect 12851 33340 14197 33368
rect 12851 33337 12863 33340
rect 12805 33331 12863 33337
rect 14185 33337 14197 33340
rect 14231 33337 14243 33371
rect 14185 33331 14243 33337
rect 3697 33303 3755 33309
rect 3697 33300 3709 33303
rect 3476 33272 3709 33300
rect 3476 33260 3482 33272
rect 3697 33269 3709 33272
rect 3743 33269 3755 33303
rect 4154 33300 4160 33312
rect 4115 33272 4160 33300
rect 3697 33263 3755 33269
rect 4154 33260 4160 33272
rect 4212 33260 4218 33312
rect 5629 33303 5687 33309
rect 5629 33269 5641 33303
rect 5675 33300 5687 33303
rect 7006 33300 7012 33312
rect 5675 33272 7012 33300
rect 5675 33269 5687 33272
rect 5629 33263 5687 33269
rect 7006 33260 7012 33272
rect 7064 33260 7070 33312
rect 12434 33260 12440 33312
rect 12492 33300 12498 33312
rect 12492 33272 12537 33300
rect 12492 33260 12498 33272
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1578 33096 1584 33108
rect 1539 33068 1584 33096
rect 1578 33056 1584 33068
rect 1636 33056 1642 33108
rect 4246 33096 4252 33108
rect 4207 33068 4252 33096
rect 4246 33056 4252 33068
rect 4304 33056 4310 33108
rect 5905 33099 5963 33105
rect 5905 33065 5917 33099
rect 5951 33096 5963 33099
rect 6638 33096 6644 33108
rect 5951 33068 6644 33096
rect 5951 33065 5963 33068
rect 5905 33059 5963 33065
rect 6638 33056 6644 33068
rect 6696 33096 6702 33108
rect 7101 33099 7159 33105
rect 7101 33096 7113 33099
rect 6696 33068 7113 33096
rect 6696 33056 6702 33068
rect 7101 33065 7113 33068
rect 7147 33065 7159 33099
rect 7558 33096 7564 33108
rect 7519 33068 7564 33096
rect 7101 33059 7159 33065
rect 7558 33056 7564 33068
rect 7616 33056 7622 33108
rect 10778 33096 10784 33108
rect 10739 33068 10784 33096
rect 10778 33056 10784 33068
rect 10836 33056 10842 33108
rect 11054 33056 11060 33108
rect 11112 33096 11118 33108
rect 11241 33099 11299 33105
rect 11241 33096 11253 33099
rect 11112 33068 11253 33096
rect 11112 33056 11118 33068
rect 11241 33065 11253 33068
rect 11287 33065 11299 33099
rect 12342 33096 12348 33108
rect 12303 33068 12348 33096
rect 11241 33059 11299 33065
rect 12342 33056 12348 33068
rect 12400 33056 12406 33108
rect 12805 33099 12863 33105
rect 12805 33065 12817 33099
rect 12851 33096 12863 33099
rect 12894 33096 12900 33108
rect 12851 33068 12900 33096
rect 12851 33065 12863 33068
rect 12805 33059 12863 33065
rect 12894 33056 12900 33068
rect 12952 33096 12958 33108
rect 15746 33096 15752 33108
rect 12952 33068 15752 33096
rect 12952 33056 12958 33068
rect 15746 33056 15752 33068
rect 15804 33056 15810 33108
rect 7282 32988 7288 33040
rect 7340 33028 7346 33040
rect 7466 33028 7472 33040
rect 7340 33000 7472 33028
rect 7340 32988 7346 33000
rect 7466 32988 7472 33000
rect 7524 32988 7530 33040
rect 12066 32988 12072 33040
rect 12124 33028 12130 33040
rect 12124 33000 12940 33028
rect 12124 32988 12130 33000
rect 1397 32963 1455 32969
rect 1397 32929 1409 32963
rect 1443 32960 1455 32963
rect 1670 32960 1676 32972
rect 1443 32932 1676 32960
rect 1443 32929 1455 32932
rect 1397 32923 1455 32929
rect 1670 32920 1676 32932
rect 1728 32920 1734 32972
rect 10042 32920 10048 32972
rect 10100 32960 10106 32972
rect 11149 32963 11207 32969
rect 11149 32960 11161 32963
rect 10100 32932 11161 32960
rect 10100 32920 10106 32932
rect 11149 32929 11161 32932
rect 11195 32960 11207 32963
rect 12342 32960 12348 32972
rect 11195 32932 12348 32960
rect 11195 32929 11207 32932
rect 11149 32923 11207 32929
rect 12342 32920 12348 32932
rect 12400 32920 12406 32972
rect 12710 32960 12716 32972
rect 12671 32932 12716 32960
rect 12710 32920 12716 32932
rect 12768 32920 12774 32972
rect 5994 32892 6000 32904
rect 5955 32864 6000 32892
rect 5994 32852 6000 32864
rect 6052 32852 6058 32904
rect 6178 32892 6184 32904
rect 6139 32864 6184 32892
rect 6178 32852 6184 32864
rect 6236 32852 6242 32904
rect 6546 32852 6552 32904
rect 6604 32892 6610 32904
rect 7006 32892 7012 32904
rect 6604 32864 7012 32892
rect 6604 32852 6610 32864
rect 7006 32852 7012 32864
rect 7064 32892 7070 32904
rect 7653 32895 7711 32901
rect 7653 32892 7665 32895
rect 7064 32864 7665 32892
rect 7064 32852 7070 32864
rect 7653 32861 7665 32864
rect 7699 32861 7711 32895
rect 7653 32855 7711 32861
rect 9582 32852 9588 32904
rect 9640 32892 9646 32904
rect 9677 32895 9735 32901
rect 9677 32892 9689 32895
rect 9640 32864 9689 32892
rect 9640 32852 9646 32864
rect 9677 32861 9689 32864
rect 9723 32861 9735 32895
rect 11422 32892 11428 32904
rect 11383 32864 11428 32892
rect 9677 32855 9735 32861
rect 11422 32852 11428 32864
rect 11480 32852 11486 32904
rect 12912 32901 12940 33000
rect 12897 32895 12955 32901
rect 12897 32861 12909 32895
rect 12943 32861 12955 32895
rect 12897 32855 12955 32861
rect 9125 32827 9183 32833
rect 9125 32793 9137 32827
rect 9171 32824 9183 32827
rect 9490 32824 9496 32836
rect 9171 32796 9496 32824
rect 9171 32793 9183 32796
rect 9125 32787 9183 32793
rect 9490 32784 9496 32796
rect 9548 32784 9554 32836
rect 10778 32784 10784 32836
rect 10836 32824 10842 32836
rect 11146 32824 11152 32836
rect 10836 32796 11152 32824
rect 10836 32784 10842 32796
rect 11146 32784 11152 32796
rect 11204 32784 11210 32836
rect 4982 32716 4988 32768
rect 5040 32756 5046 32768
rect 5169 32759 5227 32765
rect 5169 32756 5181 32759
rect 5040 32728 5181 32756
rect 5040 32716 5046 32728
rect 5169 32725 5181 32728
rect 5215 32725 5227 32759
rect 5534 32756 5540 32768
rect 5495 32728 5540 32756
rect 5169 32719 5227 32725
rect 5534 32716 5540 32728
rect 5592 32716 5598 32768
rect 7006 32756 7012 32768
rect 6967 32728 7012 32756
rect 7006 32716 7012 32728
rect 7064 32716 7070 32768
rect 8205 32759 8263 32765
rect 8205 32725 8217 32759
rect 8251 32756 8263 32759
rect 8294 32756 8300 32768
rect 8251 32728 8300 32756
rect 8251 32725 8263 32728
rect 8205 32719 8263 32725
rect 8294 32716 8300 32728
rect 8352 32716 8358 32768
rect 9398 32756 9404 32768
rect 9359 32728 9404 32756
rect 9398 32716 9404 32728
rect 9456 32716 9462 32768
rect 10413 32759 10471 32765
rect 10413 32725 10425 32759
rect 10459 32756 10471 32759
rect 10962 32756 10968 32768
rect 10459 32728 10968 32756
rect 10459 32725 10471 32728
rect 10413 32719 10471 32725
rect 10962 32716 10968 32728
rect 11020 32756 11026 32768
rect 11514 32756 11520 32768
rect 11020 32728 11520 32756
rect 11020 32716 11026 32728
rect 11514 32716 11520 32728
rect 11572 32716 11578 32768
rect 11977 32759 12035 32765
rect 11977 32725 11989 32759
rect 12023 32756 12035 32759
rect 12066 32756 12072 32768
rect 12023 32728 12072 32756
rect 12023 32725 12035 32728
rect 11977 32719 12035 32725
rect 12066 32716 12072 32728
rect 12124 32716 12130 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 7098 32512 7104 32564
rect 7156 32552 7162 32564
rect 7193 32555 7251 32561
rect 7193 32552 7205 32555
rect 7156 32524 7205 32552
rect 7156 32512 7162 32524
rect 7193 32521 7205 32524
rect 7239 32552 7251 32555
rect 7558 32552 7564 32564
rect 7239 32524 7564 32552
rect 7239 32521 7251 32524
rect 7193 32515 7251 32521
rect 7558 32512 7564 32524
rect 7616 32512 7622 32564
rect 8570 32552 8576 32564
rect 8531 32524 8576 32552
rect 8570 32512 8576 32524
rect 8628 32512 8634 32564
rect 8846 32552 8852 32564
rect 8807 32524 8852 32552
rect 8846 32512 8852 32524
rect 8904 32552 8910 32564
rect 8904 32524 9628 32552
rect 8904 32512 8910 32524
rect 1670 32484 1676 32496
rect 1631 32456 1676 32484
rect 1670 32444 1676 32456
rect 1728 32444 1734 32496
rect 5169 32487 5227 32493
rect 5169 32453 5181 32487
rect 5215 32484 5227 32487
rect 5994 32484 6000 32496
rect 5215 32456 6000 32484
rect 5215 32453 5227 32456
rect 5169 32447 5227 32453
rect 5994 32444 6000 32456
rect 6052 32444 6058 32496
rect 7466 32484 7472 32496
rect 7427 32456 7472 32484
rect 7466 32444 7472 32456
rect 7524 32444 7530 32496
rect 4341 32419 4399 32425
rect 4341 32385 4353 32419
rect 4387 32416 4399 32419
rect 5721 32419 5779 32425
rect 5721 32416 5733 32419
rect 4387 32388 5733 32416
rect 4387 32385 4399 32388
rect 4341 32379 4399 32385
rect 5721 32385 5733 32388
rect 5767 32416 5779 32419
rect 8113 32419 8171 32425
rect 5767 32388 6132 32416
rect 5767 32385 5779 32388
rect 5721 32379 5779 32385
rect 4709 32351 4767 32357
rect 4709 32317 4721 32351
rect 4755 32348 4767 32351
rect 5537 32351 5595 32357
rect 5537 32348 5549 32351
rect 4755 32320 5549 32348
rect 4755 32317 4767 32320
rect 4709 32311 4767 32317
rect 5537 32317 5549 32320
rect 5583 32348 5595 32351
rect 5810 32348 5816 32360
rect 5583 32320 5816 32348
rect 5583 32317 5595 32320
rect 5537 32311 5595 32317
rect 5810 32308 5816 32320
rect 5868 32308 5874 32360
rect 6104 32292 6132 32388
rect 8113 32385 8125 32419
rect 8159 32416 8171 32419
rect 8588 32416 8616 32512
rect 9490 32416 9496 32428
rect 8159 32388 8616 32416
rect 9451 32388 9496 32416
rect 8159 32385 8171 32388
rect 8113 32379 8171 32385
rect 9490 32376 9496 32388
rect 9548 32376 9554 32428
rect 9600 32425 9628 32524
rect 9674 32512 9680 32564
rect 9732 32552 9738 32564
rect 10134 32552 10140 32564
rect 9732 32524 10140 32552
rect 9732 32512 9738 32524
rect 10134 32512 10140 32524
rect 10192 32552 10198 32564
rect 10229 32555 10287 32561
rect 10229 32552 10241 32555
rect 10192 32524 10241 32552
rect 10192 32512 10198 32524
rect 10229 32521 10241 32524
rect 10275 32521 10287 32555
rect 10229 32515 10287 32521
rect 10781 32555 10839 32561
rect 10781 32521 10793 32555
rect 10827 32552 10839 32555
rect 10870 32552 10876 32564
rect 10827 32524 10876 32552
rect 10827 32521 10839 32524
rect 10781 32515 10839 32521
rect 9585 32419 9643 32425
rect 9585 32385 9597 32419
rect 9631 32385 9643 32419
rect 10244 32416 10272 32515
rect 10870 32512 10876 32524
rect 10928 32512 10934 32564
rect 12894 32552 12900 32564
rect 12855 32524 12900 32552
rect 12894 32512 12900 32524
rect 12952 32512 12958 32564
rect 11241 32419 11299 32425
rect 11241 32416 11253 32419
rect 10244 32388 11253 32416
rect 9585 32379 9643 32385
rect 11241 32385 11253 32388
rect 11287 32385 11299 32419
rect 11241 32379 11299 32385
rect 11425 32419 11483 32425
rect 11425 32385 11437 32419
rect 11471 32416 11483 32419
rect 12066 32416 12072 32428
rect 11471 32388 12072 32416
rect 11471 32385 11483 32388
rect 11425 32379 11483 32385
rect 12066 32376 12072 32388
rect 12124 32376 12130 32428
rect 12253 32419 12311 32425
rect 12253 32385 12265 32419
rect 12299 32416 12311 32419
rect 12437 32419 12495 32425
rect 12437 32416 12449 32419
rect 12299 32388 12449 32416
rect 12299 32385 12311 32388
rect 12253 32379 12311 32385
rect 12437 32385 12449 32388
rect 12483 32416 12495 32419
rect 12710 32416 12716 32428
rect 12483 32388 12716 32416
rect 12483 32385 12495 32388
rect 12437 32379 12495 32385
rect 12710 32376 12716 32388
rect 12768 32376 12774 32428
rect 7006 32308 7012 32360
rect 7064 32348 7070 32360
rect 7929 32351 7987 32357
rect 7929 32348 7941 32351
rect 7064 32320 7941 32348
rect 7064 32308 7070 32320
rect 7929 32317 7941 32320
rect 7975 32317 7987 32351
rect 9398 32348 9404 32360
rect 9359 32320 9404 32348
rect 7929 32311 7987 32317
rect 9398 32308 9404 32320
rect 9456 32308 9462 32360
rect 9508 32348 9536 32376
rect 9674 32348 9680 32360
rect 9508 32320 9680 32348
rect 9674 32308 9680 32320
rect 9732 32308 9738 32360
rect 4154 32240 4160 32292
rect 4212 32280 4218 32292
rect 5077 32283 5135 32289
rect 5077 32280 5089 32283
rect 4212 32252 5089 32280
rect 4212 32240 4218 32252
rect 5077 32249 5089 32252
rect 5123 32280 5135 32283
rect 5123 32252 5672 32280
rect 5123 32249 5135 32252
rect 5077 32243 5135 32249
rect 5644 32224 5672 32252
rect 6086 32240 6092 32292
rect 6144 32280 6150 32292
rect 6546 32280 6552 32292
rect 6144 32252 6552 32280
rect 6144 32240 6150 32252
rect 6546 32240 6552 32252
rect 6604 32240 6610 32292
rect 6822 32240 6828 32292
rect 6880 32280 6886 32292
rect 7837 32283 7895 32289
rect 7837 32280 7849 32283
rect 6880 32252 7849 32280
rect 6880 32240 6886 32252
rect 7837 32249 7849 32252
rect 7883 32280 7895 32283
rect 7883 32252 9076 32280
rect 7883 32249 7895 32252
rect 7837 32243 7895 32249
rect 5626 32172 5632 32224
rect 5684 32212 5690 32224
rect 6178 32212 6184 32224
rect 5684 32184 5729 32212
rect 6139 32184 6184 32212
rect 5684 32172 5690 32184
rect 6178 32172 6184 32184
rect 6236 32172 6242 32224
rect 9048 32221 9076 32252
rect 9033 32215 9091 32221
rect 9033 32181 9045 32215
rect 9079 32181 9091 32215
rect 9033 32175 9091 32181
rect 10410 32172 10416 32224
rect 10468 32212 10474 32224
rect 10689 32215 10747 32221
rect 10689 32212 10701 32215
rect 10468 32184 10701 32212
rect 10468 32172 10474 32184
rect 10689 32181 10701 32184
rect 10735 32212 10747 32215
rect 11146 32212 11152 32224
rect 10735 32184 11152 32212
rect 10735 32181 10747 32184
rect 10689 32175 10747 32181
rect 11146 32172 11152 32184
rect 11204 32172 11210 32224
rect 11885 32215 11943 32221
rect 11885 32181 11897 32215
rect 11931 32212 11943 32215
rect 12066 32212 12072 32224
rect 11931 32184 12072 32212
rect 11931 32181 11943 32184
rect 11885 32175 11943 32181
rect 12066 32172 12072 32184
rect 12124 32172 12130 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 5994 32008 6000 32020
rect 5955 31980 6000 32008
rect 5994 31968 6000 31980
rect 6052 31968 6058 32020
rect 6457 32011 6515 32017
rect 6457 31977 6469 32011
rect 6503 32008 6515 32011
rect 6638 32008 6644 32020
rect 6503 31980 6644 32008
rect 6503 31977 6515 31980
rect 6457 31971 6515 31977
rect 6638 31968 6644 31980
rect 6696 31968 6702 32020
rect 6822 32008 6828 32020
rect 6783 31980 6828 32008
rect 6822 31968 6828 31980
rect 6880 31968 6886 32020
rect 7006 31968 7012 32020
rect 7064 32008 7070 32020
rect 7377 32011 7435 32017
rect 7377 32008 7389 32011
rect 7064 31980 7389 32008
rect 7064 31968 7070 31980
rect 7377 31977 7389 31980
rect 7423 31977 7435 32011
rect 10042 32008 10048 32020
rect 10003 31980 10048 32008
rect 7377 31971 7435 31977
rect 10042 31968 10048 31980
rect 10100 31968 10106 32020
rect 10137 32011 10195 32017
rect 10137 31977 10149 32011
rect 10183 32008 10195 32011
rect 10226 32008 10232 32020
rect 10183 31980 10232 32008
rect 10183 31977 10195 31980
rect 10137 31971 10195 31977
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 10502 32008 10508 32020
rect 10463 31980 10508 32008
rect 10502 31968 10508 31980
rect 10560 31968 10566 32020
rect 11054 31968 11060 32020
rect 11112 32008 11118 32020
rect 11517 32011 11575 32017
rect 11517 32008 11529 32011
rect 11112 31980 11529 32008
rect 11112 31968 11118 31980
rect 11517 31977 11529 31980
rect 11563 31977 11575 32011
rect 11517 31971 11575 31977
rect 12066 31968 12072 32020
rect 12124 32008 12130 32020
rect 12437 32011 12495 32017
rect 12437 32008 12449 32011
rect 12124 31980 12449 32008
rect 12124 31968 12130 31980
rect 12437 31977 12449 31980
rect 12483 31977 12495 32011
rect 12437 31971 12495 31977
rect 4246 31940 4252 31952
rect 4080 31912 4252 31940
rect 4080 31884 4108 31912
rect 4246 31900 4252 31912
rect 4304 31900 4310 31952
rect 7193 31943 7251 31949
rect 7193 31909 7205 31943
rect 7239 31940 7251 31943
rect 7282 31940 7288 31952
rect 7239 31912 7288 31940
rect 7239 31909 7251 31912
rect 7193 31903 7251 31909
rect 7282 31900 7288 31912
rect 7340 31900 7346 31952
rect 4062 31872 4068 31884
rect 3975 31844 4068 31872
rect 4062 31832 4068 31844
rect 4120 31832 4126 31884
rect 4332 31875 4390 31881
rect 4332 31841 4344 31875
rect 4378 31872 4390 31875
rect 5074 31872 5080 31884
rect 4378 31844 5080 31872
rect 4378 31841 4390 31844
rect 4332 31835 4390 31841
rect 5074 31832 5080 31844
rect 5132 31832 5138 31884
rect 6178 31832 6184 31884
rect 6236 31872 6242 31884
rect 7742 31872 7748 31884
rect 6236 31844 6592 31872
rect 7703 31844 7748 31872
rect 6236 31832 6242 31844
rect 6564 31736 6592 31844
rect 7742 31832 7748 31844
rect 7800 31832 7806 31884
rect 11241 31875 11299 31881
rect 11241 31841 11253 31875
rect 11287 31872 11299 31875
rect 11422 31872 11428 31884
rect 11287 31844 11428 31872
rect 11287 31841 11299 31844
rect 11241 31835 11299 31841
rect 11422 31832 11428 31844
rect 11480 31872 11486 31884
rect 12342 31872 12348 31884
rect 11480 31844 12348 31872
rect 11480 31832 11486 31844
rect 12342 31832 12348 31844
rect 12400 31832 12406 31884
rect 7558 31764 7564 31816
rect 7616 31804 7622 31816
rect 7837 31807 7895 31813
rect 7837 31804 7849 31807
rect 7616 31776 7849 31804
rect 7616 31764 7622 31776
rect 7837 31773 7849 31776
rect 7883 31773 7895 31807
rect 8018 31804 8024 31816
rect 7931 31776 8024 31804
rect 7837 31767 7895 31773
rect 8018 31764 8024 31776
rect 8076 31804 8082 31816
rect 8846 31804 8852 31816
rect 8076 31776 8852 31804
rect 8076 31764 8082 31776
rect 8846 31764 8852 31776
rect 8904 31764 8910 31816
rect 10410 31764 10416 31816
rect 10468 31804 10474 31816
rect 10597 31807 10655 31813
rect 10597 31804 10609 31807
rect 10468 31776 10609 31804
rect 10468 31764 10474 31776
rect 10597 31773 10609 31776
rect 10643 31773 10655 31807
rect 10778 31804 10784 31816
rect 10739 31776 10784 31804
rect 10597 31767 10655 31773
rect 10778 31764 10784 31776
rect 10836 31764 10842 31816
rect 11146 31764 11152 31816
rect 11204 31804 11210 31816
rect 12066 31804 12072 31816
rect 11204 31776 12072 31804
rect 11204 31764 11210 31776
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 7650 31736 7656 31748
rect 6564 31708 7656 31736
rect 7650 31696 7656 31708
rect 7708 31696 7714 31748
rect 3050 31668 3056 31680
rect 3011 31640 3056 31668
rect 3050 31628 3056 31640
rect 3108 31628 3114 31680
rect 5442 31668 5448 31680
rect 5403 31640 5448 31668
rect 5442 31628 5448 31640
rect 5500 31628 5506 31680
rect 8294 31628 8300 31680
rect 8352 31668 8358 31680
rect 9125 31671 9183 31677
rect 9125 31668 9137 31671
rect 8352 31640 9137 31668
rect 8352 31628 8358 31640
rect 9125 31637 9137 31640
rect 9171 31668 9183 31671
rect 9306 31668 9312 31680
rect 9171 31640 9312 31668
rect 9171 31637 9183 31640
rect 9125 31631 9183 31637
rect 9306 31628 9312 31640
rect 9364 31628 9370 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 4062 31464 4068 31476
rect 4023 31436 4068 31464
rect 4062 31424 4068 31436
rect 4120 31424 4126 31476
rect 4614 31424 4620 31476
rect 4672 31464 4678 31476
rect 4890 31464 4896 31476
rect 4672 31436 4896 31464
rect 4672 31424 4678 31436
rect 4890 31424 4896 31436
rect 4948 31424 4954 31476
rect 4982 31424 4988 31476
rect 5040 31464 5046 31476
rect 5350 31464 5356 31476
rect 5040 31436 5356 31464
rect 5040 31424 5046 31436
rect 5350 31424 5356 31436
rect 5408 31424 5414 31476
rect 7742 31424 7748 31476
rect 7800 31464 7806 31476
rect 8113 31467 8171 31473
rect 8113 31464 8125 31467
rect 7800 31436 8125 31464
rect 7800 31424 7806 31436
rect 8113 31433 8125 31436
rect 8159 31433 8171 31467
rect 8113 31427 8171 31433
rect 9125 31467 9183 31473
rect 9125 31433 9137 31467
rect 9171 31464 9183 31467
rect 9398 31464 9404 31476
rect 9171 31436 9404 31464
rect 9171 31433 9183 31436
rect 9125 31427 9183 31433
rect 9398 31424 9404 31436
rect 9456 31424 9462 31476
rect 10778 31424 10784 31476
rect 10836 31464 10842 31476
rect 10873 31467 10931 31473
rect 10873 31464 10885 31467
rect 10836 31436 10885 31464
rect 10836 31424 10842 31436
rect 10873 31433 10885 31436
rect 10919 31433 10931 31467
rect 13722 31464 13728 31476
rect 13683 31436 13728 31464
rect 10873 31427 10931 31433
rect 13722 31424 13728 31436
rect 13780 31424 13786 31476
rect 7469 31399 7527 31405
rect 7469 31365 7481 31399
rect 7515 31396 7527 31399
rect 8018 31396 8024 31408
rect 7515 31368 8024 31396
rect 7515 31365 7527 31368
rect 7469 31359 7527 31365
rect 8018 31356 8024 31368
rect 8076 31356 8082 31408
rect 2869 31331 2927 31337
rect 2869 31297 2881 31331
rect 2915 31328 2927 31331
rect 3510 31328 3516 31340
rect 2915 31300 3516 31328
rect 2915 31297 2927 31300
rect 2869 31291 2927 31297
rect 3510 31288 3516 31300
rect 3568 31328 3574 31340
rect 3605 31331 3663 31337
rect 3605 31328 3617 31331
rect 3568 31300 3617 31328
rect 3568 31288 3574 31300
rect 3605 31297 3617 31300
rect 3651 31328 3663 31331
rect 4614 31328 4620 31340
rect 3651 31300 4620 31328
rect 3651 31297 3663 31300
rect 3605 31291 3663 31297
rect 4614 31288 4620 31300
rect 4672 31288 4678 31340
rect 5074 31328 5080 31340
rect 5035 31300 5080 31328
rect 5074 31288 5080 31300
rect 5132 31288 5138 31340
rect 8570 31288 8576 31340
rect 8628 31328 8634 31340
rect 8754 31328 8760 31340
rect 8628 31300 8760 31328
rect 8628 31288 8634 31300
rect 8754 31288 8760 31300
rect 8812 31288 8818 31340
rect 9306 31288 9312 31340
rect 9364 31328 9370 31340
rect 9677 31331 9735 31337
rect 9677 31328 9689 31331
rect 9364 31300 9689 31328
rect 9364 31288 9370 31300
rect 9677 31297 9689 31300
rect 9723 31328 9735 31331
rect 10226 31328 10232 31340
rect 9723 31300 10232 31328
rect 9723 31297 9735 31300
rect 9677 31291 9735 31297
rect 10226 31288 10232 31300
rect 10284 31288 10290 31340
rect 12618 31288 12624 31340
rect 12676 31328 12682 31340
rect 12894 31328 12900 31340
rect 12676 31300 12900 31328
rect 12676 31288 12682 31300
rect 12894 31288 12900 31300
rect 12952 31288 12958 31340
rect 4433 31263 4491 31269
rect 4433 31229 4445 31263
rect 4479 31260 4491 31263
rect 4982 31260 4988 31272
rect 4479 31232 4988 31260
rect 4479 31229 4491 31232
rect 4433 31223 4491 31229
rect 4982 31220 4988 31232
rect 5040 31220 5046 31272
rect 9493 31263 9551 31269
rect 9493 31229 9505 31263
rect 9539 31260 9551 31263
rect 9582 31260 9588 31272
rect 9539 31232 9588 31260
rect 9539 31229 9551 31232
rect 9493 31223 9551 31229
rect 9582 31220 9588 31232
rect 9640 31220 9646 31272
rect 13538 31260 13544 31272
rect 13499 31232 13544 31260
rect 13538 31220 13544 31232
rect 13596 31260 13602 31272
rect 14001 31263 14059 31269
rect 14001 31260 14013 31263
rect 13596 31232 14013 31260
rect 13596 31220 13602 31232
rect 14001 31229 14013 31232
rect 14047 31229 14059 31263
rect 14001 31223 14059 31229
rect 2406 31152 2412 31204
rect 2464 31192 2470 31204
rect 2501 31195 2559 31201
rect 2501 31192 2513 31195
rect 2464 31164 2513 31192
rect 2464 31152 2470 31164
rect 2501 31161 2513 31164
rect 2547 31192 2559 31195
rect 3329 31195 3387 31201
rect 3329 31192 3341 31195
rect 2547 31164 3341 31192
rect 2547 31161 2559 31164
rect 2501 31155 2559 31161
rect 3329 31161 3341 31164
rect 3375 31161 3387 31195
rect 3329 31155 3387 31161
rect 4154 31152 4160 31204
rect 4212 31192 4218 31204
rect 4893 31195 4951 31201
rect 4893 31192 4905 31195
rect 4212 31164 4905 31192
rect 4212 31152 4218 31164
rect 4893 31161 4905 31164
rect 4939 31192 4951 31195
rect 5537 31195 5595 31201
rect 5537 31192 5549 31195
rect 4939 31164 5549 31192
rect 4939 31161 4951 31164
rect 4893 31155 4951 31161
rect 5537 31161 5549 31164
rect 5583 31161 5595 31195
rect 5537 31155 5595 31161
rect 2958 31124 2964 31136
rect 2919 31096 2964 31124
rect 2958 31084 2964 31096
rect 3016 31084 3022 31136
rect 3050 31084 3056 31136
rect 3108 31124 3114 31136
rect 3421 31127 3479 31133
rect 3421 31124 3433 31127
rect 3108 31096 3433 31124
rect 3108 31084 3114 31096
rect 3421 31093 3433 31096
rect 3467 31093 3479 31127
rect 3421 31087 3479 31093
rect 4430 31084 4436 31136
rect 4488 31124 4494 31136
rect 4525 31127 4583 31133
rect 4525 31124 4537 31127
rect 4488 31096 4537 31124
rect 4488 31084 4494 31096
rect 4525 31093 4537 31096
rect 4571 31093 4583 31127
rect 4525 31087 4583 31093
rect 7558 31084 7564 31136
rect 7616 31124 7622 31136
rect 7745 31127 7803 31133
rect 7745 31124 7757 31127
rect 7616 31096 7757 31124
rect 7616 31084 7622 31096
rect 7745 31093 7757 31096
rect 7791 31093 7803 31127
rect 7745 31087 7803 31093
rect 9033 31127 9091 31133
rect 9033 31093 9045 31127
rect 9079 31124 9091 31127
rect 9306 31124 9312 31136
rect 9079 31096 9312 31124
rect 9079 31093 9091 31096
rect 9033 31087 9091 31093
rect 9306 31084 9312 31096
rect 9364 31124 9370 31136
rect 9585 31127 9643 31133
rect 9585 31124 9597 31127
rect 9364 31096 9597 31124
rect 9364 31084 9370 31096
rect 9585 31093 9597 31096
rect 9631 31093 9643 31127
rect 9585 31087 9643 31093
rect 9950 31084 9956 31136
rect 10008 31124 10014 31136
rect 10137 31127 10195 31133
rect 10137 31124 10149 31127
rect 10008 31096 10149 31124
rect 10008 31084 10014 31096
rect 10137 31093 10149 31096
rect 10183 31124 10195 31127
rect 10410 31124 10416 31136
rect 10183 31096 10416 31124
rect 10183 31093 10195 31096
rect 10137 31087 10195 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10502 31084 10508 31136
rect 10560 31124 10566 31136
rect 10597 31127 10655 31133
rect 10597 31124 10609 31127
rect 10560 31096 10609 31124
rect 10560 31084 10566 31096
rect 10597 31093 10609 31096
rect 10643 31124 10655 31127
rect 10962 31124 10968 31136
rect 10643 31096 10968 31124
rect 10643 31093 10655 31096
rect 10597 31087 10655 31093
rect 10962 31084 10968 31096
rect 11020 31084 11026 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 2406 30920 2412 30932
rect 2367 30892 2412 30920
rect 2406 30880 2412 30892
rect 2464 30880 2470 30932
rect 2774 30880 2780 30932
rect 2832 30920 2838 30932
rect 5534 30920 5540 30932
rect 2832 30892 2877 30920
rect 5495 30892 5540 30920
rect 2832 30880 2838 30892
rect 5534 30880 5540 30892
rect 5592 30880 5598 30932
rect 6733 30923 6791 30929
rect 6733 30889 6745 30923
rect 6779 30920 6791 30923
rect 6822 30920 6828 30932
rect 6779 30892 6828 30920
rect 6779 30889 6791 30892
rect 6733 30883 6791 30889
rect 6822 30880 6828 30892
rect 6880 30880 6886 30932
rect 7469 30923 7527 30929
rect 7469 30889 7481 30923
rect 7515 30920 7527 30923
rect 7650 30920 7656 30932
rect 7515 30892 7656 30920
rect 7515 30889 7527 30892
rect 7469 30883 7527 30889
rect 7650 30880 7656 30892
rect 7708 30880 7714 30932
rect 7742 30880 7748 30932
rect 7800 30920 7806 30932
rect 7929 30923 7987 30929
rect 7929 30920 7941 30923
rect 7800 30892 7941 30920
rect 7800 30880 7806 30892
rect 7929 30889 7941 30892
rect 7975 30889 7987 30923
rect 7929 30883 7987 30889
rect 8110 30880 8116 30932
rect 8168 30920 8174 30932
rect 8297 30923 8355 30929
rect 8297 30920 8309 30923
rect 8168 30892 8309 30920
rect 8168 30880 8174 30892
rect 8297 30889 8309 30892
rect 8343 30889 8355 30923
rect 9674 30920 9680 30932
rect 9635 30892 9680 30920
rect 8297 30883 8355 30889
rect 9674 30880 9680 30892
rect 9732 30880 9738 30932
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 12897 30923 12955 30929
rect 12897 30920 12909 30923
rect 12492 30892 12909 30920
rect 12492 30880 12498 30892
rect 12897 30889 12909 30892
rect 12943 30889 12955 30923
rect 12897 30883 12955 30889
rect 2222 30812 2228 30864
rect 2280 30852 2286 30864
rect 2869 30855 2927 30861
rect 2869 30852 2881 30855
rect 2280 30824 2881 30852
rect 2280 30812 2286 30824
rect 2869 30821 2881 30824
rect 2915 30852 2927 30855
rect 8570 30852 8576 30864
rect 2915 30824 8576 30852
rect 2915 30821 2927 30824
rect 2869 30815 2927 30821
rect 8570 30812 8576 30824
rect 8628 30812 8634 30864
rect 9217 30855 9275 30861
rect 9217 30821 9229 30855
rect 9263 30852 9275 30855
rect 9582 30852 9588 30864
rect 9263 30824 9588 30852
rect 9263 30821 9275 30824
rect 9217 30815 9275 30821
rect 9582 30812 9588 30824
rect 9640 30812 9646 30864
rect 11514 30812 11520 30864
rect 11572 30852 11578 30864
rect 11762 30855 11820 30861
rect 11762 30852 11774 30855
rect 11572 30824 11774 30852
rect 11572 30812 11578 30824
rect 11762 30821 11774 30824
rect 11808 30821 11820 30855
rect 11762 30815 11820 30821
rect 4338 30744 4344 30796
rect 4396 30784 4402 30796
rect 4433 30787 4491 30793
rect 4433 30784 4445 30787
rect 4396 30756 4445 30784
rect 4396 30744 4402 30756
rect 4433 30753 4445 30756
rect 4479 30753 4491 30787
rect 10042 30784 10048 30796
rect 10003 30756 10048 30784
rect 4433 30747 4491 30753
rect 10042 30744 10048 30756
rect 10100 30744 10106 30796
rect 10137 30787 10195 30793
rect 10137 30753 10149 30787
rect 10183 30784 10195 30787
rect 10686 30784 10692 30796
rect 10183 30756 10692 30784
rect 10183 30753 10195 30756
rect 10137 30747 10195 30753
rect 10686 30744 10692 30756
rect 10744 30744 10750 30796
rect 2866 30676 2872 30728
rect 2924 30716 2930 30728
rect 2961 30719 3019 30725
rect 2961 30716 2973 30719
rect 2924 30688 2973 30716
rect 2924 30676 2930 30688
rect 2961 30685 2973 30688
rect 3007 30716 3019 30719
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 3007 30688 3801 30716
rect 3007 30685 3019 30688
rect 2961 30679 3019 30685
rect 3789 30685 3801 30688
rect 3835 30716 3847 30719
rect 4522 30716 4528 30728
rect 3835 30688 4384 30716
rect 4483 30688 4528 30716
rect 3835 30685 3847 30688
rect 3789 30679 3847 30685
rect 3234 30608 3240 30660
rect 3292 30648 3298 30660
rect 3513 30651 3571 30657
rect 3513 30648 3525 30651
rect 3292 30620 3525 30648
rect 3292 30608 3298 30620
rect 3513 30617 3525 30620
rect 3559 30648 3571 30651
rect 4065 30651 4123 30657
rect 4065 30648 4077 30651
rect 3559 30620 4077 30648
rect 3559 30617 3571 30620
rect 3513 30611 3571 30617
rect 4065 30617 4077 30620
rect 4111 30617 4123 30651
rect 4356 30648 4384 30688
rect 4522 30676 4528 30688
rect 4580 30676 4586 30728
rect 4614 30676 4620 30728
rect 4672 30716 4678 30728
rect 4709 30719 4767 30725
rect 4709 30716 4721 30719
rect 4672 30688 4721 30716
rect 4672 30676 4678 30688
rect 4709 30685 4721 30688
rect 4755 30716 4767 30719
rect 5442 30716 5448 30728
rect 4755 30688 5448 30716
rect 4755 30685 4767 30688
rect 4709 30679 4767 30685
rect 5442 30676 5448 30688
rect 5500 30676 5506 30728
rect 6178 30676 6184 30728
rect 6236 30716 6242 30728
rect 6825 30719 6883 30725
rect 6825 30716 6837 30719
rect 6236 30688 6837 30716
rect 6236 30676 6242 30688
rect 6825 30685 6837 30688
rect 6871 30685 6883 30719
rect 6825 30679 6883 30685
rect 6917 30719 6975 30725
rect 6917 30685 6929 30719
rect 6963 30685 6975 30719
rect 8386 30716 8392 30728
rect 8347 30688 8392 30716
rect 6917 30679 6975 30685
rect 4982 30648 4988 30660
rect 4356 30620 4988 30648
rect 4065 30611 4123 30617
rect 4982 30608 4988 30620
rect 5040 30648 5046 30660
rect 5077 30651 5135 30657
rect 5077 30648 5089 30651
rect 5040 30620 5089 30648
rect 5040 30608 5046 30620
rect 5077 30617 5089 30620
rect 5123 30617 5135 30651
rect 5077 30611 5135 30617
rect 6086 30608 6092 30660
rect 6144 30648 6150 30660
rect 6638 30648 6644 30660
rect 6144 30620 6644 30648
rect 6144 30608 6150 30620
rect 6638 30608 6644 30620
rect 6696 30648 6702 30660
rect 6932 30648 6960 30679
rect 8386 30676 8392 30688
rect 8444 30676 8450 30728
rect 8481 30719 8539 30725
rect 8481 30685 8493 30719
rect 8527 30685 8539 30719
rect 8481 30679 8539 30685
rect 6696 30620 6960 30648
rect 6696 30608 6702 30620
rect 8294 30608 8300 30660
rect 8352 30648 8358 30660
rect 8496 30648 8524 30679
rect 10226 30676 10232 30728
rect 10284 30716 10290 30728
rect 10284 30688 10329 30716
rect 10284 30676 10290 30688
rect 11238 30676 11244 30728
rect 11296 30716 11302 30728
rect 11422 30716 11428 30728
rect 11296 30688 11428 30716
rect 11296 30676 11302 30688
rect 11422 30676 11428 30688
rect 11480 30716 11486 30728
rect 11517 30719 11575 30725
rect 11517 30716 11529 30719
rect 11480 30688 11529 30716
rect 11480 30676 11486 30688
rect 11517 30685 11529 30688
rect 11563 30685 11575 30719
rect 11517 30679 11575 30685
rect 8352 30620 8524 30648
rect 8352 30608 8358 30620
rect 5810 30580 5816 30592
rect 5771 30552 5816 30580
rect 5810 30540 5816 30552
rect 5868 30540 5874 30592
rect 6365 30583 6423 30589
rect 6365 30549 6377 30583
rect 6411 30580 6423 30583
rect 6914 30580 6920 30592
rect 6411 30552 6920 30580
rect 6411 30549 6423 30552
rect 6365 30543 6423 30549
rect 6914 30540 6920 30552
rect 6972 30540 6978 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 2133 30379 2191 30385
rect 2133 30345 2145 30379
rect 2179 30376 2191 30379
rect 2222 30376 2228 30388
rect 2179 30348 2228 30376
rect 2179 30345 2191 30348
rect 2133 30339 2191 30345
rect 2222 30336 2228 30348
rect 2280 30336 2286 30388
rect 4157 30379 4215 30385
rect 4157 30345 4169 30379
rect 4203 30376 4215 30379
rect 4614 30376 4620 30388
rect 4203 30348 4620 30376
rect 4203 30345 4215 30348
rect 4157 30339 4215 30345
rect 4614 30336 4620 30348
rect 4672 30336 4678 30388
rect 6178 30376 6184 30388
rect 6139 30348 6184 30376
rect 6178 30336 6184 30348
rect 6236 30336 6242 30388
rect 10226 30336 10232 30388
rect 10284 30376 10290 30388
rect 10965 30379 11023 30385
rect 10965 30376 10977 30379
rect 10284 30348 10977 30376
rect 10284 30336 10290 30348
rect 10965 30345 10977 30348
rect 11011 30345 11023 30379
rect 10965 30339 11023 30345
rect 11514 30336 11520 30388
rect 11572 30376 11578 30388
rect 11885 30379 11943 30385
rect 11885 30376 11897 30379
rect 11572 30348 11897 30376
rect 11572 30336 11578 30348
rect 11885 30345 11897 30348
rect 11931 30345 11943 30379
rect 11885 30339 11943 30345
rect 7834 30268 7840 30320
rect 7892 30308 7898 30320
rect 8021 30311 8079 30317
rect 8021 30308 8033 30311
rect 7892 30280 8033 30308
rect 7892 30268 7898 30280
rect 8021 30277 8033 30280
rect 8067 30308 8079 30311
rect 8110 30308 8116 30320
rect 8067 30280 8116 30308
rect 8067 30277 8079 30280
rect 8021 30271 8079 30277
rect 8110 30268 8116 30280
rect 8168 30268 8174 30320
rect 9766 30268 9772 30320
rect 9824 30308 9830 30320
rect 10042 30308 10048 30320
rect 9824 30280 10048 30308
rect 9824 30268 9830 30280
rect 10042 30268 10048 30280
rect 10100 30268 10106 30320
rect 2958 30200 2964 30252
rect 3016 30240 3022 30252
rect 3329 30243 3387 30249
rect 3329 30240 3341 30243
rect 3016 30212 3341 30240
rect 3016 30200 3022 30212
rect 3329 30209 3341 30212
rect 3375 30209 3387 30243
rect 3329 30203 3387 30209
rect 3418 30200 3424 30252
rect 3476 30240 3482 30252
rect 3476 30212 3521 30240
rect 3476 30200 3482 30212
rect 5534 30200 5540 30252
rect 5592 30240 5598 30252
rect 5629 30243 5687 30249
rect 5629 30240 5641 30243
rect 5592 30212 5641 30240
rect 5592 30200 5598 30212
rect 5629 30209 5641 30212
rect 5675 30209 5687 30243
rect 5629 30203 5687 30209
rect 5813 30243 5871 30249
rect 5813 30209 5825 30243
rect 5859 30240 5871 30243
rect 5994 30240 6000 30252
rect 5859 30212 6000 30240
rect 5859 30209 5871 30212
rect 5813 30203 5871 30209
rect 5994 30200 6000 30212
rect 6052 30200 6058 30252
rect 6914 30200 6920 30252
rect 6972 30240 6978 30252
rect 7282 30240 7288 30252
rect 6972 30212 7288 30240
rect 6972 30200 6978 30212
rect 7282 30200 7288 30212
rect 7340 30200 7346 30252
rect 7469 30243 7527 30249
rect 7469 30209 7481 30243
rect 7515 30240 7527 30243
rect 7650 30240 7656 30252
rect 7515 30212 7656 30240
rect 7515 30209 7527 30212
rect 7469 30203 7527 30209
rect 7650 30200 7656 30212
rect 7708 30200 7714 30252
rect 8757 30243 8815 30249
rect 8757 30209 8769 30243
rect 8803 30240 8815 30243
rect 10229 30243 10287 30249
rect 10229 30240 10241 30243
rect 8803 30212 10241 30240
rect 8803 30209 8815 30212
rect 8757 30203 8815 30209
rect 10229 30209 10241 30212
rect 10275 30240 10287 30243
rect 10502 30240 10508 30252
rect 10275 30212 10508 30240
rect 10275 30209 10287 30212
rect 10229 30203 10287 30209
rect 10502 30200 10508 30212
rect 10560 30200 10566 30252
rect 3234 30172 3240 30184
rect 3195 30144 3240 30172
rect 3234 30132 3240 30144
rect 3292 30132 3298 30184
rect 5902 30132 5908 30184
rect 5960 30172 5966 30184
rect 6641 30175 6699 30181
rect 6641 30172 6653 30175
rect 5960 30144 6653 30172
rect 5960 30132 5966 30144
rect 6641 30141 6653 30144
rect 6687 30172 6699 30175
rect 6687 30144 7236 30172
rect 6687 30141 6699 30144
rect 6641 30135 6699 30141
rect 5537 30107 5595 30113
rect 5537 30073 5549 30107
rect 5583 30104 5595 30107
rect 5810 30104 5816 30116
rect 5583 30076 5816 30104
rect 5583 30073 5595 30076
rect 5537 30067 5595 30073
rect 5810 30064 5816 30076
rect 5868 30104 5874 30116
rect 5868 30076 6868 30104
rect 5868 30064 5874 30076
rect 2498 30036 2504 30048
rect 2459 30008 2504 30036
rect 2498 29996 2504 30008
rect 2556 29996 2562 30048
rect 2866 30036 2872 30048
rect 2827 30008 2872 30036
rect 2866 29996 2872 30008
rect 2924 29996 2930 30048
rect 4522 30036 4528 30048
rect 4483 30008 4528 30036
rect 4522 29996 4528 30008
rect 4580 29996 4586 30048
rect 4982 30036 4988 30048
rect 4943 30008 4988 30036
rect 4982 29996 4988 30008
rect 5040 29996 5046 30048
rect 5166 30036 5172 30048
rect 5127 30008 5172 30036
rect 5166 29996 5172 30008
rect 5224 29996 5230 30048
rect 6840 30045 6868 30076
rect 7208 30048 7236 30144
rect 7926 30132 7932 30184
rect 7984 30172 7990 30184
rect 9766 30172 9772 30184
rect 7984 30144 9772 30172
rect 7984 30132 7990 30144
rect 9766 30132 9772 30144
rect 9824 30132 9830 30184
rect 9493 30107 9551 30113
rect 9493 30073 9505 30107
rect 9539 30104 9551 30107
rect 9674 30104 9680 30116
rect 9539 30076 9680 30104
rect 9539 30073 9551 30076
rect 9493 30067 9551 30073
rect 9674 30064 9680 30076
rect 9732 30104 9738 30116
rect 10045 30107 10103 30113
rect 10045 30104 10057 30107
rect 9732 30076 10057 30104
rect 9732 30064 9738 30076
rect 10045 30073 10057 30076
rect 10091 30073 10103 30107
rect 10045 30067 10103 30073
rect 10226 30064 10232 30116
rect 10284 30104 10290 30116
rect 11422 30104 11428 30116
rect 10284 30076 11428 30104
rect 10284 30064 10290 30076
rect 11422 30064 11428 30076
rect 11480 30104 11486 30116
rect 11517 30107 11575 30113
rect 11517 30104 11529 30107
rect 11480 30076 11529 30104
rect 11480 30064 11486 30076
rect 11517 30073 11529 30076
rect 11563 30073 11575 30107
rect 11517 30067 11575 30073
rect 6825 30039 6883 30045
rect 6825 30005 6837 30039
rect 6871 30005 6883 30039
rect 7190 30036 7196 30048
rect 7151 30008 7196 30036
rect 6825 29999 6883 30005
rect 7190 29996 7196 30008
rect 7248 29996 7254 30048
rect 8294 30036 8300 30048
rect 8255 30008 8300 30036
rect 8294 29996 8300 30008
rect 8352 29996 8358 30048
rect 8754 29996 8760 30048
rect 8812 30036 8818 30048
rect 9033 30039 9091 30045
rect 9033 30036 9045 30039
rect 8812 30008 9045 30036
rect 8812 29996 8818 30008
rect 9033 30005 9045 30008
rect 9079 30005 9091 30039
rect 9582 30036 9588 30048
rect 9543 30008 9588 30036
rect 9033 29999 9091 30005
rect 9582 29996 9588 30008
rect 9640 29996 9646 30048
rect 9766 29996 9772 30048
rect 9824 30036 9830 30048
rect 9953 30039 10011 30045
rect 9953 30036 9965 30039
rect 9824 30008 9965 30036
rect 9824 29996 9830 30008
rect 9953 30005 9965 30008
rect 9999 30005 10011 30039
rect 10686 30036 10692 30048
rect 10647 30008 10692 30036
rect 9953 29999 10011 30005
rect 10686 29996 10692 30008
rect 10744 29996 10750 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 2958 29792 2964 29844
rect 3016 29832 3022 29844
rect 3237 29835 3295 29841
rect 3237 29832 3249 29835
rect 3016 29804 3249 29832
rect 3016 29792 3022 29804
rect 3237 29801 3249 29804
rect 3283 29801 3295 29835
rect 4338 29832 4344 29844
rect 4299 29804 4344 29832
rect 3237 29795 3295 29801
rect 4338 29792 4344 29804
rect 4396 29792 4402 29844
rect 6914 29832 6920 29844
rect 6875 29804 6920 29832
rect 6914 29792 6920 29804
rect 6972 29792 6978 29844
rect 7282 29792 7288 29844
rect 7340 29832 7346 29844
rect 7561 29835 7619 29841
rect 7561 29832 7573 29835
rect 7340 29804 7573 29832
rect 7340 29792 7346 29804
rect 7561 29801 7573 29804
rect 7607 29801 7619 29835
rect 7561 29795 7619 29801
rect 6638 29724 6644 29776
rect 6696 29764 6702 29776
rect 7193 29767 7251 29773
rect 7193 29764 7205 29767
rect 6696 29736 7205 29764
rect 6696 29724 6702 29736
rect 7193 29733 7205 29736
rect 7239 29733 7251 29767
rect 7193 29727 7251 29733
rect 1397 29699 1455 29705
rect 1397 29665 1409 29699
rect 1443 29696 1455 29699
rect 2314 29696 2320 29708
rect 1443 29668 2320 29696
rect 1443 29665 1455 29668
rect 1397 29659 1455 29665
rect 2314 29656 2320 29668
rect 2372 29656 2378 29708
rect 2961 29699 3019 29705
rect 2961 29665 2973 29699
rect 3007 29696 3019 29699
rect 3418 29696 3424 29708
rect 3007 29668 3424 29696
rect 3007 29665 3019 29668
rect 2961 29659 3019 29665
rect 3418 29656 3424 29668
rect 3476 29656 3482 29708
rect 4982 29656 4988 29708
rect 5040 29696 5046 29708
rect 5160 29699 5218 29705
rect 5160 29696 5172 29699
rect 5040 29668 5172 29696
rect 5040 29656 5046 29668
rect 5160 29665 5172 29668
rect 5206 29696 5218 29699
rect 5994 29696 6000 29708
rect 5206 29668 6000 29696
rect 5206 29665 5218 29668
rect 5160 29659 5218 29665
rect 5994 29656 6000 29668
rect 6052 29656 6058 29708
rect 8018 29656 8024 29708
rect 8076 29696 8082 29708
rect 8113 29699 8171 29705
rect 8113 29696 8125 29699
rect 8076 29668 8125 29696
rect 8076 29656 8082 29668
rect 8113 29665 8125 29668
rect 8159 29696 8171 29699
rect 8662 29696 8668 29708
rect 8159 29668 8668 29696
rect 8159 29665 8171 29668
rect 8113 29659 8171 29665
rect 8662 29656 8668 29668
rect 8720 29656 8726 29708
rect 10502 29705 10508 29708
rect 10496 29696 10508 29705
rect 10463 29668 10508 29696
rect 10496 29659 10508 29668
rect 10502 29656 10508 29659
rect 10560 29656 10566 29708
rect 4798 29588 4804 29640
rect 4856 29628 4862 29640
rect 4893 29631 4951 29637
rect 4893 29628 4905 29631
rect 4856 29600 4905 29628
rect 4856 29588 4862 29600
rect 4893 29597 4905 29600
rect 4939 29597 4951 29631
rect 4893 29591 4951 29597
rect 7742 29588 7748 29640
rect 7800 29628 7806 29640
rect 8205 29631 8263 29637
rect 8205 29628 8217 29631
rect 7800 29600 8217 29628
rect 7800 29588 7806 29600
rect 8205 29597 8217 29600
rect 8251 29597 8263 29631
rect 8205 29591 8263 29597
rect 8389 29631 8447 29637
rect 8389 29597 8401 29631
rect 8435 29628 8447 29631
rect 8570 29628 8576 29640
rect 8435 29600 8576 29628
rect 8435 29597 8447 29600
rect 8389 29591 8447 29597
rect 8570 29588 8576 29600
rect 8628 29588 8634 29640
rect 10226 29628 10232 29640
rect 10187 29600 10232 29628
rect 10226 29588 10232 29600
rect 10284 29588 10290 29640
rect 2501 29495 2559 29501
rect 2501 29461 2513 29495
rect 2547 29492 2559 29495
rect 2774 29492 2780 29504
rect 2547 29464 2780 29492
rect 2547 29461 2559 29464
rect 2501 29455 2559 29461
rect 2774 29452 2780 29464
rect 2832 29452 2838 29504
rect 6270 29492 6276 29504
rect 6231 29464 6276 29492
rect 6270 29452 6276 29464
rect 6328 29452 6334 29504
rect 7745 29495 7803 29501
rect 7745 29461 7757 29495
rect 7791 29492 7803 29495
rect 7926 29492 7932 29504
rect 7791 29464 7932 29492
rect 7791 29461 7803 29464
rect 7745 29455 7803 29461
rect 7926 29452 7932 29464
rect 7984 29452 7990 29504
rect 8386 29452 8392 29504
rect 8444 29492 8450 29504
rect 8849 29495 8907 29501
rect 8849 29492 8861 29495
rect 8444 29464 8861 29492
rect 8444 29452 8450 29464
rect 8849 29461 8861 29464
rect 8895 29492 8907 29495
rect 9398 29492 9404 29504
rect 8895 29464 9404 29492
rect 8895 29461 8907 29464
rect 8849 29455 8907 29461
rect 9398 29452 9404 29464
rect 9456 29452 9462 29504
rect 9766 29452 9772 29504
rect 9824 29492 9830 29504
rect 9861 29495 9919 29501
rect 9861 29492 9873 29495
rect 9824 29464 9873 29492
rect 9824 29452 9830 29464
rect 9861 29461 9873 29464
rect 9907 29461 9919 29495
rect 11606 29492 11612 29504
rect 11567 29464 11612 29492
rect 9861 29455 9919 29461
rect 11606 29452 11612 29464
rect 11664 29452 11670 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 1578 29288 1584 29300
rect 1539 29260 1584 29288
rect 1578 29248 1584 29260
rect 1636 29248 1642 29300
rect 1949 29291 2007 29297
rect 1949 29257 1961 29291
rect 1995 29288 2007 29291
rect 2866 29288 2872 29300
rect 1995 29260 2872 29288
rect 1995 29257 2007 29260
rect 1949 29251 2007 29257
rect 1397 29087 1455 29093
rect 1397 29053 1409 29087
rect 1443 29084 1455 29087
rect 1964 29084 1992 29251
rect 2866 29248 2872 29260
rect 2924 29248 2930 29300
rect 4798 29248 4804 29300
rect 4856 29288 4862 29300
rect 4985 29291 5043 29297
rect 4985 29288 4997 29291
rect 4856 29260 4997 29288
rect 4856 29248 4862 29260
rect 4985 29257 4997 29260
rect 5031 29288 5043 29291
rect 5442 29288 5448 29300
rect 5031 29260 5448 29288
rect 5031 29257 5043 29260
rect 4985 29251 5043 29257
rect 5442 29248 5448 29260
rect 5500 29248 5506 29300
rect 8018 29248 8024 29300
rect 8076 29288 8082 29300
rect 8113 29291 8171 29297
rect 8113 29288 8125 29291
rect 8076 29260 8125 29288
rect 8076 29248 8082 29260
rect 8113 29257 8125 29260
rect 8159 29257 8171 29291
rect 8113 29251 8171 29257
rect 8294 29248 8300 29300
rect 8352 29288 8358 29300
rect 9677 29291 9735 29297
rect 9677 29288 9689 29291
rect 8352 29260 9689 29288
rect 8352 29248 8358 29260
rect 9677 29257 9689 29260
rect 9723 29257 9735 29291
rect 9677 29251 9735 29257
rect 2314 29220 2320 29232
rect 2227 29192 2320 29220
rect 2314 29180 2320 29192
rect 2372 29220 2378 29232
rect 5077 29223 5135 29229
rect 5077 29220 5089 29223
rect 2372 29192 5089 29220
rect 2372 29180 2378 29192
rect 5077 29189 5089 29192
rect 5123 29189 5135 29223
rect 6089 29223 6147 29229
rect 6089 29220 6101 29223
rect 5077 29183 5135 29189
rect 5552 29192 6101 29220
rect 4062 29152 4068 29164
rect 4023 29124 4068 29152
rect 4062 29112 4068 29124
rect 4120 29112 4126 29164
rect 5166 29112 5172 29164
rect 5224 29152 5230 29164
rect 5552 29161 5580 29192
rect 6089 29189 6101 29192
rect 6135 29189 6147 29223
rect 6089 29183 6147 29189
rect 7190 29180 7196 29232
rect 7248 29220 7254 29232
rect 8202 29220 8208 29232
rect 7248 29192 8208 29220
rect 7248 29180 7254 29192
rect 8202 29180 8208 29192
rect 8260 29180 8266 29232
rect 9490 29180 9496 29232
rect 9548 29220 9554 29232
rect 10781 29223 10839 29229
rect 10781 29220 10793 29223
rect 9548 29192 10793 29220
rect 9548 29180 9554 29192
rect 10781 29189 10793 29192
rect 10827 29189 10839 29223
rect 11793 29223 11851 29229
rect 11793 29220 11805 29223
rect 10781 29183 10839 29189
rect 11256 29192 11805 29220
rect 11256 29164 11284 29192
rect 11793 29189 11805 29192
rect 11839 29189 11851 29223
rect 11793 29183 11851 29189
rect 5537 29155 5595 29161
rect 5537 29152 5549 29155
rect 5224 29124 5549 29152
rect 5224 29112 5230 29124
rect 5537 29121 5549 29124
rect 5583 29121 5595 29155
rect 5537 29115 5595 29121
rect 5629 29155 5687 29161
rect 5629 29121 5641 29155
rect 5675 29152 5687 29155
rect 6270 29152 6276 29164
rect 5675 29124 6276 29152
rect 5675 29121 5687 29124
rect 5629 29115 5687 29121
rect 1443 29056 1992 29084
rect 4617 29087 4675 29093
rect 1443 29053 1455 29056
rect 1397 29047 1455 29053
rect 4617 29053 4629 29087
rect 4663 29084 4675 29087
rect 5644 29084 5672 29115
rect 6270 29112 6276 29124
rect 6328 29112 6334 29164
rect 11238 29152 11244 29164
rect 11199 29124 11244 29152
rect 11238 29112 11244 29124
rect 11296 29112 11302 29164
rect 11425 29155 11483 29161
rect 11425 29121 11437 29155
rect 11471 29152 11483 29155
rect 11606 29152 11612 29164
rect 11471 29124 11612 29152
rect 11471 29121 11483 29124
rect 11425 29115 11483 29121
rect 4663 29056 5672 29084
rect 4663 29053 4675 29056
rect 4617 29047 4675 29053
rect 7006 29044 7012 29096
rect 7064 29084 7070 29096
rect 7466 29084 7472 29096
rect 7064 29056 7472 29084
rect 7064 29044 7070 29056
rect 7466 29044 7472 29056
rect 7524 29044 7530 29096
rect 8297 29087 8355 29093
rect 8297 29053 8309 29087
rect 8343 29084 8355 29087
rect 8386 29084 8392 29096
rect 8343 29056 8392 29084
rect 8343 29053 8355 29056
rect 8297 29047 8355 29053
rect 8386 29044 8392 29056
rect 8444 29044 8450 29096
rect 11149 29087 11207 29093
rect 11149 29084 11161 29087
rect 10612 29056 11161 29084
rect 5445 29019 5503 29025
rect 5445 28985 5457 29019
rect 5491 29016 5503 29019
rect 7742 29016 7748 29028
rect 5491 28988 5580 29016
rect 7703 28988 7748 29016
rect 5491 28985 5503 28988
rect 5445 28979 5503 28985
rect 5552 28948 5580 28988
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 8570 29025 8576 29028
rect 8564 29016 8576 29025
rect 8531 28988 8576 29016
rect 8564 28979 8576 28988
rect 8570 28976 8576 28979
rect 8628 28976 8634 29028
rect 10042 29016 10048 29028
rect 9876 28988 10048 29016
rect 5902 28948 5908 28960
rect 5552 28920 5908 28948
rect 5902 28908 5908 28920
rect 5960 28908 5966 28960
rect 7466 28948 7472 28960
rect 7427 28920 7472 28948
rect 7466 28908 7472 28920
rect 7524 28908 7530 28960
rect 9876 28948 9904 28988
rect 10042 28976 10048 28988
rect 10100 28976 10106 29028
rect 10226 29016 10232 29028
rect 10187 28988 10232 29016
rect 10226 28976 10232 28988
rect 10284 28976 10290 29028
rect 10410 28976 10416 29028
rect 10468 29016 10474 29028
rect 10612 29025 10640 29056
rect 11149 29053 11161 29056
rect 11195 29053 11207 29087
rect 11149 29047 11207 29053
rect 10597 29019 10655 29025
rect 10597 29016 10609 29019
rect 10468 28988 10609 29016
rect 10468 28976 10474 28988
rect 10597 28985 10609 28988
rect 10643 28985 10655 29019
rect 11440 29016 11468 29115
rect 11606 29112 11612 29124
rect 11664 29112 11670 29164
rect 10597 28979 10655 28985
rect 11072 28988 11468 29016
rect 10778 28948 10784 28960
rect 9876 28920 10784 28948
rect 10778 28908 10784 28920
rect 10836 28908 10842 28960
rect 10870 28908 10876 28960
rect 10928 28948 10934 28960
rect 11072 28948 11100 28988
rect 10928 28920 11100 28948
rect 10928 28908 10934 28920
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 2774 28704 2780 28756
rect 2832 28744 2838 28756
rect 3053 28747 3111 28753
rect 3053 28744 3065 28747
rect 2832 28716 3065 28744
rect 2832 28704 2838 28716
rect 3053 28713 3065 28716
rect 3099 28713 3111 28747
rect 4522 28744 4528 28756
rect 4483 28716 4528 28744
rect 3053 28707 3111 28713
rect 3068 28676 3096 28707
rect 4522 28704 4528 28716
rect 4580 28704 4586 28756
rect 7466 28704 7472 28756
rect 7524 28744 7530 28756
rect 7653 28747 7711 28753
rect 7653 28744 7665 28747
rect 7524 28716 7665 28744
rect 7524 28704 7530 28716
rect 7653 28713 7665 28716
rect 7699 28744 7711 28747
rect 8570 28744 8576 28756
rect 7699 28716 8576 28744
rect 7699 28713 7711 28716
rect 7653 28707 7711 28713
rect 8570 28704 8576 28716
rect 8628 28744 8634 28756
rect 8665 28747 8723 28753
rect 8665 28744 8677 28747
rect 8628 28716 8677 28744
rect 8628 28704 8634 28716
rect 8665 28713 8677 28716
rect 8711 28744 8723 28747
rect 9401 28747 9459 28753
rect 9401 28744 9413 28747
rect 8711 28716 9413 28744
rect 8711 28713 8723 28716
rect 8665 28707 8723 28713
rect 9401 28713 9413 28716
rect 9447 28713 9459 28747
rect 10870 28744 10876 28756
rect 10831 28716 10876 28744
rect 9401 28707 9459 28713
rect 10870 28704 10876 28716
rect 10928 28704 10934 28756
rect 3510 28676 3516 28688
rect 3068 28648 3516 28676
rect 3510 28636 3516 28648
rect 3568 28676 3574 28688
rect 3568 28648 5111 28676
rect 3568 28636 3574 28648
rect 4798 28568 4804 28620
rect 4856 28608 4862 28620
rect 4893 28611 4951 28617
rect 4893 28608 4905 28611
rect 4856 28580 4905 28608
rect 4856 28568 4862 28580
rect 4893 28577 4905 28580
rect 4939 28577 4951 28611
rect 4893 28571 4951 28577
rect 4982 28540 4988 28552
rect 4943 28512 4988 28540
rect 4982 28500 4988 28512
rect 5040 28500 5046 28552
rect 5083 28549 5111 28648
rect 6178 28636 6184 28688
rect 6236 28676 6242 28688
rect 6518 28679 6576 28685
rect 6518 28676 6530 28679
rect 6236 28648 6530 28676
rect 6236 28636 6242 28648
rect 6518 28645 6530 28648
rect 6564 28645 6576 28679
rect 6518 28639 6576 28645
rect 11232 28679 11290 28685
rect 11232 28645 11244 28679
rect 11278 28676 11290 28679
rect 11422 28676 11428 28688
rect 11278 28648 11428 28676
rect 11278 28645 11290 28648
rect 11232 28639 11290 28645
rect 11422 28636 11428 28648
rect 11480 28676 11486 28688
rect 12342 28676 12348 28688
rect 11480 28648 12348 28676
rect 11480 28636 11486 28648
rect 12342 28636 12348 28648
rect 12400 28636 12406 28688
rect 5442 28568 5448 28620
rect 5500 28608 5506 28620
rect 6273 28611 6331 28617
rect 6273 28608 6285 28611
rect 5500 28580 6285 28608
rect 5500 28568 5506 28580
rect 6273 28577 6285 28580
rect 6319 28608 6331 28611
rect 6362 28608 6368 28620
rect 6319 28580 6368 28608
rect 6319 28577 6331 28580
rect 6273 28571 6331 28577
rect 6362 28568 6368 28580
rect 6420 28568 6426 28620
rect 8386 28608 8392 28620
rect 8299 28580 8392 28608
rect 8386 28568 8392 28580
rect 8444 28608 8450 28620
rect 10226 28608 10232 28620
rect 8444 28580 10232 28608
rect 8444 28568 8450 28580
rect 10226 28568 10232 28580
rect 10284 28608 10290 28620
rect 10965 28611 11023 28617
rect 10965 28608 10977 28611
rect 10284 28580 10977 28608
rect 10284 28568 10290 28580
rect 10965 28577 10977 28580
rect 11011 28608 11023 28611
rect 11054 28608 11060 28620
rect 11011 28580 11060 28608
rect 11011 28577 11023 28580
rect 10965 28571 11023 28577
rect 11054 28568 11060 28580
rect 11112 28568 11118 28620
rect 5077 28543 5135 28549
rect 5077 28509 5089 28543
rect 5123 28540 5135 28543
rect 5258 28540 5264 28552
rect 5123 28512 5264 28540
rect 5123 28509 5135 28512
rect 5077 28503 5135 28509
rect 5258 28500 5264 28512
rect 5316 28500 5322 28552
rect 5629 28475 5687 28481
rect 5629 28441 5641 28475
rect 5675 28472 5687 28475
rect 5994 28472 6000 28484
rect 5675 28444 6000 28472
rect 5675 28441 5687 28444
rect 5629 28435 5687 28441
rect 5994 28432 6000 28444
rect 6052 28432 6058 28484
rect 10321 28475 10379 28481
rect 10321 28441 10333 28475
rect 10367 28472 10379 28475
rect 10502 28472 10508 28484
rect 10367 28444 10508 28472
rect 10367 28441 10379 28444
rect 10321 28435 10379 28441
rect 10502 28432 10508 28444
rect 10560 28472 10566 28484
rect 10560 28444 10916 28472
rect 10560 28432 10566 28444
rect 5902 28404 5908 28416
rect 5863 28376 5908 28404
rect 5902 28364 5908 28376
rect 5960 28364 5966 28416
rect 10888 28404 10916 28444
rect 12345 28407 12403 28413
rect 12345 28404 12357 28407
rect 10888 28376 12357 28404
rect 12345 28373 12357 28376
rect 12391 28373 12403 28407
rect 12345 28367 12403 28373
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 2866 28200 2872 28212
rect 2827 28172 2872 28200
rect 2866 28160 2872 28172
rect 2924 28160 2930 28212
rect 3050 28200 3056 28212
rect 3011 28172 3056 28200
rect 3050 28160 3056 28172
rect 3108 28160 3114 28212
rect 4982 28200 4988 28212
rect 4943 28172 4988 28200
rect 4982 28160 4988 28172
rect 5040 28160 5046 28212
rect 5258 28200 5264 28212
rect 5219 28172 5264 28200
rect 5258 28160 5264 28172
rect 5316 28160 5322 28212
rect 5997 28203 6055 28209
rect 5997 28169 6009 28203
rect 6043 28200 6055 28203
rect 6178 28200 6184 28212
rect 6043 28172 6184 28200
rect 6043 28169 6055 28172
rect 5997 28163 6055 28169
rect 6178 28160 6184 28172
rect 6236 28160 6242 28212
rect 6362 28200 6368 28212
rect 6323 28172 6368 28200
rect 6362 28160 6368 28172
rect 6420 28160 6426 28212
rect 8386 28160 8392 28212
rect 8444 28200 8450 28212
rect 8846 28200 8852 28212
rect 8444 28172 8852 28200
rect 8444 28160 8450 28172
rect 8846 28160 8852 28172
rect 8904 28200 8910 28212
rect 9125 28203 9183 28209
rect 9125 28200 9137 28203
rect 8904 28172 9137 28200
rect 8904 28160 8910 28172
rect 9125 28169 9137 28172
rect 9171 28200 9183 28203
rect 9217 28203 9275 28209
rect 9217 28200 9229 28203
rect 9171 28172 9229 28200
rect 9171 28169 9183 28172
rect 9125 28163 9183 28169
rect 9217 28169 9229 28172
rect 9263 28169 9275 28203
rect 9398 28200 9404 28212
rect 9359 28172 9404 28200
rect 9217 28163 9275 28169
rect 9398 28160 9404 28172
rect 9456 28160 9462 28212
rect 11054 28200 11060 28212
rect 11015 28172 11060 28200
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11422 28200 11428 28212
rect 11383 28172 11428 28200
rect 11422 28160 11428 28172
rect 11480 28160 11486 28212
rect 3510 28024 3516 28076
rect 3568 28064 3574 28076
rect 3605 28067 3663 28073
rect 3605 28064 3617 28067
rect 3568 28036 3617 28064
rect 3568 28024 3574 28036
rect 3605 28033 3617 28036
rect 3651 28033 3663 28067
rect 3605 28027 3663 28033
rect 8481 28067 8539 28073
rect 8481 28033 8493 28067
rect 8527 28064 8539 28067
rect 8570 28064 8576 28076
rect 8527 28036 8576 28064
rect 8527 28033 8539 28036
rect 8481 28027 8539 28033
rect 8570 28024 8576 28036
rect 8628 28064 8634 28076
rect 8849 28067 8907 28073
rect 8849 28064 8861 28067
rect 8628 28036 8861 28064
rect 8628 28024 8634 28036
rect 8849 28033 8861 28036
rect 8895 28064 8907 28067
rect 9953 28067 10011 28073
rect 9953 28064 9965 28067
rect 8895 28036 9965 28064
rect 8895 28033 8907 28036
rect 8849 28027 8907 28033
rect 9953 28033 9965 28036
rect 9999 28033 10011 28067
rect 9953 28027 10011 28033
rect 2866 27956 2872 28008
rect 2924 27996 2930 28008
rect 3421 27999 3479 28005
rect 3421 27996 3433 27999
rect 2924 27968 3433 27996
rect 2924 27956 2930 27968
rect 3421 27965 3433 27968
rect 3467 27965 3479 27999
rect 3421 27959 3479 27965
rect 7377 27999 7435 28005
rect 7377 27965 7389 27999
rect 7423 27996 7435 27999
rect 7466 27996 7472 28008
rect 7423 27968 7472 27996
rect 7423 27965 7435 27968
rect 7377 27959 7435 27965
rect 7466 27956 7472 27968
rect 7524 27996 7530 28008
rect 8205 27999 8263 28005
rect 8205 27996 8217 27999
rect 7524 27968 8217 27996
rect 7524 27956 7530 27968
rect 8205 27965 8217 27968
rect 8251 27965 8263 27999
rect 8205 27959 8263 27965
rect 9125 27999 9183 28005
rect 9125 27965 9137 27999
rect 9171 27996 9183 27999
rect 9861 27999 9919 28005
rect 9861 27996 9873 27999
rect 9171 27968 9873 27996
rect 9171 27965 9183 27968
rect 9125 27959 9183 27965
rect 9861 27965 9873 27968
rect 9907 27965 9919 27999
rect 9861 27959 9919 27965
rect 2406 27888 2412 27940
rect 2464 27928 2470 27940
rect 2593 27931 2651 27937
rect 2593 27928 2605 27931
rect 2464 27900 2605 27928
rect 2464 27888 2470 27900
rect 2593 27897 2605 27900
rect 2639 27928 2651 27931
rect 3513 27931 3571 27937
rect 3513 27928 3525 27931
rect 2639 27900 3525 27928
rect 2639 27897 2651 27900
rect 2593 27891 2651 27897
rect 3513 27897 3525 27900
rect 3559 27897 3571 27931
rect 3513 27891 3571 27897
rect 4617 27931 4675 27937
rect 4617 27897 4629 27931
rect 4663 27928 4675 27931
rect 4798 27928 4804 27940
rect 4663 27900 4804 27928
rect 4663 27897 4675 27900
rect 4617 27891 4675 27897
rect 4798 27888 4804 27900
rect 4856 27928 4862 27940
rect 5810 27928 5816 27940
rect 4856 27900 5816 27928
rect 4856 27888 4862 27900
rect 5810 27888 5816 27900
rect 5868 27888 5874 27940
rect 7742 27928 7748 27940
rect 7655 27900 7748 27928
rect 7742 27888 7748 27900
rect 7800 27928 7806 27940
rect 7800 27900 8156 27928
rect 7800 27888 7806 27900
rect 7837 27863 7895 27869
rect 7837 27829 7849 27863
rect 7883 27860 7895 27863
rect 8018 27860 8024 27872
rect 7883 27832 8024 27860
rect 7883 27829 7895 27832
rect 7837 27823 7895 27829
rect 8018 27820 8024 27832
rect 8076 27820 8082 27872
rect 8128 27860 8156 27900
rect 9582 27888 9588 27940
rect 9640 27928 9646 27940
rect 9769 27931 9827 27937
rect 9769 27928 9781 27931
rect 9640 27900 9781 27928
rect 9640 27888 9646 27900
rect 9769 27897 9781 27900
rect 9815 27928 9827 27931
rect 11330 27928 11336 27940
rect 9815 27900 11336 27928
rect 9815 27897 9827 27900
rect 9769 27891 9827 27897
rect 11330 27888 11336 27900
rect 11388 27888 11394 27940
rect 8297 27863 8355 27869
rect 8297 27860 8309 27863
rect 8128 27832 8309 27860
rect 8297 27829 8309 27832
rect 8343 27860 8355 27863
rect 8570 27860 8576 27872
rect 8343 27832 8576 27860
rect 8343 27829 8355 27832
rect 8297 27823 8355 27829
rect 8570 27820 8576 27832
rect 8628 27820 8634 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 2406 27656 2412 27668
rect 2367 27628 2412 27656
rect 2406 27616 2412 27628
rect 2464 27616 2470 27668
rect 5258 27616 5264 27668
rect 5316 27656 5322 27668
rect 5445 27659 5503 27665
rect 5445 27656 5457 27659
rect 5316 27628 5457 27656
rect 5316 27616 5322 27628
rect 5445 27625 5457 27628
rect 5491 27625 5503 27659
rect 7558 27656 7564 27668
rect 7519 27628 7564 27656
rect 5445 27619 5503 27625
rect 7558 27616 7564 27628
rect 7616 27616 7622 27668
rect 8018 27656 8024 27668
rect 7979 27628 8024 27656
rect 8018 27616 8024 27628
rect 8076 27616 8082 27668
rect 10870 27656 10876 27668
rect 10831 27628 10876 27656
rect 10870 27616 10876 27628
rect 10928 27616 10934 27668
rect 2038 27548 2044 27600
rect 2096 27588 2102 27600
rect 2498 27588 2504 27600
rect 2096 27560 2504 27588
rect 2096 27548 2102 27560
rect 2498 27548 2504 27560
rect 2556 27588 2562 27600
rect 2869 27591 2927 27597
rect 2869 27588 2881 27591
rect 2556 27560 2881 27588
rect 2556 27548 2562 27560
rect 2869 27557 2881 27560
rect 2915 27588 2927 27591
rect 2958 27588 2964 27600
rect 2915 27560 2964 27588
rect 2915 27557 2927 27560
rect 2869 27551 2927 27557
rect 2958 27548 2964 27560
rect 3016 27548 3022 27600
rect 7926 27588 7932 27600
rect 7887 27560 7932 27588
rect 7926 27548 7932 27560
rect 7984 27548 7990 27600
rect 9493 27591 9551 27597
rect 9493 27557 9505 27591
rect 9539 27588 9551 27591
rect 9582 27588 9588 27600
rect 9539 27560 9588 27588
rect 9539 27557 9551 27560
rect 9493 27551 9551 27557
rect 9582 27548 9588 27560
rect 9640 27548 9646 27600
rect 11793 27591 11851 27597
rect 11793 27557 11805 27591
rect 11839 27588 11851 27591
rect 12130 27591 12188 27597
rect 12130 27588 12142 27591
rect 11839 27560 12142 27588
rect 11839 27557 11851 27560
rect 11793 27551 11851 27557
rect 12130 27557 12142 27560
rect 12176 27588 12188 27591
rect 12342 27588 12348 27600
rect 12176 27560 12348 27588
rect 12176 27557 12188 27560
rect 12130 27551 12188 27557
rect 12342 27548 12348 27560
rect 12400 27548 12406 27600
rect 2222 27480 2228 27532
rect 2280 27520 2286 27532
rect 2774 27520 2780 27532
rect 2280 27492 2780 27520
rect 2280 27480 2286 27492
rect 2774 27480 2780 27492
rect 2832 27520 2838 27532
rect 4338 27529 4344 27532
rect 4332 27520 4344 27529
rect 2832 27492 2877 27520
rect 3068 27492 4344 27520
rect 2832 27480 2838 27492
rect 3068 27461 3096 27492
rect 4332 27483 4344 27492
rect 4338 27480 4344 27483
rect 4396 27480 4402 27532
rect 10042 27520 10048 27532
rect 10003 27492 10048 27520
rect 10042 27480 10048 27492
rect 10100 27480 10106 27532
rect 11054 27480 11060 27532
rect 11112 27520 11118 27532
rect 11882 27520 11888 27532
rect 11112 27492 11888 27520
rect 11112 27480 11118 27492
rect 11882 27480 11888 27492
rect 11940 27480 11946 27532
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27421 3111 27455
rect 4062 27452 4068 27464
rect 4023 27424 4068 27452
rect 3053 27415 3111 27421
rect 4062 27412 4068 27424
rect 4120 27412 4126 27464
rect 8110 27452 8116 27464
rect 8071 27424 8116 27452
rect 8110 27412 8116 27424
rect 8168 27412 8174 27464
rect 8662 27412 8668 27464
rect 8720 27452 8726 27464
rect 8846 27452 8852 27464
rect 8720 27424 8852 27452
rect 8720 27412 8726 27424
rect 8846 27412 8852 27424
rect 8904 27452 8910 27464
rect 10137 27455 10195 27461
rect 10137 27452 10149 27455
rect 8904 27424 10149 27452
rect 8904 27412 8910 27424
rect 10137 27421 10149 27424
rect 10183 27421 10195 27455
rect 10137 27415 10195 27421
rect 10321 27455 10379 27461
rect 10321 27421 10333 27455
rect 10367 27452 10379 27455
rect 10870 27452 10876 27464
rect 10367 27424 10876 27452
rect 10367 27421 10379 27424
rect 10321 27415 10379 27421
rect 10870 27412 10876 27424
rect 10928 27412 10934 27464
rect 9125 27387 9183 27393
rect 9125 27353 9137 27387
rect 9171 27384 9183 27387
rect 9582 27384 9588 27396
rect 9171 27356 9588 27384
rect 9171 27353 9183 27356
rect 9125 27347 9183 27353
rect 9582 27344 9588 27356
rect 9640 27384 9646 27396
rect 9677 27387 9735 27393
rect 9677 27384 9689 27387
rect 9640 27356 9689 27384
rect 9640 27344 9646 27356
rect 9677 27353 9689 27356
rect 9723 27353 9735 27387
rect 9677 27347 9735 27353
rect 6917 27319 6975 27325
rect 6917 27285 6929 27319
rect 6963 27316 6975 27319
rect 7282 27316 7288 27328
rect 6963 27288 7288 27316
rect 6963 27285 6975 27288
rect 6917 27279 6975 27285
rect 7282 27276 7288 27288
rect 7340 27276 7346 27328
rect 13265 27319 13323 27325
rect 13265 27285 13277 27319
rect 13311 27316 13323 27319
rect 13446 27316 13452 27328
rect 13311 27288 13452 27316
rect 13311 27285 13323 27288
rect 13265 27279 13323 27285
rect 13446 27276 13452 27288
rect 13504 27276 13510 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 1765 27115 1823 27121
rect 1765 27081 1777 27115
rect 1811 27112 1823 27115
rect 3973 27115 4031 27121
rect 3973 27112 3985 27115
rect 1811 27084 3985 27112
rect 1811 27081 1823 27084
rect 1765 27075 1823 27081
rect 3973 27081 3985 27084
rect 4019 27112 4031 27115
rect 4338 27112 4344 27124
rect 4019 27084 4344 27112
rect 4019 27081 4031 27084
rect 3973 27075 4031 27081
rect 4338 27072 4344 27084
rect 4396 27112 4402 27124
rect 4893 27115 4951 27121
rect 4893 27112 4905 27115
rect 4396 27084 4905 27112
rect 4396 27072 4402 27084
rect 4893 27081 4905 27084
rect 4939 27081 4951 27115
rect 4893 27075 4951 27081
rect 8018 27072 8024 27124
rect 8076 27112 8082 27124
rect 8205 27115 8263 27121
rect 8205 27112 8217 27115
rect 8076 27084 8217 27112
rect 8076 27072 8082 27084
rect 8205 27081 8217 27084
rect 8251 27081 8263 27115
rect 8205 27075 8263 27081
rect 10134 27072 10140 27124
rect 10192 27112 10198 27124
rect 10229 27115 10287 27121
rect 10229 27112 10241 27115
rect 10192 27084 10241 27112
rect 10192 27072 10198 27084
rect 10229 27081 10241 27084
rect 10275 27081 10287 27115
rect 10229 27075 10287 27081
rect 2133 27047 2191 27053
rect 2133 27013 2145 27047
rect 2179 27044 2191 27047
rect 2222 27044 2228 27056
rect 2179 27016 2228 27044
rect 2179 27013 2191 27016
rect 2133 27007 2191 27013
rect 2222 27004 2228 27016
rect 2280 27004 2286 27056
rect 2498 27044 2504 27056
rect 2459 27016 2504 27044
rect 2498 27004 2504 27016
rect 2556 27004 2562 27056
rect 4062 27004 4068 27056
rect 4120 27044 4126 27056
rect 4617 27047 4675 27053
rect 4617 27044 4629 27047
rect 4120 27016 4629 27044
rect 4120 27004 4126 27016
rect 4617 27013 4629 27016
rect 4663 27044 4675 27047
rect 5442 27044 5448 27056
rect 4663 27016 5448 27044
rect 4663 27013 4675 27016
rect 4617 27007 4675 27013
rect 5442 27004 5448 27016
rect 5500 27004 5506 27056
rect 6178 27004 6184 27056
rect 6236 27044 6242 27056
rect 6273 27047 6331 27053
rect 6273 27044 6285 27047
rect 6236 27016 6285 27044
rect 6236 27004 6242 27016
rect 6273 27013 6285 27016
rect 6319 27044 6331 27047
rect 7929 27047 7987 27053
rect 6319 27016 7512 27044
rect 6319 27013 6331 27016
rect 6273 27007 6331 27013
rect 2593 26911 2651 26917
rect 2593 26877 2605 26911
rect 2639 26908 2651 26911
rect 2682 26908 2688 26920
rect 2639 26880 2688 26908
rect 2639 26877 2651 26880
rect 2593 26871 2651 26877
rect 2682 26868 2688 26880
rect 2740 26908 2746 26920
rect 4080 26908 4108 27004
rect 7282 26976 7288 26988
rect 7243 26948 7288 26976
rect 7282 26936 7288 26948
rect 7340 26936 7346 26988
rect 7484 26985 7512 27016
rect 7929 27013 7941 27047
rect 7975 27044 7987 27047
rect 8110 27044 8116 27056
rect 7975 27016 8116 27044
rect 7975 27013 7987 27016
rect 7929 27007 7987 27013
rect 8110 27004 8116 27016
rect 8168 27004 8174 27056
rect 11882 27004 11888 27056
rect 11940 27044 11946 27056
rect 13449 27047 13507 27053
rect 13449 27044 13461 27047
rect 11940 27016 13461 27044
rect 11940 27004 11946 27016
rect 13449 27013 13461 27016
rect 13495 27013 13507 27047
rect 13449 27007 13507 27013
rect 7469 26979 7527 26985
rect 7469 26945 7481 26979
rect 7515 26976 7527 26979
rect 7650 26976 7656 26988
rect 7515 26948 7656 26976
rect 7515 26945 7527 26948
rect 7469 26939 7527 26945
rect 7650 26936 7656 26948
rect 7708 26936 7714 26988
rect 8757 26979 8815 26985
rect 8757 26945 8769 26979
rect 8803 26976 8815 26979
rect 9490 26976 9496 26988
rect 8803 26948 9496 26976
rect 8803 26945 8815 26948
rect 8757 26939 8815 26945
rect 9490 26936 9496 26948
rect 9548 26976 9554 26988
rect 9677 26979 9735 26985
rect 9677 26976 9689 26979
rect 9548 26948 9689 26976
rect 9548 26936 9554 26948
rect 9677 26945 9689 26948
rect 9723 26945 9735 26979
rect 9858 26976 9864 26988
rect 9819 26948 9864 26976
rect 9677 26939 9735 26945
rect 9858 26936 9864 26948
rect 9916 26936 9922 26988
rect 10870 26936 10876 26988
rect 10928 26976 10934 26988
rect 11238 26976 11244 26988
rect 10928 26948 11244 26976
rect 10928 26936 10934 26948
rect 11238 26936 11244 26948
rect 11296 26976 11302 26988
rect 11333 26979 11391 26985
rect 11333 26976 11345 26979
rect 11296 26948 11345 26976
rect 11296 26936 11302 26948
rect 11333 26945 11345 26948
rect 11379 26945 11391 26979
rect 12986 26976 12992 26988
rect 12947 26948 12992 26976
rect 11333 26939 11391 26945
rect 12986 26936 12992 26948
rect 13044 26936 13050 26988
rect 9582 26908 9588 26920
rect 2740 26880 4108 26908
rect 9543 26880 9588 26908
rect 2740 26868 2746 26880
rect 9582 26868 9588 26880
rect 9640 26868 9646 26920
rect 10778 26868 10784 26920
rect 10836 26908 10842 26920
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 10836 26880 12909 26908
rect 10836 26868 10842 26880
rect 2860 26843 2918 26849
rect 2860 26809 2872 26843
rect 2906 26840 2918 26843
rect 2958 26840 2964 26852
rect 2906 26812 2964 26840
rect 2906 26809 2918 26812
rect 2860 26803 2918 26809
rect 2958 26800 2964 26812
rect 3016 26800 3022 26852
rect 6641 26843 6699 26849
rect 6641 26809 6653 26843
rect 6687 26840 6699 26843
rect 11241 26843 11299 26849
rect 11241 26840 11253 26843
rect 6687 26812 7236 26840
rect 6687 26809 6699 26812
rect 6641 26803 6699 26809
rect 6822 26772 6828 26784
rect 6783 26744 6828 26772
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 7208 26781 7236 26812
rect 10612 26812 11253 26840
rect 7193 26775 7251 26781
rect 7193 26741 7205 26775
rect 7239 26772 7251 26775
rect 7374 26772 7380 26784
rect 7239 26744 7380 26772
rect 7239 26741 7251 26744
rect 7193 26735 7251 26741
rect 7374 26732 7380 26744
rect 7432 26772 7438 26784
rect 8478 26772 8484 26784
rect 7432 26744 8484 26772
rect 7432 26732 7438 26744
rect 8478 26732 8484 26744
rect 8536 26732 8542 26784
rect 8846 26732 8852 26784
rect 8904 26772 8910 26784
rect 9033 26775 9091 26781
rect 9033 26772 9045 26775
rect 8904 26744 9045 26772
rect 8904 26732 8910 26744
rect 9033 26741 9045 26744
rect 9079 26741 9091 26775
rect 9033 26735 9091 26741
rect 9217 26775 9275 26781
rect 9217 26741 9229 26775
rect 9263 26772 9275 26775
rect 9306 26772 9312 26784
rect 9263 26744 9312 26772
rect 9263 26741 9275 26744
rect 9217 26735 9275 26741
rect 9306 26732 9312 26744
rect 9364 26732 9370 26784
rect 10410 26732 10416 26784
rect 10468 26772 10474 26784
rect 10612 26781 10640 26812
rect 11241 26809 11253 26812
rect 11287 26840 11299 26843
rect 11330 26840 11336 26852
rect 11287 26812 11336 26840
rect 11287 26809 11299 26812
rect 11241 26803 11299 26809
rect 11330 26800 11336 26812
rect 11388 26800 11394 26852
rect 11532 26784 11560 26880
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 12897 26871 12955 26877
rect 12250 26840 12256 26852
rect 12211 26812 12256 26840
rect 12250 26800 12256 26812
rect 12308 26800 12314 26852
rect 12802 26840 12808 26852
rect 12763 26812 12808 26840
rect 12802 26800 12808 26812
rect 12860 26800 12866 26852
rect 10597 26775 10655 26781
rect 10597 26772 10609 26775
rect 10468 26744 10609 26772
rect 10468 26732 10474 26744
rect 10597 26741 10609 26744
rect 10643 26741 10655 26775
rect 10778 26772 10784 26784
rect 10739 26744 10784 26772
rect 10597 26735 10655 26741
rect 10778 26732 10784 26744
rect 10836 26732 10842 26784
rect 10870 26732 10876 26784
rect 10928 26772 10934 26784
rect 11149 26775 11207 26781
rect 11149 26772 11161 26775
rect 10928 26744 11161 26772
rect 10928 26732 10934 26744
rect 11149 26741 11161 26744
rect 11195 26741 11207 26775
rect 11149 26735 11207 26741
rect 11514 26732 11520 26784
rect 11572 26772 11578 26784
rect 11793 26775 11851 26781
rect 11793 26772 11805 26775
rect 11572 26744 11805 26772
rect 11572 26732 11578 26744
rect 11793 26741 11805 26744
rect 11839 26741 11851 26775
rect 11793 26735 11851 26741
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 12492 26744 12537 26772
rect 12492 26732 12498 26744
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 2222 26528 2228 26580
rect 2280 26568 2286 26580
rect 2682 26568 2688 26580
rect 2280 26540 2688 26568
rect 2280 26528 2286 26540
rect 2682 26528 2688 26540
rect 2740 26528 2746 26580
rect 2958 26568 2964 26580
rect 2919 26540 2964 26568
rect 2958 26528 2964 26540
rect 3016 26528 3022 26580
rect 5813 26571 5871 26577
rect 5813 26537 5825 26571
rect 5859 26568 5871 26571
rect 6365 26571 6423 26577
rect 6365 26568 6377 26571
rect 5859 26540 6377 26568
rect 5859 26537 5871 26540
rect 5813 26531 5871 26537
rect 6365 26537 6377 26540
rect 6411 26568 6423 26571
rect 6822 26568 6828 26580
rect 6411 26540 6828 26568
rect 6411 26537 6423 26540
rect 6365 26531 6423 26537
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 7926 26568 7932 26580
rect 7887 26540 7932 26568
rect 7926 26528 7932 26540
rect 7984 26528 7990 26580
rect 9953 26571 10011 26577
rect 9953 26537 9965 26571
rect 9999 26568 10011 26571
rect 10870 26568 10876 26580
rect 9999 26540 10876 26568
rect 9999 26537 10011 26540
rect 9953 26531 10011 26537
rect 10870 26528 10876 26540
rect 10928 26528 10934 26580
rect 12342 26568 12348 26580
rect 12303 26540 12348 26568
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 11238 26509 11244 26512
rect 10505 26503 10563 26509
rect 10505 26469 10517 26503
rect 10551 26500 10563 26503
rect 11232 26500 11244 26509
rect 10551 26472 11244 26500
rect 10551 26469 10563 26472
rect 10505 26463 10563 26469
rect 11232 26463 11244 26472
rect 11296 26500 11302 26512
rect 12986 26500 12992 26512
rect 11296 26472 12992 26500
rect 11238 26460 11244 26463
rect 11296 26460 11302 26472
rect 12986 26460 12992 26472
rect 13044 26460 13050 26512
rect 5445 26435 5503 26441
rect 5445 26401 5457 26435
rect 5491 26432 5503 26435
rect 6273 26435 6331 26441
rect 6273 26432 6285 26435
rect 5491 26404 6285 26432
rect 5491 26401 5503 26404
rect 5445 26395 5503 26401
rect 6273 26401 6285 26404
rect 6319 26432 6331 26435
rect 6822 26432 6828 26444
rect 6319 26404 6828 26432
rect 6319 26401 6331 26404
rect 6273 26395 6331 26401
rect 6822 26392 6828 26404
rect 6880 26392 6886 26444
rect 10870 26392 10876 26444
rect 10928 26432 10934 26444
rect 12342 26432 12348 26444
rect 10928 26404 12348 26432
rect 10928 26392 10934 26404
rect 12342 26392 12348 26404
rect 12400 26392 12406 26444
rect 5994 26324 6000 26376
rect 6052 26364 6058 26376
rect 6457 26367 6515 26373
rect 6457 26364 6469 26367
rect 6052 26336 6469 26364
rect 6052 26324 6058 26336
rect 6457 26333 6469 26336
rect 6503 26333 6515 26367
rect 6457 26327 6515 26333
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26364 7067 26367
rect 7190 26364 7196 26376
rect 7055 26336 7196 26364
rect 7055 26333 7067 26336
rect 7009 26327 7067 26333
rect 7190 26324 7196 26336
rect 7248 26364 7254 26376
rect 7469 26367 7527 26373
rect 7469 26364 7481 26367
rect 7248 26336 7481 26364
rect 7248 26324 7254 26336
rect 7469 26333 7481 26336
rect 7515 26333 7527 26367
rect 7469 26327 7527 26333
rect 10965 26367 11023 26373
rect 10965 26333 10977 26367
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 5902 26296 5908 26308
rect 5863 26268 5908 26296
rect 5902 26256 5908 26268
rect 5960 26256 5966 26308
rect 9309 26299 9367 26305
rect 9309 26265 9321 26299
rect 9355 26296 9367 26299
rect 9355 26268 9628 26296
rect 9355 26265 9367 26268
rect 9309 26259 9367 26265
rect 4617 26231 4675 26237
rect 4617 26197 4629 26231
rect 4663 26228 4675 26231
rect 4982 26228 4988 26240
rect 4663 26200 4988 26228
rect 4663 26197 4675 26200
rect 4617 26191 4675 26197
rect 4982 26188 4988 26200
rect 5040 26228 5046 26240
rect 6730 26228 6736 26240
rect 5040 26200 6736 26228
rect 5040 26188 5046 26200
rect 6730 26188 6736 26200
rect 6788 26188 6794 26240
rect 8662 26228 8668 26240
rect 8623 26200 8668 26228
rect 8662 26188 8668 26200
rect 8720 26188 8726 26240
rect 9600 26228 9628 26268
rect 9858 26228 9864 26240
rect 9600 26200 9864 26228
rect 9858 26188 9864 26200
rect 9916 26188 9922 26240
rect 10980 26228 11008 26327
rect 11146 26228 11152 26240
rect 10980 26200 11152 26228
rect 11146 26188 11152 26200
rect 11204 26188 11210 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 1578 26024 1584 26036
rect 1539 25996 1584 26024
rect 1578 25984 1584 25996
rect 1636 25984 1642 26036
rect 6178 26024 6184 26036
rect 6139 25996 6184 26024
rect 6178 25984 6184 25996
rect 6236 25984 6242 26036
rect 6822 26024 6828 26036
rect 6783 25996 6828 26024
rect 6822 25984 6828 25996
rect 6880 25984 6886 26036
rect 9858 25984 9864 26036
rect 9916 26024 9922 26036
rect 10045 26027 10103 26033
rect 10045 26024 10057 26027
rect 9916 25996 10057 26024
rect 9916 25984 9922 25996
rect 10045 25993 10057 25996
rect 10091 26024 10103 26027
rect 10091 25996 10732 26024
rect 10091 25993 10103 25996
rect 10045 25987 10103 25993
rect 5077 25891 5135 25897
rect 5077 25888 5089 25891
rect 5000 25860 5089 25888
rect 1397 25823 1455 25829
rect 1397 25789 1409 25823
rect 1443 25820 1455 25823
rect 1443 25792 1992 25820
rect 1443 25789 1455 25792
rect 1397 25783 1455 25789
rect 1964 25696 1992 25792
rect 4338 25780 4344 25832
rect 4396 25820 4402 25832
rect 4893 25823 4951 25829
rect 4893 25820 4905 25823
rect 4396 25792 4905 25820
rect 4396 25780 4402 25792
rect 4893 25789 4905 25792
rect 4939 25789 4951 25823
rect 4893 25783 4951 25789
rect 5000 25752 5028 25860
rect 5077 25857 5089 25860
rect 5123 25857 5135 25891
rect 6196 25888 6224 25984
rect 8570 25956 8576 25968
rect 8531 25928 8576 25956
rect 8570 25916 8576 25928
rect 8628 25916 8634 25968
rect 10137 25959 10195 25965
rect 10137 25925 10149 25959
rect 10183 25925 10195 25959
rect 10137 25919 10195 25925
rect 7377 25891 7435 25897
rect 7377 25888 7389 25891
rect 6196 25860 7389 25888
rect 5077 25851 5135 25857
rect 7377 25857 7389 25860
rect 7423 25857 7435 25891
rect 7377 25851 7435 25857
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25888 8539 25891
rect 9217 25891 9275 25897
rect 9217 25888 9229 25891
rect 8527 25860 9229 25888
rect 8527 25857 8539 25860
rect 8481 25851 8539 25857
rect 9217 25857 9229 25860
rect 9263 25888 9275 25891
rect 9398 25888 9404 25900
rect 9263 25860 9404 25888
rect 9263 25857 9275 25860
rect 9217 25851 9275 25857
rect 9398 25848 9404 25860
rect 9456 25848 9462 25900
rect 7190 25820 7196 25832
rect 7151 25792 7196 25820
rect 7190 25780 7196 25792
rect 7248 25780 7254 25832
rect 8662 25780 8668 25832
rect 8720 25820 8726 25832
rect 8941 25823 8999 25829
rect 8941 25820 8953 25823
rect 8720 25792 8953 25820
rect 8720 25780 8726 25792
rect 8941 25789 8953 25792
rect 8987 25820 8999 25823
rect 10152 25820 10180 25919
rect 10594 25888 10600 25900
rect 10555 25860 10600 25888
rect 10594 25848 10600 25860
rect 10652 25848 10658 25900
rect 10704 25897 10732 25996
rect 11054 25984 11060 26036
rect 11112 26024 11118 26036
rect 11149 26027 11207 26033
rect 11149 26024 11161 26027
rect 11112 25996 11161 26024
rect 11112 25984 11118 25996
rect 11149 25993 11161 25996
rect 11195 25993 11207 26027
rect 11149 25987 11207 25993
rect 11238 25984 11244 26036
rect 11296 26024 11302 26036
rect 11517 26027 11575 26033
rect 11517 26024 11529 26027
rect 11296 25996 11529 26024
rect 11296 25984 11302 25996
rect 11517 25993 11529 25996
rect 11563 25993 11575 26027
rect 11517 25987 11575 25993
rect 10689 25891 10747 25897
rect 10689 25857 10701 25891
rect 10735 25888 10747 25891
rect 10870 25888 10876 25900
rect 10735 25860 10876 25888
rect 10735 25857 10747 25860
rect 10689 25851 10747 25857
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 8987 25792 10180 25820
rect 10505 25823 10563 25829
rect 8987 25789 8999 25792
rect 8941 25783 8999 25789
rect 10505 25789 10517 25823
rect 10551 25820 10563 25823
rect 10778 25820 10784 25832
rect 10551 25792 10784 25820
rect 10551 25789 10563 25792
rect 10505 25783 10563 25789
rect 4080 25724 5028 25752
rect 9033 25755 9091 25761
rect 4080 25696 4108 25724
rect 9033 25721 9045 25755
rect 9079 25752 9091 25755
rect 9306 25752 9312 25764
rect 9079 25724 9312 25752
rect 9079 25721 9091 25724
rect 9033 25715 9091 25721
rect 9306 25712 9312 25724
rect 9364 25712 9370 25764
rect 9677 25755 9735 25761
rect 9677 25721 9689 25755
rect 9723 25752 9735 25755
rect 10520 25752 10548 25783
rect 10778 25780 10784 25792
rect 10836 25780 10842 25832
rect 9723 25724 10548 25752
rect 9723 25721 9735 25724
rect 9677 25715 9735 25721
rect 1946 25684 1952 25696
rect 1907 25656 1952 25684
rect 1946 25644 1952 25656
rect 2004 25644 2010 25696
rect 4062 25684 4068 25696
rect 4023 25656 4068 25684
rect 4062 25644 4068 25656
rect 4120 25644 4126 25696
rect 4338 25684 4344 25696
rect 4299 25656 4344 25684
rect 4338 25644 4344 25656
rect 4396 25644 4402 25696
rect 4522 25684 4528 25696
rect 4483 25656 4528 25684
rect 4522 25644 4528 25656
rect 4580 25644 4586 25696
rect 4982 25684 4988 25696
rect 4943 25656 4988 25684
rect 4982 25644 4988 25656
rect 5040 25644 5046 25696
rect 5902 25684 5908 25696
rect 5863 25656 5908 25684
rect 5902 25644 5908 25656
rect 5960 25644 5966 25696
rect 6641 25687 6699 25693
rect 6641 25653 6653 25687
rect 6687 25684 6699 25687
rect 7282 25684 7288 25696
rect 6687 25656 7288 25684
rect 6687 25653 6699 25656
rect 6641 25647 6699 25653
rect 7282 25644 7288 25656
rect 7340 25644 7346 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 1946 25440 1952 25492
rect 2004 25480 2010 25492
rect 2317 25483 2375 25489
rect 2317 25480 2329 25483
rect 2004 25452 2329 25480
rect 2004 25440 2010 25452
rect 2317 25449 2329 25452
rect 2363 25449 2375 25483
rect 2317 25443 2375 25449
rect 4246 25440 4252 25492
rect 4304 25480 4310 25492
rect 4982 25480 4988 25492
rect 4304 25452 4988 25480
rect 4304 25440 4310 25452
rect 4982 25440 4988 25452
rect 5040 25440 5046 25492
rect 5902 25440 5908 25492
rect 5960 25480 5966 25492
rect 6549 25483 6607 25489
rect 6549 25480 6561 25483
rect 5960 25452 6561 25480
rect 5960 25440 5966 25452
rect 6549 25449 6561 25452
rect 6595 25449 6607 25483
rect 6549 25443 6607 25449
rect 8665 25483 8723 25489
rect 8665 25449 8677 25483
rect 8711 25480 8723 25483
rect 9306 25480 9312 25492
rect 8711 25452 9312 25480
rect 8711 25449 8723 25452
rect 8665 25443 8723 25449
rect 9306 25440 9312 25452
rect 9364 25440 9370 25492
rect 10229 25483 10287 25489
rect 10229 25449 10241 25483
rect 10275 25480 10287 25483
rect 10594 25480 10600 25492
rect 10275 25452 10600 25480
rect 10275 25449 10287 25452
rect 10229 25443 10287 25449
rect 10594 25440 10600 25452
rect 10652 25440 10658 25492
rect 2685 25415 2743 25421
rect 2685 25381 2697 25415
rect 2731 25412 2743 25415
rect 2774 25412 2780 25424
rect 2731 25384 2780 25412
rect 2731 25381 2743 25384
rect 2685 25375 2743 25381
rect 2774 25372 2780 25384
rect 2832 25372 2838 25424
rect 5436 25415 5494 25421
rect 5436 25381 5448 25415
rect 5482 25412 5494 25415
rect 6178 25412 6184 25424
rect 5482 25384 6184 25412
rect 5482 25381 5494 25384
rect 5436 25375 5494 25381
rect 6178 25372 6184 25384
rect 6236 25372 6242 25424
rect 2682 25236 2688 25288
rect 2740 25276 2746 25288
rect 2777 25279 2835 25285
rect 2777 25276 2789 25279
rect 2740 25248 2789 25276
rect 2740 25236 2746 25248
rect 2777 25245 2789 25248
rect 2823 25245 2835 25279
rect 2958 25276 2964 25288
rect 2919 25248 2964 25276
rect 2777 25239 2835 25245
rect 2958 25236 2964 25248
rect 3016 25236 3022 25288
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25276 4215 25279
rect 4617 25279 4675 25285
rect 4617 25276 4629 25279
rect 4203 25248 4629 25276
rect 4203 25245 4215 25248
rect 4157 25239 4215 25245
rect 4617 25245 4629 25248
rect 4663 25276 4675 25279
rect 4982 25276 4988 25288
rect 4663 25248 4988 25276
rect 4663 25245 4675 25248
rect 4617 25239 4675 25245
rect 4982 25236 4988 25248
rect 5040 25236 5046 25288
rect 5169 25279 5227 25285
rect 5169 25245 5181 25279
rect 5215 25245 5227 25279
rect 5169 25239 5227 25245
rect 2590 25168 2596 25220
rect 2648 25208 2654 25220
rect 2976 25208 3004 25236
rect 2648 25180 3004 25208
rect 2648 25168 2654 25180
rect 2225 25143 2283 25149
rect 2225 25109 2237 25143
rect 2271 25140 2283 25143
rect 2406 25140 2412 25152
rect 2271 25112 2412 25140
rect 2271 25109 2283 25112
rect 2225 25103 2283 25109
rect 2406 25100 2412 25112
rect 2464 25100 2470 25152
rect 5184 25140 5212 25239
rect 5442 25140 5448 25152
rect 5184 25112 5448 25140
rect 5442 25100 5448 25112
rect 5500 25100 5506 25152
rect 7926 25140 7932 25152
rect 7887 25112 7932 25140
rect 7926 25100 7932 25112
rect 7984 25100 7990 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 4062 24936 4068 24948
rect 4023 24908 4068 24936
rect 4062 24896 4068 24908
rect 4120 24896 4126 24948
rect 6089 24939 6147 24945
rect 6089 24905 6101 24939
rect 6135 24936 6147 24939
rect 6178 24936 6184 24948
rect 6135 24908 6184 24936
rect 6135 24905 6147 24908
rect 6089 24899 6147 24905
rect 6178 24896 6184 24908
rect 6236 24896 6242 24948
rect 4080 24868 4108 24896
rect 4614 24868 4620 24880
rect 4080 24840 4620 24868
rect 4614 24828 4620 24840
rect 4672 24868 4678 24880
rect 4672 24840 5212 24868
rect 4672 24828 4678 24840
rect 4525 24803 4583 24809
rect 4525 24769 4537 24803
rect 4571 24800 4583 24803
rect 5074 24800 5080 24812
rect 4571 24772 5080 24800
rect 4571 24769 4583 24772
rect 4525 24763 4583 24769
rect 5074 24760 5080 24772
rect 5132 24760 5138 24812
rect 5184 24809 5212 24840
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24769 5227 24803
rect 5169 24763 5227 24769
rect 2041 24735 2099 24741
rect 2041 24701 2053 24735
rect 2087 24732 2099 24735
rect 2133 24735 2191 24741
rect 2133 24732 2145 24735
rect 2087 24704 2145 24732
rect 2087 24701 2099 24704
rect 2041 24695 2099 24701
rect 2133 24701 2145 24704
rect 2179 24732 2191 24735
rect 2222 24732 2228 24744
rect 2179 24704 2228 24732
rect 2179 24701 2191 24704
rect 2133 24695 2191 24701
rect 2222 24692 2228 24704
rect 2280 24692 2286 24744
rect 2406 24741 2412 24744
rect 2400 24732 2412 24741
rect 2367 24704 2412 24732
rect 2400 24695 2412 24704
rect 2406 24692 2412 24695
rect 2464 24692 2470 24744
rect 4982 24732 4988 24744
rect 4943 24704 4988 24732
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 5442 24692 5448 24744
rect 5500 24732 5506 24744
rect 5721 24735 5779 24741
rect 5721 24732 5733 24735
rect 5500 24704 5733 24732
rect 5500 24692 5506 24704
rect 5721 24701 5733 24704
rect 5767 24732 5779 24735
rect 7745 24735 7803 24741
rect 7745 24732 7757 24735
rect 5767 24704 7757 24732
rect 5767 24701 5779 24704
rect 5721 24695 5779 24701
rect 7745 24701 7757 24704
rect 7791 24732 7803 24735
rect 7837 24735 7895 24741
rect 7837 24732 7849 24735
rect 7791 24704 7849 24732
rect 7791 24701 7803 24704
rect 7745 24695 7803 24701
rect 7837 24701 7849 24704
rect 7883 24701 7895 24735
rect 7837 24695 7895 24701
rect 2682 24664 2688 24676
rect 2516 24636 2688 24664
rect 1673 24599 1731 24605
rect 1673 24565 1685 24599
rect 1719 24596 1731 24599
rect 2516 24596 2544 24636
rect 2682 24624 2688 24636
rect 2740 24624 2746 24676
rect 7852 24664 7880 24695
rect 7926 24692 7932 24744
rect 7984 24732 7990 24744
rect 8093 24735 8151 24741
rect 8093 24732 8105 24735
rect 7984 24704 8105 24732
rect 7984 24692 7990 24704
rect 8093 24701 8105 24704
rect 8139 24701 8151 24735
rect 8093 24695 8151 24701
rect 8662 24664 8668 24676
rect 7852 24636 8668 24664
rect 8662 24624 8668 24636
rect 8720 24624 8726 24676
rect 10226 24624 10232 24676
rect 10284 24664 10290 24676
rect 10870 24664 10876 24676
rect 10284 24636 10876 24664
rect 10284 24624 10290 24636
rect 10870 24624 10876 24636
rect 10928 24624 10934 24676
rect 1719 24568 2544 24596
rect 1719 24565 1731 24568
rect 1673 24559 1731 24565
rect 2590 24556 2596 24608
rect 2648 24596 2654 24608
rect 3513 24599 3571 24605
rect 3513 24596 3525 24599
rect 2648 24568 3525 24596
rect 2648 24556 2654 24568
rect 3513 24565 3525 24568
rect 3559 24565 3571 24599
rect 3513 24559 3571 24565
rect 4617 24599 4675 24605
rect 4617 24565 4629 24599
rect 4663 24596 4675 24599
rect 4798 24596 4804 24608
rect 4663 24568 4804 24596
rect 4663 24565 4675 24568
rect 4617 24559 4675 24565
rect 4798 24556 4804 24568
rect 4856 24556 4862 24608
rect 8018 24556 8024 24608
rect 8076 24596 8082 24608
rect 9217 24599 9275 24605
rect 9217 24596 9229 24599
rect 8076 24568 9229 24596
rect 8076 24556 8082 24568
rect 9217 24565 9229 24568
rect 9263 24565 9275 24599
rect 9217 24559 9275 24565
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 2409 24395 2467 24401
rect 2409 24361 2421 24395
rect 2455 24392 2467 24395
rect 2590 24392 2596 24404
rect 2455 24364 2596 24392
rect 2455 24361 2467 24364
rect 2409 24355 2467 24361
rect 2590 24352 2596 24364
rect 2648 24352 2654 24404
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 4065 24395 4123 24401
rect 4065 24392 4077 24395
rect 2832 24364 4077 24392
rect 2832 24352 2838 24364
rect 4065 24361 4077 24364
rect 4111 24361 4123 24395
rect 4522 24392 4528 24404
rect 4483 24364 4528 24392
rect 4065 24355 4123 24361
rect 4522 24352 4528 24364
rect 4580 24352 4586 24404
rect 7285 24395 7343 24401
rect 7285 24361 7297 24395
rect 7331 24392 7343 24395
rect 7837 24395 7895 24401
rect 7837 24392 7849 24395
rect 7331 24364 7849 24392
rect 7331 24361 7343 24364
rect 7285 24355 7343 24361
rect 7837 24361 7849 24364
rect 7883 24392 7895 24395
rect 9677 24395 9735 24401
rect 9677 24392 9689 24395
rect 7883 24364 9689 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 9677 24361 9689 24364
rect 9723 24361 9735 24395
rect 9677 24355 9735 24361
rect 10137 24395 10195 24401
rect 10137 24361 10149 24395
rect 10183 24392 10195 24395
rect 10226 24392 10232 24404
rect 10183 24364 10232 24392
rect 10183 24361 10195 24364
rect 10137 24355 10195 24361
rect 5534 24284 5540 24336
rect 5592 24324 5598 24336
rect 7742 24324 7748 24336
rect 5592 24296 7748 24324
rect 5592 24284 5598 24296
rect 7742 24284 7748 24296
rect 7800 24284 7806 24336
rect 9306 24284 9312 24336
rect 9364 24324 9370 24336
rect 10152 24324 10180 24355
rect 10226 24352 10232 24364
rect 10284 24352 10290 24404
rect 9364 24296 10180 24324
rect 9364 24284 9370 24296
rect 4433 24259 4491 24265
rect 4433 24225 4445 24259
rect 4479 24256 4491 24259
rect 4798 24256 4804 24268
rect 4479 24228 4804 24256
rect 4479 24225 4491 24228
rect 4433 24219 4491 24225
rect 4798 24216 4804 24228
rect 4856 24216 4862 24268
rect 10045 24259 10103 24265
rect 10045 24225 10057 24259
rect 10091 24256 10103 24259
rect 10134 24256 10140 24268
rect 10091 24228 10140 24256
rect 10091 24225 10103 24228
rect 10045 24219 10103 24225
rect 10134 24216 10140 24228
rect 10192 24216 10198 24268
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11330 24256 11336 24268
rect 11112 24228 11336 24256
rect 11112 24216 11118 24228
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 11600 24259 11658 24265
rect 11600 24225 11612 24259
rect 11646 24256 11658 24259
rect 12342 24256 12348 24268
rect 11646 24228 12348 24256
rect 11646 24225 11658 24228
rect 11600 24219 11658 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 4154 24148 4160 24200
rect 4212 24188 4218 24200
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 4212 24160 4629 24188
rect 4212 24148 4218 24160
rect 4617 24157 4629 24160
rect 4663 24157 4675 24191
rect 8018 24188 8024 24200
rect 7979 24160 8024 24188
rect 4617 24151 4675 24157
rect 8018 24148 8024 24160
rect 8076 24148 8082 24200
rect 10226 24148 10232 24200
rect 10284 24188 10290 24200
rect 10284 24160 10329 24188
rect 10284 24148 10290 24160
rect 6914 24052 6920 24064
rect 6875 24024 6920 24052
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 7190 24012 7196 24064
rect 7248 24052 7254 24064
rect 7377 24055 7435 24061
rect 7377 24052 7389 24055
rect 7248 24024 7389 24052
rect 7248 24012 7254 24024
rect 7377 24021 7389 24024
rect 7423 24021 7435 24055
rect 8386 24052 8392 24064
rect 8347 24024 8392 24052
rect 7377 24015 7435 24021
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 9217 24055 9275 24061
rect 9217 24021 9229 24055
rect 9263 24052 9275 24055
rect 9398 24052 9404 24064
rect 9263 24024 9404 24052
rect 9263 24021 9275 24024
rect 9217 24015 9275 24021
rect 9398 24012 9404 24024
rect 9456 24012 9462 24064
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 12713 24055 12771 24061
rect 12713 24052 12725 24055
rect 12492 24024 12725 24052
rect 12492 24012 12498 24024
rect 12713 24021 12725 24024
rect 12759 24021 12771 24055
rect 12713 24015 12771 24021
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 4154 23848 4160 23860
rect 4115 23820 4160 23848
rect 4154 23808 4160 23820
rect 4212 23808 4218 23860
rect 4522 23848 4528 23860
rect 4483 23820 4528 23848
rect 4522 23808 4528 23820
rect 4580 23808 4586 23860
rect 4798 23848 4804 23860
rect 4759 23820 4804 23848
rect 4798 23808 4804 23820
rect 4856 23808 4862 23860
rect 7282 23808 7288 23860
rect 7340 23848 7346 23860
rect 7742 23848 7748 23860
rect 7340 23820 7748 23848
rect 7340 23808 7346 23820
rect 7742 23808 7748 23820
rect 7800 23848 7806 23860
rect 7837 23851 7895 23857
rect 7837 23848 7849 23851
rect 7800 23820 7849 23848
rect 7800 23808 7806 23820
rect 7837 23817 7849 23820
rect 7883 23817 7895 23851
rect 7837 23811 7895 23817
rect 7926 23808 7932 23860
rect 7984 23848 7990 23860
rect 8573 23851 8631 23857
rect 8573 23848 8585 23851
rect 7984 23820 8585 23848
rect 7984 23808 7990 23820
rect 8573 23817 8585 23820
rect 8619 23848 8631 23851
rect 10226 23848 10232 23860
rect 8619 23820 10232 23848
rect 8619 23817 8631 23820
rect 8573 23811 8631 23817
rect 10226 23808 10232 23820
rect 10284 23848 10290 23860
rect 10505 23851 10563 23857
rect 10505 23848 10517 23851
rect 10284 23820 10517 23848
rect 10284 23808 10290 23820
rect 10505 23817 10517 23820
rect 10551 23817 10563 23851
rect 10505 23811 10563 23817
rect 11330 23808 11336 23860
rect 11388 23848 11394 23860
rect 11425 23851 11483 23857
rect 11425 23848 11437 23851
rect 11388 23820 11437 23848
rect 11388 23808 11394 23820
rect 11425 23817 11437 23820
rect 11471 23817 11483 23851
rect 11425 23811 11483 23817
rect 8018 23740 8024 23792
rect 8076 23780 8082 23792
rect 8205 23783 8263 23789
rect 8205 23780 8217 23783
rect 8076 23752 8217 23780
rect 8076 23740 8082 23752
rect 8205 23749 8217 23752
rect 8251 23749 8263 23783
rect 8205 23743 8263 23749
rect 10134 23740 10140 23792
rect 10192 23780 10198 23792
rect 11057 23783 11115 23789
rect 11057 23780 11069 23783
rect 10192 23752 11069 23780
rect 10192 23740 10198 23752
rect 11057 23749 11069 23752
rect 11103 23780 11115 23783
rect 11514 23780 11520 23792
rect 11103 23752 11520 23780
rect 11103 23749 11115 23752
rect 11057 23743 11115 23749
rect 11514 23740 11520 23752
rect 11572 23740 11578 23792
rect 6914 23672 6920 23724
rect 6972 23712 6978 23724
rect 7285 23715 7343 23721
rect 7285 23712 7297 23715
rect 6972 23684 7297 23712
rect 6972 23672 6978 23684
rect 7285 23681 7297 23684
rect 7331 23681 7343 23715
rect 7285 23675 7343 23681
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 6273 23647 6331 23653
rect 6273 23613 6285 23647
rect 6319 23644 6331 23647
rect 7190 23644 7196 23656
rect 6319 23616 7196 23644
rect 6319 23613 6331 23616
rect 6273 23607 6331 23613
rect 7190 23604 7196 23616
rect 7248 23604 7254 23656
rect 6641 23579 6699 23585
rect 6641 23545 6653 23579
rect 6687 23576 6699 23579
rect 7392 23576 7420 23675
rect 8662 23604 8668 23656
rect 8720 23644 8726 23656
rect 9122 23644 9128 23656
rect 8720 23616 9128 23644
rect 8720 23604 8726 23616
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 9398 23653 9404 23656
rect 9392 23644 9404 23653
rect 9359 23616 9404 23644
rect 9392 23607 9404 23616
rect 9398 23604 9404 23607
rect 9456 23604 9462 23656
rect 8110 23576 8116 23588
rect 6687 23548 8116 23576
rect 6687 23545 6699 23548
rect 6641 23539 6699 23545
rect 8110 23536 8116 23548
rect 8168 23536 8174 23588
rect 5810 23508 5816 23520
rect 5771 23480 5816 23508
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 6822 23508 6828 23520
rect 6783 23480 6828 23508
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 9033 23511 9091 23517
rect 9033 23477 9045 23511
rect 9079 23508 9091 23511
rect 9306 23508 9312 23520
rect 9079 23480 9312 23508
rect 9079 23477 9091 23480
rect 9033 23471 9091 23477
rect 9306 23468 9312 23480
rect 9364 23468 9370 23520
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12342 23508 12348 23520
rect 11931 23480 12348 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 5629 23307 5687 23313
rect 5629 23273 5641 23307
rect 5675 23304 5687 23307
rect 6181 23307 6239 23313
rect 6181 23304 6193 23307
rect 5675 23276 6193 23304
rect 5675 23273 5687 23276
rect 5629 23267 5687 23273
rect 6181 23273 6193 23276
rect 6227 23304 6239 23307
rect 6822 23304 6828 23316
rect 6227 23276 6828 23304
rect 6227 23273 6239 23276
rect 6181 23267 6239 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 6914 23264 6920 23316
rect 6972 23304 6978 23316
rect 7837 23307 7895 23313
rect 7837 23304 7849 23307
rect 6972 23276 7849 23304
rect 6972 23264 6978 23276
rect 7837 23273 7849 23276
rect 7883 23273 7895 23307
rect 7837 23267 7895 23273
rect 8205 23307 8263 23313
rect 8205 23273 8217 23307
rect 8251 23304 8263 23307
rect 8386 23304 8392 23316
rect 8251 23276 8392 23304
rect 8251 23273 8263 23276
rect 8205 23267 8263 23273
rect 8386 23264 8392 23276
rect 8444 23264 8450 23316
rect 11054 23304 11060 23316
rect 11015 23276 11060 23304
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 12526 23264 12532 23316
rect 12584 23304 12590 23316
rect 12621 23307 12679 23313
rect 12621 23304 12633 23307
rect 12584 23276 12633 23304
rect 12584 23264 12590 23276
rect 12621 23273 12633 23276
rect 12667 23273 12679 23307
rect 12621 23267 12679 23273
rect 4430 23236 4436 23248
rect 4343 23208 4436 23236
rect 4430 23196 4436 23208
rect 4488 23236 4494 23248
rect 7098 23236 7104 23248
rect 4488 23208 7104 23236
rect 4488 23196 4494 23208
rect 7098 23196 7104 23208
rect 7156 23196 7162 23248
rect 8294 23196 8300 23248
rect 8352 23236 8358 23248
rect 8662 23236 8668 23248
rect 8352 23208 8668 23236
rect 8352 23196 8358 23208
rect 8662 23196 8668 23208
rect 8720 23196 8726 23248
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 1670 23168 1676 23180
rect 1443 23140 1676 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 1670 23128 1676 23140
rect 1728 23128 1734 23180
rect 4522 23168 4528 23180
rect 4483 23140 4528 23168
rect 4522 23128 4528 23140
rect 4580 23128 4586 23180
rect 5810 23128 5816 23180
rect 5868 23168 5874 23180
rect 6089 23171 6147 23177
rect 6089 23168 6101 23171
rect 5868 23140 6101 23168
rect 5868 23128 5874 23140
rect 6089 23137 6101 23140
rect 6135 23168 6147 23171
rect 7374 23168 7380 23180
rect 6135 23140 7380 23168
rect 6135 23137 6147 23140
rect 6089 23131 6147 23137
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 7650 23128 7656 23180
rect 7708 23168 7714 23180
rect 7745 23171 7803 23177
rect 7745 23168 7757 23171
rect 7708 23140 7757 23168
rect 7708 23128 7714 23140
rect 7745 23137 7757 23140
rect 7791 23168 7803 23171
rect 8018 23168 8024 23180
rect 7791 23140 8024 23168
rect 7791 23137 7803 23140
rect 7745 23131 7803 23137
rect 8018 23128 8024 23140
rect 8076 23168 8082 23180
rect 9944 23171 10002 23177
rect 8076 23140 8432 23168
rect 8076 23128 8082 23140
rect 4614 23100 4620 23112
rect 4575 23072 4620 23100
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 6270 23100 6276 23112
rect 6231 23072 6276 23100
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 7101 23103 7159 23109
rect 7101 23069 7113 23103
rect 7147 23100 7159 23103
rect 7668 23100 7696 23128
rect 8294 23100 8300 23112
rect 7147 23072 7696 23100
rect 8255 23072 8300 23100
rect 7147 23069 7159 23072
rect 7101 23063 7159 23069
rect 8294 23060 8300 23072
rect 8352 23060 8358 23112
rect 8404 23109 8432 23140
rect 9944 23137 9956 23171
rect 9990 23168 10002 23171
rect 12434 23168 12440 23180
rect 9990 23140 12440 23168
rect 9990 23137 10002 23140
rect 9944 23131 10002 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 12529 23171 12587 23177
rect 12529 23137 12541 23171
rect 12575 23168 12587 23171
rect 12802 23168 12808 23180
rect 12575 23140 12808 23168
rect 12575 23137 12587 23140
rect 12529 23131 12587 23137
rect 12802 23128 12808 23140
rect 12860 23128 12866 23180
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23069 8447 23103
rect 8389 23063 8447 23069
rect 9122 23060 9128 23112
rect 9180 23100 9186 23112
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 9180 23072 9229 23100
rect 9180 23060 9186 23072
rect 9217 23069 9229 23072
rect 9263 23100 9275 23103
rect 9677 23103 9735 23109
rect 9677 23100 9689 23103
rect 9263 23072 9689 23100
rect 9263 23069 9275 23072
rect 9217 23063 9275 23069
rect 9677 23069 9689 23072
rect 9723 23069 9735 23103
rect 9677 23063 9735 23069
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 2777 22967 2835 22973
rect 2777 22933 2789 22967
rect 2823 22964 2835 22967
rect 3142 22964 3148 22976
rect 2823 22936 3148 22964
rect 2823 22933 2835 22936
rect 2777 22927 2835 22933
rect 3142 22924 3148 22936
rect 3200 22964 3206 22976
rect 4065 22967 4123 22973
rect 4065 22964 4077 22967
rect 3200 22936 4077 22964
rect 3200 22924 3206 22936
rect 4065 22933 4077 22936
rect 4111 22933 4123 22967
rect 5718 22964 5724 22976
rect 5679 22936 5724 22964
rect 4065 22927 4123 22933
rect 5718 22924 5724 22936
rect 5776 22924 5782 22976
rect 9692 22964 9720 23063
rect 12342 22992 12348 23044
rect 12400 23032 12406 23044
rect 12728 23032 12756 23063
rect 12400 23004 12756 23032
rect 12400 22992 12406 23004
rect 11330 22964 11336 22976
rect 9692 22936 11336 22964
rect 11330 22924 11336 22936
rect 11388 22924 11394 22976
rect 11974 22924 11980 22976
rect 12032 22964 12038 22976
rect 12161 22967 12219 22973
rect 12161 22964 12173 22967
rect 12032 22936 12173 22964
rect 12032 22924 12038 22936
rect 12161 22933 12173 22936
rect 12207 22933 12219 22967
rect 12728 22964 12756 23004
rect 13170 22964 13176 22976
rect 12728 22936 13176 22964
rect 12161 22927 12219 22933
rect 13170 22924 13176 22936
rect 13228 22924 13234 22976
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2406 22720 2412 22772
rect 2464 22760 2470 22772
rect 2501 22763 2559 22769
rect 2501 22760 2513 22763
rect 2464 22732 2513 22760
rect 2464 22720 2470 22732
rect 2501 22729 2513 22732
rect 2547 22729 2559 22763
rect 2682 22760 2688 22772
rect 2643 22732 2688 22760
rect 2501 22723 2559 22729
rect 1670 22692 1676 22704
rect 1631 22664 1676 22692
rect 1670 22652 1676 22664
rect 1728 22652 1734 22704
rect 2516 22692 2544 22723
rect 2682 22720 2688 22732
rect 2740 22720 2746 22772
rect 4157 22763 4215 22769
rect 4157 22729 4169 22763
rect 4203 22760 4215 22763
rect 4430 22760 4436 22772
rect 4203 22732 4436 22760
rect 4203 22729 4215 22732
rect 4157 22723 4215 22729
rect 4430 22720 4436 22732
rect 4488 22720 4494 22772
rect 4614 22720 4620 22772
rect 4672 22760 4678 22772
rect 5629 22763 5687 22769
rect 5629 22760 5641 22763
rect 4672 22732 5641 22760
rect 4672 22720 4678 22732
rect 5629 22729 5641 22732
rect 5675 22729 5687 22763
rect 6270 22760 6276 22772
rect 6231 22732 6276 22760
rect 5629 22723 5687 22729
rect 6270 22720 6276 22732
rect 6328 22720 6334 22772
rect 7926 22720 7932 22772
rect 7984 22760 7990 22772
rect 8021 22763 8079 22769
rect 8021 22760 8033 22763
rect 7984 22732 8033 22760
rect 7984 22720 7990 22732
rect 8021 22729 8033 22732
rect 8067 22729 8079 22763
rect 8021 22723 8079 22729
rect 7009 22695 7067 22701
rect 2516 22664 3372 22692
rect 3142 22624 3148 22636
rect 3103 22596 3148 22624
rect 3142 22584 3148 22596
rect 3200 22584 3206 22636
rect 3344 22633 3372 22664
rect 7009 22661 7021 22695
rect 7055 22692 7067 22695
rect 7742 22692 7748 22704
rect 7055 22664 7748 22692
rect 7055 22661 7067 22664
rect 7009 22655 7067 22661
rect 7742 22652 7748 22664
rect 7800 22652 7806 22704
rect 3329 22627 3387 22633
rect 3329 22593 3341 22627
rect 3375 22624 3387 22627
rect 4062 22624 4068 22636
rect 3375 22596 4068 22624
rect 3375 22593 3387 22596
rect 3329 22587 3387 22593
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 7466 22624 7472 22636
rect 7427 22596 7472 22624
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 7650 22624 7656 22636
rect 7611 22596 7656 22624
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 8036 22624 8064 22723
rect 8386 22720 8392 22772
rect 8444 22760 8450 22772
rect 8573 22763 8631 22769
rect 8573 22760 8585 22763
rect 8444 22732 8585 22760
rect 8444 22720 8450 22732
rect 8573 22729 8585 22732
rect 8619 22729 8631 22763
rect 8573 22723 8631 22729
rect 9953 22763 10011 22769
rect 9953 22729 9965 22763
rect 9999 22760 10011 22763
rect 10502 22760 10508 22772
rect 9999 22732 10508 22760
rect 9999 22729 10011 22732
rect 9953 22723 10011 22729
rect 10502 22720 10508 22732
rect 10560 22760 10566 22772
rect 11241 22763 11299 22769
rect 10560 22732 10916 22760
rect 10560 22720 10566 22732
rect 8481 22695 8539 22701
rect 8481 22661 8493 22695
rect 8527 22692 8539 22695
rect 8662 22692 8668 22704
rect 8527 22664 8668 22692
rect 8527 22661 8539 22664
rect 8481 22655 8539 22661
rect 8662 22652 8668 22664
rect 8720 22652 8726 22704
rect 9125 22627 9183 22633
rect 9125 22624 9137 22627
rect 8036 22596 9137 22624
rect 9125 22593 9137 22596
rect 9171 22624 9183 22627
rect 10689 22627 10747 22633
rect 10689 22624 10701 22627
rect 9171 22596 10701 22624
rect 9171 22593 9183 22596
rect 9125 22587 9183 22593
rect 10689 22593 10701 22596
rect 10735 22624 10747 22627
rect 10778 22624 10784 22636
rect 10735 22596 10784 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 10778 22584 10784 22596
rect 10836 22584 10842 22636
rect 4249 22559 4307 22565
rect 4249 22525 4261 22559
rect 4295 22556 4307 22559
rect 5350 22556 5356 22568
rect 4295 22528 5356 22556
rect 4295 22525 4307 22528
rect 4249 22519 4307 22525
rect 5350 22516 5356 22528
rect 5408 22516 5414 22568
rect 6641 22559 6699 22565
rect 6641 22525 6653 22559
rect 6687 22556 6699 22559
rect 7377 22559 7435 22565
rect 7377 22556 7389 22559
rect 6687 22528 7389 22556
rect 6687 22525 6699 22528
rect 6641 22519 6699 22525
rect 7377 22525 7389 22528
rect 7423 22556 7435 22559
rect 7834 22556 7840 22568
rect 7423 22528 7840 22556
rect 7423 22525 7435 22528
rect 7377 22519 7435 22525
rect 7834 22516 7840 22528
rect 7892 22516 7898 22568
rect 8662 22516 8668 22568
rect 8720 22556 8726 22568
rect 9033 22559 9091 22565
rect 9033 22556 9045 22559
rect 8720 22528 9045 22556
rect 8720 22516 8726 22528
rect 9033 22525 9045 22528
rect 9079 22525 9091 22559
rect 9033 22519 9091 22525
rect 3053 22491 3111 22497
rect 3053 22488 3065 22491
rect 2424 22460 3065 22488
rect 2424 22432 2452 22460
rect 3053 22457 3065 22460
rect 3099 22457 3111 22491
rect 3053 22451 3111 22457
rect 3789 22491 3847 22497
rect 3789 22457 3801 22491
rect 3835 22488 3847 22491
rect 4494 22491 4552 22497
rect 4494 22488 4506 22491
rect 3835 22460 4506 22488
rect 3835 22457 3847 22460
rect 3789 22451 3847 22457
rect 4494 22457 4506 22460
rect 4540 22488 4552 22491
rect 5902 22488 5908 22500
rect 4540 22460 5908 22488
rect 4540 22457 4552 22460
rect 4494 22451 4552 22457
rect 5902 22448 5908 22460
rect 5960 22448 5966 22500
rect 9677 22491 9735 22497
rect 9677 22457 9689 22491
rect 9723 22488 9735 22491
rect 9766 22488 9772 22500
rect 9723 22460 9772 22488
rect 9723 22457 9735 22460
rect 9677 22451 9735 22457
rect 9766 22448 9772 22460
rect 9824 22488 9830 22500
rect 10042 22488 10048 22500
rect 9824 22460 10048 22488
rect 9824 22448 9830 22460
rect 10042 22448 10048 22460
rect 10100 22488 10106 22500
rect 10505 22491 10563 22497
rect 10505 22488 10517 22491
rect 10100 22460 10517 22488
rect 10100 22448 10106 22460
rect 10505 22457 10517 22460
rect 10551 22457 10563 22491
rect 10505 22451 10563 22457
rect 10888 22432 10916 22732
rect 11241 22729 11253 22763
rect 11287 22760 11299 22763
rect 11330 22760 11336 22772
rect 11287 22732 11336 22760
rect 11287 22729 11299 22732
rect 11241 22723 11299 22729
rect 11330 22720 11336 22732
rect 11388 22760 11394 22772
rect 11514 22760 11520 22772
rect 11388 22732 11520 22760
rect 11388 22720 11394 22732
rect 11514 22720 11520 22732
rect 11572 22720 11578 22772
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 12250 22760 12256 22772
rect 11931 22732 12256 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 12250 22720 12256 22732
rect 12308 22760 12314 22772
rect 12526 22760 12532 22772
rect 12308 22732 12532 22760
rect 12308 22720 12314 22732
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 12894 22624 12900 22636
rect 12728 22596 12900 22624
rect 12158 22448 12164 22500
rect 12216 22488 12222 22500
rect 12253 22491 12311 22497
rect 12253 22488 12265 22491
rect 12216 22460 12265 22488
rect 12216 22448 12222 22460
rect 12253 22457 12265 22460
rect 12299 22488 12311 22491
rect 12728 22488 12756 22596
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 12986 22584 12992 22636
rect 13044 22624 13050 22636
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 13044 22596 13093 22624
rect 13044 22584 13050 22596
rect 13081 22593 13093 22596
rect 13127 22624 13139 22627
rect 13170 22624 13176 22636
rect 13127 22596 13176 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13170 22584 13176 22596
rect 13228 22624 13234 22636
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 13228 22596 13829 22624
rect 13228 22584 13234 22596
rect 13817 22593 13829 22596
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 12802 22516 12808 22568
rect 12860 22556 12866 22568
rect 13449 22559 13507 22565
rect 13449 22556 13461 22559
rect 12860 22528 13461 22556
rect 12860 22516 12866 22528
rect 13449 22525 13461 22528
rect 13495 22525 13507 22559
rect 13449 22519 13507 22525
rect 12299 22460 12756 22488
rect 12299 22457 12311 22460
rect 12253 22451 12311 22457
rect 2225 22423 2283 22429
rect 2225 22389 2237 22423
rect 2271 22420 2283 22423
rect 2406 22420 2412 22432
rect 2271 22392 2412 22420
rect 2271 22389 2283 22392
rect 2225 22383 2283 22389
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 8754 22380 8760 22432
rect 8812 22420 8818 22432
rect 8941 22423 8999 22429
rect 8941 22420 8953 22423
rect 8812 22392 8953 22420
rect 8812 22380 8818 22392
rect 8941 22389 8953 22392
rect 8987 22389 8999 22423
rect 10134 22420 10140 22432
rect 10095 22392 10140 22420
rect 8941 22383 8999 22389
rect 10134 22380 10140 22392
rect 10192 22380 10198 22432
rect 10597 22423 10655 22429
rect 10597 22389 10609 22423
rect 10643 22420 10655 22423
rect 10870 22420 10876 22432
rect 10643 22392 10876 22420
rect 10643 22389 10655 22392
rect 10597 22383 10655 22389
rect 10870 22380 10876 22392
rect 10928 22380 10934 22432
rect 12342 22380 12348 22432
rect 12400 22420 12406 22432
rect 12437 22423 12495 22429
rect 12437 22420 12449 22423
rect 12400 22392 12449 22420
rect 12400 22380 12406 22392
rect 12437 22389 12449 22392
rect 12483 22389 12495 22423
rect 12728 22420 12756 22460
rect 12897 22491 12955 22497
rect 12897 22457 12909 22491
rect 12943 22488 12955 22491
rect 13078 22488 13084 22500
rect 12943 22460 13084 22488
rect 12943 22457 12955 22460
rect 12897 22451 12955 22457
rect 13078 22448 13084 22460
rect 13136 22448 13142 22500
rect 12805 22423 12863 22429
rect 12805 22420 12817 22423
rect 12728 22392 12817 22420
rect 12437 22383 12495 22389
rect 12805 22389 12817 22392
rect 12851 22389 12863 22423
rect 12805 22383 12863 22389
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 2406 22216 2412 22228
rect 2367 22188 2412 22216
rect 2406 22176 2412 22188
rect 2464 22176 2470 22228
rect 2498 22176 2504 22228
rect 2556 22216 2562 22228
rect 2777 22219 2835 22225
rect 2777 22216 2789 22219
rect 2556 22188 2789 22216
rect 2556 22176 2562 22188
rect 2777 22185 2789 22188
rect 2823 22216 2835 22219
rect 3050 22216 3056 22228
rect 2823 22188 3056 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 3050 22176 3056 22188
rect 3108 22216 3114 22228
rect 3418 22216 3424 22228
rect 3108 22188 3424 22216
rect 3108 22176 3114 22188
rect 3418 22176 3424 22188
rect 3476 22176 3482 22228
rect 5902 22176 5908 22228
rect 5960 22216 5966 22228
rect 6181 22219 6239 22225
rect 6181 22216 6193 22219
rect 5960 22188 6193 22216
rect 5960 22176 5966 22188
rect 6181 22185 6193 22188
rect 6227 22185 6239 22219
rect 6181 22179 6239 22185
rect 7101 22219 7159 22225
rect 7101 22185 7113 22219
rect 7147 22216 7159 22219
rect 7466 22216 7472 22228
rect 7147 22188 7472 22216
rect 7147 22185 7159 22188
rect 7101 22179 7159 22185
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 10045 22219 10103 22225
rect 10045 22185 10057 22219
rect 10091 22216 10103 22219
rect 10686 22216 10692 22228
rect 10091 22188 10692 22216
rect 10091 22185 10103 22188
rect 10045 22179 10103 22185
rect 10686 22176 10692 22188
rect 10744 22216 10750 22228
rect 10744 22188 10916 22216
rect 10744 22176 10750 22188
rect 2869 22151 2927 22157
rect 2869 22117 2881 22151
rect 2915 22148 2927 22151
rect 2958 22148 2964 22160
rect 2915 22120 2964 22148
rect 2915 22117 2927 22120
rect 2869 22111 2927 22117
rect 2958 22108 2964 22120
rect 3016 22108 3022 22160
rect 5350 22148 5356 22160
rect 4816 22120 5356 22148
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 1670 22080 1676 22092
rect 1443 22052 1676 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 1670 22040 1676 22052
rect 1728 22040 1734 22092
rect 4614 22080 4620 22092
rect 3068 22052 4620 22080
rect 3068 22024 3096 22052
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 3050 22012 3056 22024
rect 2963 21984 3056 22012
rect 3050 21972 3056 21984
rect 3108 21972 3114 22024
rect 4816 22021 4844 22120
rect 5350 22108 5356 22120
rect 5408 22108 5414 22160
rect 10134 22148 10140 22160
rect 9876 22120 10140 22148
rect 5074 22089 5080 22092
rect 5068 22080 5080 22089
rect 5035 22052 5080 22080
rect 5068 22043 5080 22052
rect 5074 22040 5080 22043
rect 5132 22040 5138 22092
rect 6086 22040 6092 22092
rect 6144 22080 6150 22092
rect 6730 22080 6736 22092
rect 6144 22052 6736 22080
rect 6144 22040 6150 22052
rect 6730 22040 6736 22052
rect 6788 22040 6794 22092
rect 7650 22080 7656 22092
rect 7611 22052 7656 22080
rect 7650 22040 7656 22052
rect 7708 22040 7714 22092
rect 7742 22040 7748 22092
rect 7800 22080 7806 22092
rect 8018 22080 8024 22092
rect 7800 22052 8024 22080
rect 7800 22040 7806 22052
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 8294 22040 8300 22092
rect 8352 22080 8358 22092
rect 8941 22083 8999 22089
rect 8941 22080 8953 22083
rect 8352 22052 8953 22080
rect 8352 22040 8358 22052
rect 8941 22049 8953 22052
rect 8987 22080 8999 22083
rect 9876 22080 9904 22120
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 10226 22108 10232 22160
rect 10284 22148 10290 22160
rect 10778 22148 10784 22160
rect 10284 22120 10456 22148
rect 10739 22120 10784 22148
rect 10284 22108 10290 22120
rect 8987 22052 9904 22080
rect 9968 22052 10272 22080
rect 8987 22049 8999 22052
rect 8941 22043 8999 22049
rect 4341 22015 4399 22021
rect 4341 21981 4353 22015
rect 4387 22012 4399 22015
rect 4801 22015 4859 22021
rect 4801 22012 4813 22015
rect 4387 21984 4813 22012
rect 4387 21981 4399 21984
rect 4341 21975 4399 21981
rect 4801 21981 4813 21984
rect 4847 21981 4859 22015
rect 4801 21975 4859 21981
rect 7929 22015 7987 22021
rect 7929 21981 7941 22015
rect 7975 22012 7987 22015
rect 8110 22012 8116 22024
rect 7975 21984 8116 22012
rect 7975 21981 7987 21984
rect 7929 21975 7987 21981
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 1578 21944 1584 21956
rect 1539 21916 1584 21944
rect 1578 21904 1584 21916
rect 1636 21904 1642 21956
rect 7285 21947 7343 21953
rect 7285 21913 7297 21947
rect 7331 21944 7343 21947
rect 7374 21944 7380 21956
rect 7331 21916 7380 21944
rect 7331 21913 7343 21916
rect 7285 21907 7343 21913
rect 7374 21904 7380 21916
rect 7432 21904 7438 21956
rect 9493 21947 9551 21953
rect 9493 21913 9505 21947
rect 9539 21944 9551 21947
rect 9968 21944 9996 22052
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 9539 21916 9996 21944
rect 9539 21913 9551 21916
rect 9493 21907 9551 21913
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 4246 21876 4252 21888
rect 3927 21848 4252 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 4246 21836 4252 21848
rect 4304 21836 4310 21888
rect 8665 21879 8723 21885
rect 8665 21845 8677 21879
rect 8711 21876 8723 21879
rect 8754 21876 8760 21888
rect 8711 21848 8760 21876
rect 8711 21845 8723 21848
rect 8665 21839 8723 21845
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 9677 21879 9735 21885
rect 9677 21845 9689 21879
rect 9723 21876 9735 21879
rect 9766 21876 9772 21888
rect 9723 21848 9772 21876
rect 9723 21845 9735 21848
rect 9677 21839 9735 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 10152 21876 10180 21975
rect 10244 21944 10272 22052
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10428 22012 10456 22120
rect 10778 22108 10784 22120
rect 10836 22108 10842 22160
rect 10686 22012 10692 22024
rect 10367 21984 10692 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 10888 22012 10916 22188
rect 11054 22176 11060 22228
rect 11112 22216 11118 22228
rect 11609 22219 11667 22225
rect 11609 22216 11621 22219
rect 11112 22188 11621 22216
rect 11112 22176 11118 22188
rect 11609 22185 11621 22188
rect 11655 22216 11667 22219
rect 11974 22216 11980 22228
rect 11655 22188 11980 22216
rect 11655 22185 11667 22188
rect 11609 22179 11667 22185
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12802 22216 12808 22228
rect 12763 22188 12808 22216
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 11149 22083 11207 22089
rect 11149 22049 11161 22083
rect 11195 22080 11207 22083
rect 11701 22083 11759 22089
rect 11701 22080 11713 22083
rect 11195 22052 11713 22080
rect 11195 22049 11207 22052
rect 11149 22043 11207 22049
rect 11701 22049 11713 22052
rect 11747 22080 11759 22083
rect 12342 22080 12348 22092
rect 11747 22052 12348 22080
rect 11747 22049 11759 22052
rect 11701 22043 11759 22049
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 10888 21984 11284 22012
rect 11256 21953 11284 21984
rect 11330 21972 11336 22024
rect 11388 22012 11394 22024
rect 11885 22015 11943 22021
rect 11885 22012 11897 22015
rect 11388 21984 11897 22012
rect 11388 21972 11394 21984
rect 11885 21981 11897 21984
rect 11931 22012 11943 22015
rect 12434 22012 12440 22024
rect 11931 21984 12440 22012
rect 11931 21981 11943 21984
rect 11885 21975 11943 21981
rect 12434 21972 12440 21984
rect 12492 21972 12498 22024
rect 11241 21947 11299 21953
rect 10244 21916 10916 21944
rect 10318 21876 10324 21888
rect 10152 21848 10324 21876
rect 10318 21836 10324 21848
rect 10376 21836 10382 21888
rect 10888 21876 10916 21916
rect 11241 21913 11253 21947
rect 11287 21913 11299 21947
rect 11241 21907 11299 21913
rect 11330 21876 11336 21888
rect 10888 21848 11336 21876
rect 11330 21836 11336 21848
rect 11388 21836 11394 21888
rect 12529 21879 12587 21885
rect 12529 21845 12541 21879
rect 12575 21876 12587 21879
rect 13078 21876 13084 21888
rect 12575 21848 13084 21876
rect 12575 21845 12587 21848
rect 12529 21839 12587 21845
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 2133 21675 2191 21681
rect 2133 21641 2145 21675
rect 2179 21672 2191 21675
rect 2682 21672 2688 21684
rect 2179 21644 2688 21672
rect 2179 21641 2191 21644
rect 2133 21635 2191 21641
rect 2682 21632 2688 21644
rect 2740 21632 2746 21684
rect 4062 21672 4068 21684
rect 4023 21644 4068 21672
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 4246 21632 4252 21684
rect 4304 21672 4310 21684
rect 4522 21672 4528 21684
rect 4304 21644 4528 21672
rect 4304 21632 4310 21644
rect 4522 21632 4528 21644
rect 4580 21672 4586 21684
rect 5169 21675 5227 21681
rect 5169 21672 5181 21675
rect 4580 21644 5181 21672
rect 4580 21632 4586 21644
rect 5169 21641 5181 21644
rect 5215 21641 5227 21675
rect 5169 21635 5227 21641
rect 5902 21632 5908 21684
rect 5960 21672 5966 21684
rect 6181 21675 6239 21681
rect 6181 21672 6193 21675
rect 5960 21644 6193 21672
rect 5960 21632 5966 21644
rect 6181 21641 6193 21644
rect 6227 21641 6239 21675
rect 6181 21635 6239 21641
rect 7466 21632 7472 21684
rect 7524 21672 7530 21684
rect 8202 21672 8208 21684
rect 7524 21644 8208 21672
rect 7524 21632 7530 21644
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 10686 21672 10692 21684
rect 10428 21644 10692 21672
rect 2498 21604 2504 21616
rect 2459 21576 2504 21604
rect 2498 21564 2504 21576
rect 2556 21564 2562 21616
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 5920 21536 5948 21632
rect 9033 21607 9091 21613
rect 9033 21573 9045 21607
rect 9079 21604 9091 21607
rect 10137 21607 10195 21613
rect 10137 21604 10149 21607
rect 9079 21576 10149 21604
rect 9079 21573 9091 21576
rect 9033 21567 9091 21573
rect 10137 21573 10149 21576
rect 10183 21604 10195 21607
rect 10318 21604 10324 21616
rect 10183 21576 10324 21604
rect 10183 21573 10195 21576
rect 10137 21567 10195 21573
rect 10318 21564 10324 21576
rect 10376 21564 10382 21616
rect 5859 21508 5948 21536
rect 9769 21539 9827 21545
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 9769 21505 9781 21539
rect 9815 21536 9827 21539
rect 10428 21536 10456 21644
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11238 21632 11244 21684
rect 11296 21672 11302 21684
rect 11514 21672 11520 21684
rect 11296 21644 11520 21672
rect 11296 21632 11302 21644
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 11882 21632 11888 21684
rect 11940 21672 11946 21684
rect 12069 21675 12127 21681
rect 12069 21672 12081 21675
rect 11940 21644 12081 21672
rect 11940 21632 11946 21644
rect 12069 21641 12081 21644
rect 12115 21672 12127 21675
rect 12161 21675 12219 21681
rect 12161 21672 12173 21675
rect 12115 21644 12173 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 12161 21641 12173 21644
rect 12207 21641 12219 21675
rect 12161 21635 12219 21641
rect 12437 21607 12495 21613
rect 12437 21604 12449 21607
rect 9815 21508 10456 21536
rect 10520 21576 12449 21604
rect 9815 21505 9827 21508
rect 9769 21499 9827 21505
rect 10520 21480 10548 21576
rect 12437 21573 12449 21576
rect 12483 21573 12495 21607
rect 12437 21567 12495 21573
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 11146 21536 11152 21548
rect 10827 21508 11152 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 11146 21496 11152 21508
rect 11204 21536 11210 21548
rect 11330 21536 11336 21548
rect 11204 21508 11336 21536
rect 11204 21496 11210 21508
rect 11330 21496 11336 21508
rect 11388 21496 11394 21548
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21536 12127 21539
rect 12986 21536 12992 21548
rect 12115 21508 12848 21536
rect 12947 21508 12992 21536
rect 12115 21505 12127 21508
rect 12069 21499 12127 21505
rect 2682 21468 2688 21480
rect 2595 21440 2688 21468
rect 2682 21428 2688 21440
rect 2740 21468 2746 21480
rect 2740 21440 4752 21468
rect 2740 21428 2746 21440
rect 1765 21403 1823 21409
rect 1765 21369 1777 21403
rect 1811 21400 1823 21403
rect 2952 21403 3010 21409
rect 2952 21400 2964 21403
rect 1811 21372 2964 21400
rect 1811 21369 1823 21372
rect 1765 21363 1823 21369
rect 2952 21369 2964 21372
rect 2998 21400 3010 21403
rect 3050 21400 3056 21412
rect 2998 21372 3056 21400
rect 2998 21369 3010 21372
rect 2952 21363 3010 21369
rect 3050 21360 3056 21372
rect 3108 21360 3114 21412
rect 4724 21341 4752 21440
rect 5350 21428 5356 21480
rect 5408 21468 5414 21480
rect 6549 21471 6607 21477
rect 6549 21468 6561 21471
rect 5408 21440 6561 21468
rect 5408 21428 5414 21440
rect 6549 21437 6561 21440
rect 6595 21468 6607 21471
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6595 21440 6837 21468
rect 6595 21437 6607 21440
rect 6549 21431 6607 21437
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 7092 21471 7150 21477
rect 7092 21437 7104 21471
rect 7138 21468 7150 21471
rect 7558 21468 7564 21480
rect 7138 21440 7564 21468
rect 7138 21437 7150 21440
rect 7092 21431 7150 21437
rect 7558 21428 7564 21440
rect 7616 21428 7622 21480
rect 10042 21428 10048 21480
rect 10100 21468 10106 21480
rect 10318 21468 10324 21480
rect 10100 21440 10324 21468
rect 10100 21428 10106 21440
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 10502 21468 10508 21480
rect 10415 21440 10508 21468
rect 10502 21428 10508 21440
rect 10560 21428 10566 21480
rect 12820 21468 12848 21508
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 12820 21440 13032 21468
rect 5077 21403 5135 21409
rect 5077 21369 5089 21403
rect 5123 21400 5135 21403
rect 5123 21372 5672 21400
rect 5123 21369 5135 21372
rect 5077 21363 5135 21369
rect 4709 21335 4767 21341
rect 4709 21301 4721 21335
rect 4755 21332 4767 21335
rect 5350 21332 5356 21344
rect 4755 21304 5356 21332
rect 4755 21301 4767 21304
rect 4709 21295 4767 21301
rect 5350 21292 5356 21304
rect 5408 21292 5414 21344
rect 5534 21332 5540 21344
rect 5495 21304 5540 21332
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 5644 21341 5672 21372
rect 7282 21360 7288 21412
rect 7340 21400 7346 21412
rect 9306 21400 9312 21412
rect 7340 21372 9312 21400
rect 7340 21360 7346 21372
rect 9306 21360 9312 21372
rect 9364 21360 9370 21412
rect 9401 21403 9459 21409
rect 9401 21369 9413 21403
rect 9447 21400 9459 21403
rect 12897 21403 12955 21409
rect 12897 21400 12909 21403
rect 9447 21372 10640 21400
rect 9447 21369 9459 21372
rect 9401 21363 9459 21369
rect 10612 21344 10640 21372
rect 11808 21372 12909 21400
rect 5629 21335 5687 21341
rect 5629 21301 5641 21335
rect 5675 21332 5687 21335
rect 5902 21332 5908 21344
rect 5675 21304 5908 21332
rect 5675 21301 5687 21304
rect 5629 21295 5687 21301
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 7650 21292 7656 21344
rect 7708 21332 7714 21344
rect 8110 21332 8116 21344
rect 7708 21304 8116 21332
rect 7708 21292 7714 21304
rect 8110 21292 8116 21304
rect 8168 21332 8174 21344
rect 8205 21335 8263 21341
rect 8205 21332 8217 21335
rect 8168 21304 8217 21332
rect 8168 21292 8174 21304
rect 8205 21301 8217 21304
rect 8251 21301 8263 21335
rect 8205 21295 8263 21301
rect 10594 21292 10600 21344
rect 10652 21332 10658 21344
rect 10652 21304 10697 21332
rect 10652 21292 10658 21304
rect 11514 21292 11520 21344
rect 11572 21332 11578 21344
rect 11808 21341 11836 21372
rect 12897 21369 12909 21372
rect 12943 21369 12955 21403
rect 12897 21363 12955 21369
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11572 21304 11805 21332
rect 11572 21292 11578 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 12805 21335 12863 21341
rect 12805 21301 12817 21335
rect 12851 21332 12863 21335
rect 13004 21332 13032 21440
rect 13354 21332 13360 21344
rect 12851 21304 13360 21332
rect 12851 21301 12863 21304
rect 12805 21295 12863 21301
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 2682 21128 2688 21140
rect 2643 21100 2688 21128
rect 2682 21088 2688 21100
rect 2740 21088 2746 21140
rect 3050 21128 3056 21140
rect 3011 21100 3056 21128
rect 3050 21088 3056 21100
rect 3108 21088 3114 21140
rect 4893 21131 4951 21137
rect 4893 21097 4905 21131
rect 4939 21128 4951 21131
rect 5074 21128 5080 21140
rect 4939 21100 5080 21128
rect 4939 21097 4951 21100
rect 4893 21091 4951 21097
rect 5074 21088 5080 21100
rect 5132 21128 5138 21140
rect 6178 21128 6184 21140
rect 5132 21100 6184 21128
rect 5132 21088 5138 21100
rect 6178 21088 6184 21100
rect 6236 21128 6242 21140
rect 6733 21131 6791 21137
rect 6733 21128 6745 21131
rect 6236 21100 6745 21128
rect 6236 21088 6242 21100
rect 6733 21097 6745 21100
rect 6779 21097 6791 21131
rect 6733 21091 6791 21097
rect 7377 21131 7435 21137
rect 7377 21097 7389 21131
rect 7423 21128 7435 21131
rect 7558 21128 7564 21140
rect 7423 21100 7564 21128
rect 7423 21097 7435 21100
rect 7377 21091 7435 21097
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 8018 21088 8024 21140
rect 8076 21128 8082 21140
rect 8849 21131 8907 21137
rect 8849 21128 8861 21131
rect 8076 21100 8861 21128
rect 8076 21088 8082 21100
rect 8849 21097 8861 21100
rect 8895 21097 8907 21131
rect 9398 21128 9404 21140
rect 9359 21100 9404 21128
rect 8849 21091 8907 21097
rect 9398 21088 9404 21100
rect 9456 21088 9462 21140
rect 10502 21128 10508 21140
rect 10463 21100 10508 21128
rect 10502 21088 10508 21100
rect 10560 21088 10566 21140
rect 11054 21128 11060 21140
rect 11015 21100 11060 21128
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 11149 21131 11207 21137
rect 11149 21097 11161 21131
rect 11195 21128 11207 21131
rect 11514 21128 11520 21140
rect 11195 21100 11520 21128
rect 11195 21097 11207 21100
rect 11149 21091 11207 21097
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 12529 21131 12587 21137
rect 12529 21097 12541 21131
rect 12575 21128 12587 21131
rect 12897 21131 12955 21137
rect 12897 21128 12909 21131
rect 12575 21100 12909 21128
rect 12575 21097 12587 21100
rect 12529 21091 12587 21097
rect 12897 21097 12909 21100
rect 12943 21128 12955 21131
rect 12986 21128 12992 21140
rect 12943 21100 12992 21128
rect 12943 21097 12955 21100
rect 12897 21091 12955 21097
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 5261 21063 5319 21069
rect 5261 21029 5273 21063
rect 5307 21060 5319 21063
rect 5534 21060 5540 21072
rect 5307 21032 5540 21060
rect 5307 21029 5319 21032
rect 5261 21023 5319 21029
rect 5534 21020 5540 21032
rect 5592 21020 5598 21072
rect 7576 21060 7604 21088
rect 7576 21032 8432 21060
rect 5626 21001 5632 21004
rect 5620 20992 5632 21001
rect 5587 20964 5632 20992
rect 5620 20955 5632 20964
rect 5684 20992 5690 21004
rect 7650 20992 7656 21004
rect 5684 20964 7656 20992
rect 5626 20952 5632 20955
rect 5684 20952 5690 20964
rect 7650 20952 7656 20964
rect 7708 20952 7714 21004
rect 8202 20992 8208 21004
rect 8163 20964 8208 20992
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 1670 20924 1676 20936
rect 1631 20896 1676 20924
rect 1670 20884 1676 20896
rect 1728 20884 1734 20936
rect 5350 20924 5356 20936
rect 5311 20896 5356 20924
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 7742 20884 7748 20936
rect 7800 20924 7806 20936
rect 8404 20933 8432 21032
rect 9766 21020 9772 21072
rect 9824 21060 9830 21072
rect 11330 21060 11336 21072
rect 9824 21032 11336 21060
rect 9824 21020 9830 21032
rect 11330 21020 11336 21032
rect 11388 21060 11394 21072
rect 11609 21063 11667 21069
rect 11609 21060 11621 21063
rect 11388 21032 11621 21060
rect 11388 21020 11394 21032
rect 11609 21029 11621 21032
rect 11655 21029 11667 21063
rect 11609 21023 11667 21029
rect 9214 20952 9220 21004
rect 9272 20992 9278 21004
rect 9398 20992 9404 21004
rect 9272 20964 9404 20992
rect 9272 20952 9278 20964
rect 9398 20952 9404 20964
rect 9456 20952 9462 21004
rect 10229 20995 10287 21001
rect 10229 20961 10241 20995
rect 10275 20992 10287 20995
rect 11146 20992 11152 21004
rect 10275 20964 11152 20992
rect 10275 20961 10287 20964
rect 10229 20955 10287 20961
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 11422 20952 11428 21004
rect 11480 20992 11486 21004
rect 11517 20995 11575 21001
rect 11517 20992 11529 20995
rect 11480 20964 11529 20992
rect 11480 20952 11486 20964
rect 11517 20961 11529 20964
rect 11563 20961 11575 20995
rect 11517 20955 11575 20961
rect 13078 20952 13084 21004
rect 13136 20992 13142 21004
rect 13262 20992 13268 21004
rect 13136 20964 13268 20992
rect 13136 20952 13142 20964
rect 13262 20952 13268 20964
rect 13320 20952 13326 21004
rect 8297 20927 8355 20933
rect 8297 20924 8309 20927
rect 7800 20896 8309 20924
rect 7800 20884 7806 20896
rect 8297 20893 8309 20896
rect 8343 20893 8355 20927
rect 8297 20887 8355 20893
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20893 8447 20927
rect 8389 20887 8447 20893
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 9582 20924 9588 20936
rect 8720 20896 9588 20924
rect 8720 20884 8726 20896
rect 9582 20884 9588 20896
rect 9640 20884 9646 20936
rect 11790 20924 11796 20936
rect 11751 20896 11796 20924
rect 11790 20884 11796 20896
rect 11848 20884 11854 20936
rect 7834 20788 7840 20800
rect 7795 20760 7840 20788
rect 7834 20748 7840 20760
rect 7892 20748 7898 20800
rect 13170 20788 13176 20800
rect 13131 20760 13176 20788
rect 13170 20748 13176 20760
rect 13228 20748 13234 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 5626 20544 5632 20596
rect 5684 20584 5690 20596
rect 5721 20587 5779 20593
rect 5721 20584 5733 20587
rect 5684 20556 5733 20584
rect 5684 20544 5690 20556
rect 5721 20553 5733 20556
rect 5767 20553 5779 20587
rect 5721 20547 5779 20553
rect 7285 20587 7343 20593
rect 7285 20553 7297 20587
rect 7331 20584 7343 20587
rect 7834 20584 7840 20596
rect 7331 20556 7840 20584
rect 7331 20553 7343 20556
rect 7285 20547 7343 20553
rect 7834 20544 7840 20556
rect 7892 20544 7898 20596
rect 8202 20584 8208 20596
rect 8163 20556 8208 20584
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 10413 20587 10471 20593
rect 10413 20553 10425 20587
rect 10459 20584 10471 20587
rect 11790 20584 11796 20596
rect 10459 20556 11796 20584
rect 10459 20553 10471 20556
rect 10413 20547 10471 20553
rect 11790 20544 11796 20556
rect 11848 20584 11854 20596
rect 11885 20587 11943 20593
rect 11885 20584 11897 20587
rect 11848 20556 11897 20584
rect 11848 20544 11854 20556
rect 11885 20553 11897 20556
rect 11931 20553 11943 20587
rect 11885 20547 11943 20553
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 12492 20556 12537 20584
rect 12492 20544 12498 20556
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20448 7435 20451
rect 8220 20448 8248 20544
rect 11241 20519 11299 20525
rect 11241 20485 11253 20519
rect 11287 20516 11299 20519
rect 11330 20516 11336 20528
rect 11287 20488 11336 20516
rect 11287 20485 11299 20488
rect 11241 20479 11299 20485
rect 11330 20476 11336 20488
rect 11388 20476 11394 20528
rect 12986 20448 12992 20460
rect 7423 20420 8248 20448
rect 12947 20420 12992 20448
rect 7423 20417 7435 20420
rect 7377 20411 7435 20417
rect 12986 20408 12992 20420
rect 13044 20408 13050 20460
rect 9033 20383 9091 20389
rect 9033 20380 9045 20383
rect 8864 20352 9045 20380
rect 5350 20244 5356 20256
rect 5311 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 7742 20204 7748 20256
rect 7800 20244 7806 20256
rect 7837 20247 7895 20253
rect 7837 20244 7849 20247
rect 7800 20216 7849 20244
rect 7800 20204 7806 20216
rect 7837 20213 7849 20216
rect 7883 20213 7895 20247
rect 7837 20207 7895 20213
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 8864 20253 8892 20352
rect 9033 20349 9045 20352
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20380 12863 20383
rect 13170 20380 13176 20392
rect 12851 20352 13176 20380
rect 12851 20349 12863 20352
rect 12805 20343 12863 20349
rect 13170 20340 13176 20352
rect 13228 20340 13234 20392
rect 9300 20315 9358 20321
rect 9300 20281 9312 20315
rect 9346 20312 9358 20315
rect 9490 20312 9496 20324
rect 9346 20284 9496 20312
rect 9346 20281 9358 20284
rect 9300 20275 9358 20281
rect 9490 20272 9496 20284
rect 9548 20272 9554 20324
rect 12894 20312 12900 20324
rect 12855 20284 12900 20312
rect 12894 20272 12900 20284
rect 12952 20312 12958 20324
rect 13449 20315 13507 20321
rect 13449 20312 13461 20315
rect 12952 20284 13461 20312
rect 12952 20272 12958 20284
rect 13449 20281 13461 20284
rect 13495 20281 13507 20315
rect 13449 20275 13507 20281
rect 8849 20247 8907 20253
rect 8849 20244 8861 20247
rect 8352 20216 8861 20244
rect 8352 20204 8358 20216
rect 8849 20213 8861 20216
rect 8895 20213 8907 20247
rect 8849 20207 8907 20213
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11480 20216 11529 20244
rect 11480 20204 11486 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 7558 20000 7564 20052
rect 7616 20040 7622 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 7616 20012 7849 20040
rect 7616 20000 7622 20012
rect 7837 20009 7849 20012
rect 7883 20009 7895 20043
rect 10042 20040 10048 20052
rect 10003 20012 10048 20040
rect 7837 20003 7895 20009
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 10502 20040 10508 20052
rect 10463 20012 10508 20040
rect 10502 20000 10508 20012
rect 10560 20000 10566 20052
rect 12986 20040 12992 20052
rect 12947 20012 12992 20040
rect 12986 20000 12992 20012
rect 13044 20000 13050 20052
rect 11876 19975 11934 19981
rect 11876 19941 11888 19975
rect 11922 19972 11934 19975
rect 11974 19972 11980 19984
rect 11922 19944 11980 19972
rect 11922 19941 11934 19944
rect 11876 19935 11934 19941
rect 11974 19932 11980 19944
rect 12032 19932 12038 19984
rect 10042 19864 10048 19916
rect 10100 19904 10106 19916
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 10100 19876 10425 19904
rect 10100 19864 10106 19876
rect 10413 19873 10425 19876
rect 10459 19904 10471 19907
rect 10962 19904 10968 19916
rect 10459 19876 10968 19904
rect 10459 19873 10471 19876
rect 10413 19867 10471 19873
rect 10962 19864 10968 19876
rect 11020 19864 11026 19916
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11609 19907 11667 19913
rect 11609 19904 11621 19907
rect 11296 19876 11621 19904
rect 11296 19864 11302 19876
rect 11609 19873 11621 19876
rect 11655 19873 11667 19907
rect 11609 19867 11667 19873
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19836 10747 19839
rect 11146 19836 11152 19848
rect 10735 19808 11152 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 9953 19771 10011 19777
rect 9953 19737 9965 19771
rect 9999 19768 10011 19771
rect 10704 19768 10732 19799
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 9999 19740 10732 19768
rect 9999 19737 10011 19740
rect 9953 19731 10011 19737
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7282 19700 7288 19712
rect 6963 19672 7288 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8846 19700 8852 19712
rect 8527 19672 8852 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9125 19703 9183 19709
rect 9125 19669 9137 19703
rect 9171 19700 9183 19703
rect 9490 19700 9496 19712
rect 9171 19672 9496 19700
rect 9171 19669 9183 19672
rect 9125 19663 9183 19669
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 11238 19456 11244 19508
rect 11296 19496 11302 19508
rect 11885 19499 11943 19505
rect 11885 19496 11897 19499
rect 11296 19468 11897 19496
rect 11296 19456 11302 19468
rect 11885 19465 11897 19468
rect 11931 19465 11943 19499
rect 11885 19459 11943 19465
rect 6641 19431 6699 19437
rect 6641 19397 6653 19431
rect 6687 19428 6699 19431
rect 6687 19400 7512 19428
rect 6687 19397 6699 19400
rect 6641 19391 6699 19397
rect 7484 19372 7512 19400
rect 7466 19360 7472 19372
rect 7427 19332 7472 19360
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19329 8999 19363
rect 11146 19360 11152 19372
rect 11107 19332 11152 19360
rect 8941 19323 8999 19329
rect 8018 19252 8024 19304
rect 8076 19292 8082 19304
rect 8202 19292 8208 19304
rect 8076 19264 8208 19292
rect 8076 19252 8082 19264
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 8386 19292 8392 19304
rect 8343 19264 8392 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 8386 19252 8392 19264
rect 8444 19292 8450 19304
rect 8956 19292 8984 19323
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 8444 19264 8984 19292
rect 8444 19252 8450 19264
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 10686 19292 10692 19304
rect 9916 19264 10692 19292
rect 9916 19252 9922 19264
rect 10686 19252 10692 19264
rect 10744 19292 10750 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 10744 19264 10977 19292
rect 10744 19252 10750 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 6273 19227 6331 19233
rect 6273 19193 6285 19227
rect 6319 19224 6331 19227
rect 6638 19224 6644 19236
rect 6319 19196 6644 19224
rect 6319 19193 6331 19196
rect 6273 19187 6331 19193
rect 6638 19184 6644 19196
rect 6696 19184 6702 19236
rect 7929 19227 7987 19233
rect 7929 19193 7941 19227
rect 7975 19224 7987 19227
rect 10137 19227 10195 19233
rect 7975 19196 8800 19224
rect 7975 19193 7987 19196
rect 7929 19187 7987 19193
rect 8772 19168 8800 19196
rect 10137 19193 10149 19227
rect 10183 19224 10195 19227
rect 10594 19224 10600 19236
rect 10183 19196 10600 19224
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 10594 19184 10600 19196
rect 10652 19184 10658 19236
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 10873 19227 10931 19233
rect 10873 19224 10885 19227
rect 10836 19196 10885 19224
rect 10836 19184 10842 19196
rect 10873 19193 10885 19196
rect 10919 19224 10931 19227
rect 11514 19224 11520 19236
rect 10919 19196 11520 19224
rect 10919 19193 10931 19196
rect 10873 19187 10931 19193
rect 11514 19184 11520 19196
rect 11572 19184 11578 19236
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7190 19156 7196 19168
rect 6880 19128 6925 19156
rect 7151 19128 7196 19156
rect 6880 19116 6886 19128
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 7340 19128 7385 19156
rect 7340 19116 7346 19128
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 8389 19159 8447 19165
rect 8389 19156 8401 19159
rect 8352 19128 8401 19156
rect 8352 19116 8358 19128
rect 8389 19125 8401 19128
rect 8435 19125 8447 19159
rect 8754 19156 8760 19168
rect 8715 19128 8760 19156
rect 8389 19119 8447 19125
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 8849 19159 8907 19165
rect 8849 19125 8861 19159
rect 8895 19156 8907 19159
rect 9030 19156 9036 19168
rect 8895 19128 9036 19156
rect 8895 19125 8907 19128
rect 8849 19119 8907 19125
rect 9030 19116 9036 19128
rect 9088 19156 9094 19168
rect 9582 19156 9588 19168
rect 9088 19128 9588 19156
rect 9088 19116 9094 19128
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 9769 19159 9827 19165
rect 9769 19125 9781 19159
rect 9815 19156 9827 19159
rect 9858 19156 9864 19168
rect 9815 19128 9864 19156
rect 9815 19125 9827 19128
rect 9769 19119 9827 19125
rect 9858 19116 9864 19128
rect 9916 19156 9922 19168
rect 10042 19156 10048 19168
rect 9916 19128 10048 19156
rect 9916 19116 9922 19128
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10502 19156 10508 19168
rect 10463 19128 10508 19156
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 6638 18912 6644 18964
rect 6696 18952 6702 18964
rect 7190 18952 7196 18964
rect 6696 18924 7196 18952
rect 6696 18912 6702 18924
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10318 18952 10324 18964
rect 10091 18924 10324 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 10686 18952 10692 18964
rect 10647 18924 10692 18952
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 11146 18952 11152 18964
rect 11059 18924 11152 18952
rect 11146 18912 11152 18924
rect 11204 18952 11210 18964
rect 11701 18955 11759 18961
rect 11701 18952 11713 18955
rect 11204 18924 11713 18952
rect 11204 18912 11210 18924
rect 11701 18921 11713 18924
rect 11747 18952 11759 18955
rect 11974 18952 11980 18964
rect 11747 18924 11980 18952
rect 11747 18921 11759 18924
rect 11701 18915 11759 18921
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18816 5227 18819
rect 5258 18816 5264 18828
rect 5215 18788 5264 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5442 18825 5448 18828
rect 5436 18816 5448 18825
rect 5403 18788 5448 18816
rect 5436 18779 5448 18788
rect 5442 18776 5448 18779
rect 5500 18776 5506 18828
rect 8202 18816 8208 18828
rect 8163 18788 8208 18816
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 10594 18816 10600 18828
rect 9916 18788 10600 18816
rect 9916 18776 9922 18788
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 8294 18748 8300 18760
rect 8255 18720 8300 18748
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 10137 18751 10195 18757
rect 10137 18717 10149 18751
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10962 18748 10968 18760
rect 10367 18720 10968 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 7650 18640 7656 18692
rect 7708 18680 7714 18692
rect 8404 18680 8432 18711
rect 9490 18680 9496 18692
rect 7708 18652 9496 18680
rect 7708 18640 7714 18652
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 9858 18640 9864 18692
rect 9916 18680 9922 18692
rect 10152 18680 10180 18711
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 10870 18680 10876 18692
rect 9916 18652 10876 18680
rect 9916 18640 9922 18652
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 6178 18572 6184 18624
rect 6236 18612 6242 18624
rect 6549 18615 6607 18621
rect 6549 18612 6561 18615
rect 6236 18584 6561 18612
rect 6236 18572 6242 18584
rect 6549 18581 6561 18584
rect 6595 18581 6607 18615
rect 7834 18612 7840 18624
rect 7795 18584 7840 18612
rect 6549 18575 6607 18581
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 9674 18612 9680 18624
rect 9635 18584 9680 18612
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 7285 18411 7343 18417
rect 7285 18377 7297 18411
rect 7331 18408 7343 18411
rect 8294 18408 8300 18420
rect 7331 18380 8300 18408
rect 7331 18377 7343 18380
rect 7285 18371 7343 18377
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 9490 18408 9496 18420
rect 9451 18380 9496 18408
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 10413 18411 10471 18417
rect 10413 18408 10425 18411
rect 10376 18380 10425 18408
rect 10376 18368 10382 18380
rect 10413 18377 10425 18380
rect 10459 18377 10471 18411
rect 10413 18371 10471 18377
rect 7650 18340 7656 18352
rect 7611 18312 7656 18340
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 1946 18272 1952 18284
rect 1412 18244 1952 18272
rect 1412 18213 1440 18244
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 5350 18232 5356 18284
rect 5408 18272 5414 18284
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5408 18244 5641 18272
rect 5408 18232 5414 18244
rect 5629 18241 5641 18244
rect 5675 18272 5687 18275
rect 5902 18272 5908 18284
rect 5675 18244 5908 18272
rect 5675 18241 5687 18244
rect 5629 18235 5687 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18173 1455 18207
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 1397 18167 1455 18173
rect 3528 18176 3617 18204
rect 3528 18080 3556 18176
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 3605 18167 3663 18173
rect 8018 18164 8024 18216
rect 8076 18204 8082 18216
rect 8113 18207 8171 18213
rect 8113 18204 8125 18207
rect 8076 18176 8125 18204
rect 8076 18164 8082 18176
rect 8113 18173 8125 18176
rect 8159 18173 8171 18207
rect 8113 18167 8171 18173
rect 3878 18145 3884 18148
rect 3872 18136 3884 18145
rect 3839 18108 3884 18136
rect 3872 18099 3884 18108
rect 3878 18096 3884 18099
rect 3936 18096 3942 18148
rect 5442 18136 5448 18148
rect 5000 18108 5448 18136
rect 3510 18068 3516 18080
rect 3471 18040 3516 18068
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 4062 18028 4068 18080
rect 4120 18068 4126 18080
rect 5000 18077 5028 18108
rect 5442 18096 5448 18108
rect 5500 18136 5506 18148
rect 5905 18139 5963 18145
rect 5905 18136 5917 18139
rect 5500 18108 5917 18136
rect 5500 18096 5506 18108
rect 5905 18105 5917 18108
rect 5951 18105 5963 18139
rect 5905 18099 5963 18105
rect 4985 18071 5043 18077
rect 4985 18068 4997 18071
rect 4120 18040 4997 18068
rect 4120 18028 4126 18040
rect 4985 18037 4997 18040
rect 5031 18037 5043 18071
rect 4985 18031 5043 18037
rect 8021 18071 8079 18077
rect 8021 18037 8033 18071
rect 8067 18068 8079 18071
rect 8128 18068 8156 18167
rect 8386 18145 8392 18148
rect 8380 18136 8392 18145
rect 8347 18108 8392 18136
rect 8380 18099 8392 18108
rect 8386 18096 8392 18099
rect 8444 18096 8450 18148
rect 8294 18068 8300 18080
rect 8067 18040 8300 18068
rect 8067 18037 8079 18040
rect 8021 18031 8079 18037
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9916 18040 10057 18068
rect 9916 18028 9922 18040
rect 10045 18037 10057 18040
rect 10091 18037 10103 18071
rect 10045 18031 10103 18037
rect 10873 18071 10931 18077
rect 10873 18037 10885 18071
rect 10919 18068 10931 18071
rect 10962 18068 10968 18080
rect 10919 18040 10968 18068
rect 10919 18037 10931 18040
rect 10873 18031 10931 18037
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 7466 17864 7472 17876
rect 7423 17836 7472 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 9732 17836 10149 17864
rect 9732 17824 9738 17836
rect 10137 17833 10149 17836
rect 10183 17864 10195 17867
rect 11146 17864 11152 17876
rect 10183 17836 11152 17864
rect 10183 17833 10195 17836
rect 10137 17827 10195 17833
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 6178 17756 6184 17808
rect 6236 17805 6242 17808
rect 6236 17799 6300 17805
rect 6236 17765 6254 17799
rect 6288 17765 6300 17799
rect 6236 17759 6300 17765
rect 6236 17756 6242 17759
rect 11974 17756 11980 17808
rect 12032 17805 12038 17808
rect 12032 17799 12096 17805
rect 12032 17765 12050 17799
rect 12084 17765 12096 17799
rect 12032 17759 12096 17765
rect 12032 17756 12038 17759
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4798 17728 4804 17740
rect 4387 17700 4804 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 4890 17688 4896 17740
rect 4948 17728 4954 17740
rect 4948 17700 4993 17728
rect 4948 17688 4954 17700
rect 5718 17688 5724 17740
rect 5776 17728 5782 17740
rect 6086 17728 6092 17740
rect 5776 17700 6092 17728
rect 5776 17688 5782 17700
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9824 17700 10057 17728
rect 9824 17688 9830 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5902 17620 5908 17672
rect 5960 17660 5966 17672
rect 5997 17663 6055 17669
rect 5997 17660 6009 17663
rect 5960 17632 6009 17660
rect 5960 17620 5966 17632
rect 5997 17629 6009 17632
rect 6043 17629 6055 17663
rect 5997 17623 6055 17629
rect 8202 17620 8208 17672
rect 8260 17660 8266 17672
rect 8481 17663 8539 17669
rect 8481 17660 8493 17663
rect 8260 17632 8493 17660
rect 8260 17620 8266 17632
rect 8481 17629 8493 17632
rect 8527 17629 8539 17663
rect 10318 17660 10324 17672
rect 10279 17632 10324 17660
rect 8481 17623 8539 17629
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 11422 17620 11428 17672
rect 11480 17660 11486 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11480 17632 11805 17660
rect 11480 17620 11486 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 3697 17595 3755 17601
rect 3697 17561 3709 17595
rect 3743 17592 3755 17595
rect 3878 17592 3884 17604
rect 3743 17564 3884 17592
rect 3743 17561 3755 17564
rect 3697 17555 3755 17561
rect 3878 17552 3884 17564
rect 3936 17592 3942 17604
rect 5000 17592 5028 17620
rect 8386 17592 8392 17604
rect 3936 17564 5028 17592
rect 8220 17564 8392 17592
rect 3936 17552 3942 17564
rect 3970 17484 3976 17536
rect 4028 17524 4034 17536
rect 4433 17527 4491 17533
rect 4433 17524 4445 17527
rect 4028 17496 4445 17524
rect 4028 17484 4034 17496
rect 4433 17493 4445 17496
rect 4479 17493 4491 17527
rect 4433 17487 4491 17493
rect 8018 17484 8024 17536
rect 8076 17524 8082 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 8076 17496 8125 17524
rect 8076 17484 8082 17496
rect 8113 17493 8125 17496
rect 8159 17524 8171 17527
rect 8220 17524 8248 17564
rect 8386 17552 8392 17564
rect 8444 17552 8450 17604
rect 9674 17592 9680 17604
rect 9635 17564 9680 17592
rect 9674 17552 9680 17564
rect 9732 17552 9738 17604
rect 8159 17496 8248 17524
rect 9309 17527 9367 17533
rect 8159 17493 8171 17496
rect 8113 17487 8171 17493
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9490 17524 9496 17536
rect 9355 17496 9496 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9490 17484 9496 17496
rect 9548 17484 9554 17536
rect 13170 17524 13176 17536
rect 13131 17496 13176 17524
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 4798 17280 4804 17332
rect 4856 17320 4862 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 4856 17292 6837 17320
rect 4856 17280 4862 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 6825 17283 6883 17289
rect 10318 17280 10324 17332
rect 10376 17320 10382 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 10376 17292 10609 17320
rect 10376 17280 10382 17292
rect 10597 17289 10609 17292
rect 10643 17289 10655 17323
rect 11146 17320 11152 17332
rect 11107 17292 11152 17320
rect 10597 17283 10655 17289
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 12032 17292 12173 17320
rect 12032 17280 12038 17292
rect 12161 17289 12173 17292
rect 12207 17289 12219 17323
rect 12161 17283 12219 17289
rect 5721 17255 5779 17261
rect 5721 17221 5733 17255
rect 5767 17252 5779 17255
rect 6178 17252 6184 17264
rect 5767 17224 6184 17252
rect 5767 17221 5779 17224
rect 5721 17215 5779 17221
rect 6178 17212 6184 17224
rect 6236 17212 6242 17264
rect 6288 17224 7512 17252
rect 5902 17184 5908 17196
rect 5736 17156 5908 17184
rect 3510 17116 3516 17128
rect 3423 17088 3516 17116
rect 3510 17076 3516 17088
rect 3568 17116 3574 17128
rect 3605 17119 3663 17125
rect 3605 17116 3617 17119
rect 3568 17088 3617 17116
rect 3568 17076 3574 17088
rect 3605 17085 3617 17088
rect 3651 17116 3663 17119
rect 5736 17116 5764 17156
rect 5902 17144 5908 17156
rect 5960 17184 5966 17196
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 5960 17156 6101 17184
rect 5960 17144 5966 17156
rect 6089 17153 6101 17156
rect 6135 17184 6147 17187
rect 6288 17184 6316 17224
rect 6135 17156 6316 17184
rect 6135 17153 6147 17156
rect 6089 17147 6147 17153
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6822 17184 6828 17196
rect 6696 17156 6828 17184
rect 6696 17144 6702 17156
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17153 7435 17187
rect 7484 17184 7512 17224
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 8662 17252 8668 17264
rect 8352 17224 8668 17252
rect 8352 17212 8358 17224
rect 8662 17212 8668 17224
rect 8720 17212 8726 17264
rect 7484 17156 8432 17184
rect 7377 17147 7435 17153
rect 3651 17088 5764 17116
rect 3651 17085 3663 17088
rect 3605 17079 3663 17085
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 7392 17116 7420 17147
rect 8404 17128 8432 17156
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 5868 17088 7849 17116
rect 5868 17076 5874 17088
rect 7837 17085 7849 17088
rect 7883 17085 7895 17119
rect 7837 17079 7895 17085
rect 8386 17076 8392 17128
rect 8444 17116 8450 17128
rect 9214 17116 9220 17128
rect 8444 17088 9220 17116
rect 8444 17076 8450 17088
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 9490 17125 9496 17128
rect 9484 17116 9496 17125
rect 9451 17088 9496 17116
rect 9484 17079 9496 17088
rect 9490 17076 9496 17079
rect 9548 17076 9554 17128
rect 3872 17051 3930 17057
rect 3872 17017 3884 17051
rect 3918 17048 3930 17051
rect 4246 17048 4252 17060
rect 3918 17020 4252 17048
rect 3918 17017 3930 17020
rect 3872 17011 3930 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 6730 17048 6736 17060
rect 6564 17020 6736 17048
rect 4614 16940 4620 16992
rect 4672 16980 4678 16992
rect 4982 16980 4988 16992
rect 4672 16952 4988 16980
rect 4672 16940 4678 16952
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 5902 16940 5908 16992
rect 5960 16980 5966 16992
rect 6564 16989 6592 17020
rect 6730 17008 6736 17020
rect 6788 17048 6794 17060
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 6788 17020 7297 17048
rect 6788 17008 6794 17020
rect 7285 17017 7297 17020
rect 7331 17017 7343 17051
rect 7285 17011 7343 17017
rect 7466 17008 7472 17060
rect 7524 17048 7530 17060
rect 9033 17051 9091 17057
rect 9033 17048 9045 17051
rect 7524 17020 9045 17048
rect 7524 17008 7530 17020
rect 9033 17017 9045 17020
rect 9079 17048 9091 17051
rect 9766 17048 9772 17060
rect 9079 17020 9772 17048
rect 9079 17017 9091 17020
rect 9033 17011 9091 17017
rect 9766 17008 9772 17020
rect 9824 17008 9830 17060
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 5960 16952 6561 16980
rect 5960 16940 5966 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7193 16983 7251 16989
rect 7193 16980 7205 16983
rect 6972 16952 7205 16980
rect 6972 16940 6978 16952
rect 7193 16949 7205 16952
rect 7239 16949 7251 16983
rect 7193 16943 7251 16949
rect 8478 16940 8484 16992
rect 8536 16980 8542 16992
rect 9490 16980 9496 16992
rect 8536 16952 9496 16980
rect 8536 16940 8542 16952
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11480 16952 11805 16980
rect 11480 16940 11486 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 11793 16943 11851 16949
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 4890 16776 4896 16788
rect 4851 16748 4896 16776
rect 4890 16736 4896 16748
rect 4948 16776 4954 16788
rect 5261 16779 5319 16785
rect 5261 16776 5273 16779
rect 4948 16748 5273 16776
rect 4948 16736 4954 16748
rect 5261 16745 5273 16748
rect 5307 16745 5319 16779
rect 5261 16739 5319 16745
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6457 16779 6515 16785
rect 6457 16776 6469 16779
rect 6236 16748 6469 16776
rect 6236 16736 6242 16748
rect 6457 16745 6469 16748
rect 6503 16745 6515 16779
rect 6457 16739 6515 16745
rect 7193 16779 7251 16785
rect 7193 16745 7205 16779
rect 7239 16776 7251 16779
rect 7282 16776 7288 16788
rect 7239 16748 7288 16776
rect 7239 16745 7251 16748
rect 7193 16739 7251 16745
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 7708 16748 7753 16776
rect 7708 16736 7714 16748
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 9306 16776 9312 16788
rect 8720 16748 9312 16776
rect 8720 16736 8726 16748
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9953 16779 10011 16785
rect 9953 16745 9965 16779
rect 9999 16776 10011 16779
rect 10318 16776 10324 16788
rect 9999 16748 10324 16776
rect 9999 16745 10011 16748
rect 9953 16739 10011 16745
rect 5534 16668 5540 16720
rect 5592 16708 5598 16720
rect 5721 16711 5779 16717
rect 5721 16708 5733 16711
rect 5592 16680 5733 16708
rect 5592 16668 5598 16680
rect 5721 16677 5733 16680
rect 5767 16677 5779 16711
rect 5721 16671 5779 16677
rect 8849 16711 8907 16717
rect 8849 16677 8861 16711
rect 8895 16708 8907 16711
rect 9582 16708 9588 16720
rect 8895 16680 9588 16708
rect 8895 16677 8907 16680
rect 8849 16671 8907 16677
rect 9582 16668 9588 16680
rect 9640 16708 9646 16720
rect 9968 16708 9996 16739
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11885 16779 11943 16785
rect 11885 16776 11897 16779
rect 11020 16748 11897 16776
rect 11020 16736 11026 16748
rect 11885 16745 11897 16748
rect 11931 16745 11943 16779
rect 11885 16739 11943 16745
rect 11422 16708 11428 16720
rect 9640 16680 9996 16708
rect 10520 16680 11428 16708
rect 9640 16668 9646 16680
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 5626 16640 5632 16652
rect 4396 16612 5632 16640
rect 4396 16600 4402 16612
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16640 7619 16643
rect 7607 16612 8340 16640
rect 7607 16609 7619 16612
rect 7561 16603 7619 16609
rect 5810 16572 5816 16584
rect 5723 16544 5816 16572
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 7742 16572 7748 16584
rect 7703 16544 7748 16572
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 8312 16572 8340 16612
rect 9214 16600 9220 16652
rect 9272 16640 9278 16652
rect 10520 16649 10548 16680
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 10778 16649 10784 16652
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 9272 16612 9321 16640
rect 9272 16600 9278 16612
rect 9309 16609 9321 16612
rect 9355 16640 9367 16643
rect 10505 16643 10563 16649
rect 10505 16640 10517 16643
rect 9355 16612 10517 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 10505 16609 10517 16612
rect 10551 16609 10563 16643
rect 10772 16640 10784 16649
rect 10739 16612 10784 16640
rect 10505 16603 10563 16609
rect 10772 16603 10784 16612
rect 10778 16600 10784 16603
rect 10836 16600 10842 16652
rect 8386 16572 8392 16584
rect 8312 16544 8392 16572
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 5828 16504 5856 16532
rect 4264 16476 5856 16504
rect 4264 16448 4292 16476
rect 3697 16439 3755 16445
rect 3697 16405 3709 16439
rect 3743 16436 3755 16439
rect 4246 16436 4252 16448
rect 3743 16408 4252 16436
rect 3743 16405 3755 16408
rect 3697 16399 3755 16405
rect 4246 16396 4252 16408
rect 4304 16396 4310 16448
rect 4525 16439 4583 16445
rect 4525 16405 4537 16439
rect 4571 16436 4583 16439
rect 4614 16436 4620 16448
rect 4571 16408 4620 16436
rect 4571 16405 4583 16408
rect 4525 16399 4583 16405
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 10413 16439 10471 16445
rect 10413 16405 10425 16439
rect 10459 16436 10471 16439
rect 10778 16436 10784 16448
rect 10459 16408 10784 16436
rect 10459 16405 10471 16408
rect 10413 16399 10471 16405
rect 10778 16396 10784 16408
rect 10836 16396 10842 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 7190 16232 7196 16244
rect 7151 16204 7196 16232
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 7558 16232 7564 16244
rect 7340 16204 7564 16232
rect 7340 16192 7346 16204
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8386 16232 8392 16244
rect 8343 16204 8392 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8754 16232 8760 16244
rect 8715 16204 8760 16232
rect 8754 16192 8760 16204
rect 8812 16192 8818 16244
rect 8846 16192 8852 16244
rect 8904 16232 8910 16244
rect 8904 16204 9260 16232
rect 8904 16192 8910 16204
rect 2317 16167 2375 16173
rect 2317 16133 2329 16167
rect 2363 16164 2375 16167
rect 3513 16167 3571 16173
rect 3513 16164 3525 16167
rect 2363 16136 3525 16164
rect 2363 16133 2375 16136
rect 2317 16127 2375 16133
rect 1946 16096 1952 16108
rect 1412 16068 1952 16096
rect 1412 16037 1440 16068
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 2424 16037 2452 16136
rect 3513 16133 3525 16136
rect 3559 16133 3571 16167
rect 3513 16127 3571 16133
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16096 3479 16099
rect 4062 16096 4068 16108
rect 3467 16068 4068 16096
rect 3467 16065 3479 16068
rect 3421 16059 3479 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 6822 16096 6828 16108
rect 5583 16068 6828 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16096 7159 16099
rect 7282 16096 7288 16108
rect 7147 16068 7288 16096
rect 7147 16065 7159 16068
rect 7101 16059 7159 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 7742 16096 7748 16108
rect 7703 16068 7748 16096
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 9232 16105 9260 16204
rect 10226 16192 10232 16244
rect 10284 16232 10290 16244
rect 10594 16232 10600 16244
rect 10284 16204 10600 16232
rect 10284 16192 10290 16204
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 10318 16164 10324 16176
rect 10279 16136 10324 16164
rect 10318 16124 10324 16136
rect 10376 16124 10382 16176
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16096 9367 16099
rect 9582 16096 9588 16108
rect 9355 16068 9588 16096
rect 9355 16065 9367 16068
rect 9309 16059 9367 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 15997 2467 16031
rect 2409 15991 2467 15997
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3099 16000 3893 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 3881 15997 3893 16000
rect 3927 16028 3939 16031
rect 3970 16028 3976 16040
rect 3927 16000 3976 16028
rect 3927 15997 3939 16000
rect 3881 15991 3939 15997
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 8711 16000 9137 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 9125 15997 9137 16000
rect 9171 16028 9183 16031
rect 9398 16028 9404 16040
rect 9171 16000 9404 16028
rect 9171 15997 9183 16000
rect 9125 15991 9183 15997
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 5534 15960 5540 15972
rect 3896 15932 5540 15960
rect 3896 15904 3924 15932
rect 5534 15920 5540 15932
rect 5592 15960 5598 15972
rect 5997 15963 6055 15969
rect 5997 15960 6009 15963
rect 5592 15932 6009 15960
rect 5592 15920 5598 15932
rect 5997 15929 6009 15932
rect 6043 15929 6055 15963
rect 7558 15960 7564 15972
rect 7471 15932 7564 15960
rect 5997 15923 6055 15929
rect 7558 15920 7564 15932
rect 7616 15960 7622 15972
rect 8846 15960 8852 15972
rect 7616 15932 8852 15960
rect 7616 15920 7622 15932
rect 8846 15920 8852 15932
rect 8904 15920 8910 15972
rect 9306 15920 9312 15972
rect 9364 15960 9370 15972
rect 9508 15960 9536 16068
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 10870 16096 10876 16108
rect 10275 16068 10876 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 9364 15932 9536 15960
rect 9861 15963 9919 15969
rect 9364 15920 9370 15932
rect 9861 15929 9873 15963
rect 9907 15960 9919 15963
rect 10686 15960 10692 15972
rect 9907 15932 10692 15960
rect 9907 15929 9919 15932
rect 9861 15923 9919 15929
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 2593 15895 2651 15901
rect 2593 15861 2605 15895
rect 2639 15892 2651 15895
rect 2774 15892 2780 15904
rect 2639 15864 2780 15892
rect 2639 15861 2651 15864
rect 2593 15855 2651 15861
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 3878 15852 3884 15904
rect 3936 15852 3942 15904
rect 3973 15895 4031 15901
rect 3973 15861 3985 15895
rect 4019 15892 4031 15895
rect 4062 15892 4068 15904
rect 4019 15864 4068 15892
rect 4019 15861 4031 15864
rect 3973 15855 4031 15861
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4246 15852 4252 15904
rect 4304 15892 4310 15904
rect 4706 15892 4712 15904
rect 4304 15864 4712 15892
rect 4304 15852 4310 15864
rect 4706 15852 4712 15864
rect 4764 15892 4770 15904
rect 4893 15895 4951 15901
rect 4893 15892 4905 15895
rect 4764 15864 4905 15892
rect 4764 15852 4770 15864
rect 4893 15861 4905 15864
rect 4939 15861 4951 15895
rect 4893 15855 4951 15861
rect 5074 15852 5080 15904
rect 5132 15892 5138 15904
rect 5261 15895 5319 15901
rect 5261 15892 5273 15895
rect 5132 15864 5273 15892
rect 5132 15852 5138 15864
rect 5261 15861 5273 15864
rect 5307 15892 5319 15895
rect 5626 15892 5632 15904
rect 5307 15864 5632 15892
rect 5307 15861 5319 15864
rect 5261 15855 5319 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7466 15892 7472 15904
rect 6687 15864 7472 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7466 15852 7472 15864
rect 7524 15892 7530 15904
rect 7653 15895 7711 15901
rect 7653 15892 7665 15895
rect 7524 15864 7665 15892
rect 7524 15852 7530 15864
rect 7653 15861 7665 15864
rect 7699 15861 7711 15895
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 7653 15855 7711 15861
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11422 15892 11428 15904
rect 11383 15864 11428 15892
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 3605 15691 3663 15697
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 4062 15688 4068 15700
rect 3651 15660 4068 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 6178 15648 6184 15700
rect 6236 15688 6242 15700
rect 6641 15691 6699 15697
rect 6641 15688 6653 15691
rect 6236 15660 6653 15688
rect 6236 15648 6242 15660
rect 6641 15657 6653 15660
rect 6687 15657 6699 15691
rect 6641 15651 6699 15657
rect 7101 15691 7159 15697
rect 7101 15657 7113 15691
rect 7147 15688 7159 15691
rect 7282 15688 7288 15700
rect 7147 15660 7288 15688
rect 7147 15657 7159 15660
rect 7101 15651 7159 15657
rect 4430 15552 4436 15564
rect 4391 15524 4436 15552
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 4246 15444 4252 15496
rect 4304 15484 4310 15496
rect 4525 15487 4583 15493
rect 4525 15484 4537 15487
rect 4304 15456 4537 15484
rect 4304 15444 4310 15456
rect 4525 15453 4537 15456
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 6656 15484 6684 15651
rect 7282 15648 7288 15660
rect 7340 15688 7346 15700
rect 7558 15688 7564 15700
rect 7340 15660 7564 15688
rect 7340 15648 7346 15660
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 8846 15688 8852 15700
rect 7708 15660 7753 15688
rect 8807 15660 8852 15688
rect 7708 15648 7714 15660
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 10597 15691 10655 15697
rect 10597 15657 10609 15691
rect 10643 15688 10655 15691
rect 10870 15688 10876 15700
rect 10643 15660 10876 15688
rect 10643 15657 10655 15660
rect 10597 15651 10655 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11793 15623 11851 15629
rect 11793 15589 11805 15623
rect 11839 15620 11851 15623
rect 12253 15623 12311 15629
rect 12253 15620 12265 15623
rect 11839 15592 12265 15620
rect 11839 15589 11851 15592
rect 11793 15583 11851 15589
rect 12253 15589 12265 15592
rect 12299 15620 12311 15623
rect 12342 15620 12348 15632
rect 12299 15592 12348 15620
rect 12299 15589 12311 15592
rect 12253 15583 12311 15589
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 7558 15552 7564 15564
rect 7519 15524 7564 15552
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 8846 15552 8852 15564
rect 8444 15524 8852 15552
rect 8444 15512 8450 15524
rect 8846 15512 8852 15524
rect 8904 15512 8910 15564
rect 7742 15484 7748 15496
rect 4672 15456 4765 15484
rect 6656 15456 7748 15484
rect 4672 15444 4678 15456
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 9677 15487 9735 15493
rect 9677 15484 9689 15487
rect 9640 15456 9689 15484
rect 9640 15444 9646 15456
rect 9677 15453 9689 15456
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 12308 15456 12357 15484
rect 12308 15444 12314 15456
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 12575 15456 13032 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 4632 15416 4660 15444
rect 4120 15388 4660 15416
rect 12360 15416 12388 15447
rect 12894 15416 12900 15428
rect 12360 15388 12900 15416
rect 4120 15376 4126 15388
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 13004 15360 13032 15456
rect 5166 15348 5172 15360
rect 5127 15320 5172 15348
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 7190 15348 7196 15360
rect 7151 15320 7196 15348
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11882 15348 11888 15360
rect 11843 15320 11888 15348
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 12986 15348 12992 15360
rect 12947 15320 12992 15348
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 3421 15147 3479 15153
rect 3421 15113 3433 15147
rect 3467 15144 3479 15147
rect 3605 15147 3663 15153
rect 3605 15144 3617 15147
rect 3467 15116 3617 15144
rect 3467 15113 3479 15116
rect 3421 15107 3479 15113
rect 3605 15113 3617 15116
rect 3651 15144 3663 15147
rect 4246 15144 4252 15156
rect 3651 15116 4252 15144
rect 3651 15113 3663 15116
rect 3605 15107 3663 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15144 7895 15147
rect 7926 15144 7932 15156
rect 7883 15116 7932 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 10686 15104 10692 15156
rect 10744 15144 10750 15156
rect 10781 15147 10839 15153
rect 10781 15144 10793 15147
rect 10744 15116 10793 15144
rect 10744 15104 10750 15116
rect 10781 15113 10793 15116
rect 10827 15113 10839 15147
rect 12158 15144 12164 15156
rect 12119 15116 12164 15144
rect 10781 15107 10839 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 12710 15144 12716 15156
rect 12268 15116 12716 15144
rect 3973 15079 4031 15085
rect 3973 15045 3985 15079
rect 4019 15076 4031 15079
rect 4062 15076 4068 15088
rect 4019 15048 4068 15076
rect 4019 15045 4031 15048
rect 3973 15039 4031 15045
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 6273 15079 6331 15085
rect 6273 15045 6285 15079
rect 6319 15076 6331 15079
rect 6319 15048 7420 15076
rect 6319 15045 6331 15048
rect 6273 15039 6331 15045
rect 7392 15020 7420 15048
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11793 15079 11851 15085
rect 11793 15076 11805 15079
rect 11204 15048 11805 15076
rect 11204 15036 11210 15048
rect 11793 15045 11805 15048
rect 11839 15076 11851 15079
rect 12268 15076 12296 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 12952 15116 13461 15144
rect 12952 15104 12958 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 11839 15048 12296 15076
rect 11839 15045 11851 15048
rect 11793 15039 11851 15045
rect 5166 14968 5172 15020
rect 5224 15008 5230 15020
rect 5353 15011 5411 15017
rect 5353 15008 5365 15011
rect 5224 14980 5365 15008
rect 5224 14968 5230 14980
rect 5353 14977 5365 14980
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 7190 15008 7196 15020
rect 5951 14980 7196 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 8444 14980 8585 15008
rect 8444 14968 8450 14980
rect 8573 14977 8585 14980
rect 8619 15008 8631 15011
rect 9306 15008 9312 15020
rect 8619 14980 9312 15008
rect 8619 14977 8631 14980
rect 8573 14971 8631 14977
rect 9306 14968 9312 14980
rect 9364 15008 9370 15020
rect 9585 15011 9643 15017
rect 9585 15008 9597 15011
rect 9364 14980 9597 15008
rect 9364 14968 9370 14980
rect 9585 14977 9597 14980
rect 9631 14977 9643 15011
rect 9585 14971 9643 14977
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 15008 10747 15011
rect 10870 15008 10876 15020
rect 10735 14980 10876 15008
rect 10735 14977 10747 14980
rect 10689 14971 10747 14977
rect 10870 14968 10876 14980
rect 10928 15008 10934 15020
rect 11425 15011 11483 15017
rect 11425 15008 11437 15011
rect 10928 14980 11437 15008
rect 10928 14968 10934 14980
rect 11425 14977 11437 14980
rect 11471 15008 11483 15011
rect 11974 15008 11980 15020
rect 11471 14980 11980 15008
rect 11471 14977 11483 14980
rect 11425 14971 11483 14977
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12986 15008 12992 15020
rect 12492 14980 12992 15008
rect 12492 14968 12498 14980
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 7208 14940 7236 14968
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 4387 14912 5396 14940
rect 7208 14912 7297 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 3237 14875 3295 14881
rect 3237 14841 3249 14875
rect 3283 14872 3295 14875
rect 4430 14872 4436 14884
rect 3283 14844 4436 14872
rect 3283 14841 3295 14844
rect 3237 14835 3295 14841
rect 4430 14832 4436 14844
rect 4488 14832 4494 14884
rect 4614 14872 4620 14884
rect 4575 14844 4620 14872
rect 4614 14832 4620 14844
rect 4672 14872 4678 14884
rect 5261 14875 5319 14881
rect 5261 14872 5273 14875
rect 4672 14844 5273 14872
rect 4672 14832 4678 14844
rect 5261 14841 5273 14844
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 5368 14816 5396 14912
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14940 8999 14943
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 8987 14912 9505 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 9493 14909 9505 14912
rect 9539 14940 9551 14943
rect 9674 14940 9680 14952
rect 9539 14912 9680 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 9674 14900 9680 14912
rect 9732 14940 9738 14952
rect 10410 14940 10416 14952
rect 9732 14912 10416 14940
rect 9732 14900 9738 14912
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 11238 14940 11244 14952
rect 11195 14912 11244 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 11238 14900 11244 14912
rect 11296 14940 11302 14952
rect 11882 14940 11888 14952
rect 11296 14912 11888 14940
rect 11296 14900 11302 14912
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 12158 14900 12164 14952
rect 12216 14940 12222 14952
rect 12216 14912 12848 14940
rect 12216 14900 12222 14912
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 9401 14875 9459 14881
rect 6687 14844 7052 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7024 14816 7052 14844
rect 9401 14841 9413 14875
rect 9447 14872 9459 14875
rect 9582 14872 9588 14884
rect 9447 14844 9588 14872
rect 9447 14841 9459 14844
rect 9401 14835 9459 14841
rect 9582 14832 9588 14844
rect 9640 14832 9646 14884
rect 12820 14881 12848 14912
rect 12805 14875 12863 14881
rect 11256 14844 12480 14872
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 3421 14807 3479 14813
rect 3421 14804 3433 14807
rect 2740 14776 3433 14804
rect 2740 14764 2746 14776
rect 3421 14773 3433 14776
rect 3467 14773 3479 14807
rect 4798 14804 4804 14816
rect 4759 14776 4804 14804
rect 3421 14767 3479 14773
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5169 14807 5227 14813
rect 5169 14773 5181 14807
rect 5215 14804 5227 14807
rect 5350 14804 5356 14816
rect 5215 14776 5356 14804
rect 5215 14773 5227 14776
rect 5169 14767 5227 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 7064 14776 7205 14804
rect 7064 14764 7070 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 9033 14807 9091 14813
rect 9033 14773 9045 14807
rect 9079 14804 9091 14807
rect 9306 14804 9312 14816
rect 9079 14776 9312 14804
rect 9079 14773 9091 14776
rect 9033 14767 9091 14773
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 10318 14804 10324 14816
rect 10279 14776 10324 14804
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 11256 14813 11284 14844
rect 12452 14813 12480 14844
rect 12805 14841 12817 14875
rect 12851 14872 12863 14875
rect 13722 14872 13728 14884
rect 12851 14844 13728 14872
rect 12851 14841 12863 14844
rect 12805 14835 12863 14841
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 11112 14776 11253 14804
rect 11112 14764 11118 14776
rect 11241 14773 11253 14776
rect 11287 14773 11299 14807
rect 11241 14767 11299 14773
rect 12437 14807 12495 14813
rect 12437 14773 12449 14807
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12768 14776 12909 14804
rect 12768 14764 12774 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 4249 14603 4307 14609
rect 4249 14569 4261 14603
rect 4295 14600 4307 14603
rect 4430 14600 4436 14612
rect 4295 14572 4436 14600
rect 4295 14569 4307 14572
rect 4249 14563 4307 14569
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4709 14603 4767 14609
rect 4709 14569 4721 14603
rect 4755 14600 4767 14603
rect 4798 14600 4804 14612
rect 4755 14572 4804 14600
rect 4755 14569 4767 14572
rect 4709 14563 4767 14569
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6822 14600 6828 14612
rect 6595 14572 6828 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7285 14603 7343 14609
rect 7285 14569 7297 14603
rect 7331 14600 7343 14603
rect 7558 14600 7564 14612
rect 7331 14572 7564 14600
rect 7331 14569 7343 14572
rect 7285 14563 7343 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 7653 14603 7711 14609
rect 7653 14569 7665 14603
rect 7699 14600 7711 14603
rect 7742 14600 7748 14612
rect 7699 14572 7748 14600
rect 7699 14569 7711 14572
rect 7653 14563 7711 14569
rect 7742 14560 7748 14572
rect 7800 14560 7806 14612
rect 8021 14603 8079 14609
rect 8021 14569 8033 14603
rect 8067 14600 8079 14603
rect 8202 14600 8208 14612
rect 8067 14572 8208 14600
rect 8067 14569 8079 14572
rect 8021 14563 8079 14569
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 9125 14603 9183 14609
rect 9125 14569 9137 14603
rect 9171 14600 9183 14603
rect 9582 14600 9588 14612
rect 9171 14572 9588 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 10229 14603 10287 14609
rect 10229 14569 10241 14603
rect 10275 14600 10287 14603
rect 10778 14600 10784 14612
rect 10275 14572 10784 14600
rect 10275 14569 10287 14572
rect 10229 14563 10287 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11238 14600 11244 14612
rect 11199 14572 11244 14600
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 13173 14603 13231 14609
rect 13173 14600 13185 14603
rect 12032 14572 13185 14600
rect 12032 14560 12038 14572
rect 13173 14569 13185 14572
rect 13219 14569 13231 14603
rect 13173 14563 13231 14569
rect 6638 14532 6644 14544
rect 6599 14504 6644 14532
rect 6638 14492 6644 14504
rect 6696 14492 6702 14544
rect 12060 14535 12118 14541
rect 12060 14501 12072 14535
rect 12106 14532 12118 14535
rect 12158 14532 12164 14544
rect 12106 14504 12164 14532
rect 12106 14501 12118 14504
rect 12060 14495 12118 14501
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 4982 14464 4988 14476
rect 4663 14436 4988 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 9306 14464 9312 14476
rect 8435 14436 9312 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 10597 14467 10655 14473
rect 10597 14464 10609 14467
rect 10376 14436 10609 14464
rect 10376 14424 10382 14436
rect 10597 14433 10609 14436
rect 10643 14464 10655 14467
rect 10962 14464 10968 14476
rect 10643 14436 10968 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 4801 14399 4859 14405
rect 4801 14396 4813 14399
rect 4764 14368 4813 14396
rect 4764 14356 4770 14368
rect 4801 14365 4813 14368
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 6788 14368 6833 14396
rect 6788 14356 6794 14368
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 7926 14396 7932 14408
rect 7616 14368 7932 14396
rect 7616 14356 7622 14368
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8478 14396 8484 14408
rect 8439 14368 8484 14396
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 8754 14396 8760 14408
rect 8711 14368 8760 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 10410 14396 10416 14408
rect 10183 14368 10416 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10410 14356 10416 14368
rect 10468 14396 10474 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10468 14368 10701 14396
rect 10468 14356 10474 14368
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 10870 14396 10876 14408
rect 10831 14368 10876 14396
rect 10689 14359 10747 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 11790 14396 11796 14408
rect 11480 14368 11796 14396
rect 11480 14356 11486 14368
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 7466 14288 7472 14340
rect 7524 14328 7530 14340
rect 7650 14328 7656 14340
rect 7524 14300 7656 14328
rect 7524 14288 7530 14300
rect 7650 14288 7656 14300
rect 7708 14288 7714 14340
rect 3053 14263 3111 14269
rect 3053 14229 3065 14263
rect 3099 14260 3111 14263
rect 3326 14260 3332 14272
rect 3099 14232 3332 14260
rect 3099 14229 3111 14232
rect 3053 14223 3111 14229
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5684 14232 6193 14260
rect 5684 14220 5690 14232
rect 6181 14229 6193 14232
rect 6227 14229 6239 14263
rect 6181 14223 6239 14229
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12158 14260 12164 14272
rect 11747 14232 12164 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12158 14220 12164 14232
rect 12216 14260 12222 14272
rect 12434 14260 12440 14272
rect 12216 14232 12440 14260
rect 12216 14220 12222 14232
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 6822 14056 6828 14068
rect 5951 14028 6828 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8202 14056 8208 14068
rect 8076 14028 8208 14056
rect 8076 14016 8082 14028
rect 8202 14016 8208 14028
rect 8260 14056 8266 14068
rect 8754 14056 8760 14068
rect 8260 14028 8760 14056
rect 8260 14016 8266 14028
rect 8754 14016 8760 14028
rect 8812 14056 8818 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 8812 14028 9229 14056
rect 8812 14016 8818 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 10410 14056 10416 14068
rect 10371 14028 10416 14056
rect 9217 14019 9275 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11974 14056 11980 14068
rect 11563 14028 11980 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12161 14059 12219 14065
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 12434 14056 12440 14068
rect 12207 14028 12440 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 4341 13991 4399 13997
rect 4341 13957 4353 13991
rect 4387 13988 4399 13991
rect 5166 13988 5172 14000
rect 4387 13960 5172 13988
rect 4387 13957 4399 13960
rect 4341 13951 4399 13957
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 6638 13988 6644 14000
rect 6599 13960 6644 13988
rect 6638 13948 6644 13960
rect 6696 13948 6702 14000
rect 10321 13991 10379 13997
rect 10321 13957 10333 13991
rect 10367 13988 10379 13991
rect 10594 13988 10600 14000
rect 10367 13960 10600 13988
rect 10367 13957 10379 13960
rect 10321 13951 10379 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 9953 13923 10011 13929
rect 7423 13892 7972 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7944 13864 7972 13892
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 9999 13892 11069 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 11057 13889 11069 13892
rect 11103 13920 11115 13923
rect 12176 13920 12204 14019
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 11103 13892 12204 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 2314 13812 2320 13864
rect 2372 13852 2378 13864
rect 2869 13855 2927 13861
rect 2869 13852 2881 13855
rect 2372 13824 2881 13852
rect 2372 13812 2378 13824
rect 2869 13821 2881 13824
rect 2915 13852 2927 13855
rect 2961 13855 3019 13861
rect 2961 13852 2973 13855
rect 2915 13824 2973 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 2961 13821 2973 13824
rect 3007 13852 3019 13855
rect 4982 13852 4988 13864
rect 3007 13824 4844 13852
rect 4943 13824 4988 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3228 13787 3286 13793
rect 3228 13753 3240 13787
rect 3274 13784 3286 13787
rect 3326 13784 3332 13796
rect 3274 13756 3332 13784
rect 3274 13753 3286 13756
rect 3228 13747 3286 13753
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 4816 13784 4844 13824
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 5534 13852 5540 13864
rect 5399 13824 5540 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 6273 13855 6331 13861
rect 6273 13821 6285 13855
rect 6319 13852 6331 13855
rect 6730 13852 6736 13864
rect 6319 13824 6736 13852
rect 6319 13821 6331 13824
rect 6273 13815 6331 13821
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 4890 13784 4896 13796
rect 4816 13756 4896 13784
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 7098 13744 7104 13796
rect 7156 13784 7162 13796
rect 7745 13787 7803 13793
rect 7745 13784 7757 13787
rect 7156 13756 7757 13784
rect 7156 13744 7162 13756
rect 7745 13753 7757 13756
rect 7791 13784 7803 13787
rect 7852 13784 7880 13815
rect 7926 13812 7932 13864
rect 7984 13852 7990 13864
rect 8104 13855 8162 13861
rect 8104 13852 8116 13855
rect 7984 13824 8116 13852
rect 7984 13812 7990 13824
rect 8104 13821 8116 13824
rect 8150 13852 8162 13855
rect 8386 13852 8392 13864
rect 8150 13824 8392 13852
rect 8150 13821 8162 13824
rect 8104 13815 8162 13821
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 10594 13812 10600 13864
rect 10652 13852 10658 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10652 13824 10793 13852
rect 10652 13812 10658 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 11790 13852 11796 13864
rect 10781 13815 10839 13821
rect 10980 13824 11796 13852
rect 10980 13796 11008 13824
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 10962 13784 10968 13796
rect 7791 13756 10968 13784
rect 7791 13753 7803 13756
rect 7745 13747 7803 13753
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 12342 13744 12348 13796
rect 12400 13784 12406 13796
rect 12437 13787 12495 13793
rect 12437 13784 12449 13787
rect 12400 13756 12449 13784
rect 12400 13744 12406 13756
rect 12437 13753 12449 13756
rect 12483 13753 12495 13787
rect 12437 13747 12495 13753
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 10928 13688 10973 13716
rect 10928 13676 10934 13688
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2682 13512 2688 13524
rect 2455 13484 2688 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 4709 13515 4767 13521
rect 4709 13481 4721 13515
rect 4755 13512 4767 13515
rect 4798 13512 4804 13524
rect 4755 13484 4804 13512
rect 4755 13481 4767 13484
rect 4709 13475 4767 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 7926 13512 7932 13524
rect 7887 13484 7932 13512
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 8021 13515 8079 13521
rect 8021 13481 8033 13515
rect 8067 13512 8079 13515
rect 8478 13512 8484 13524
rect 8067 13484 8484 13512
rect 8067 13481 8079 13484
rect 8021 13475 8079 13481
rect 8478 13472 8484 13484
rect 8536 13512 8542 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8536 13484 9045 13512
rect 8536 13472 8542 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 9364 13484 9413 13512
rect 9364 13472 9370 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 9401 13475 9459 13481
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10870 13512 10876 13524
rect 10183 13484 10876 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10870 13472 10876 13484
rect 10928 13512 10934 13524
rect 11149 13515 11207 13521
rect 11149 13512 11161 13515
rect 10928 13484 11161 13512
rect 10928 13472 10934 13484
rect 11149 13481 11161 13484
rect 11195 13481 11207 13515
rect 12066 13512 12072 13524
rect 12027 13484 12072 13512
rect 11149 13475 11207 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 1762 13404 1768 13456
rect 1820 13444 1826 13456
rect 2869 13447 2927 13453
rect 2869 13444 2881 13447
rect 1820 13416 2881 13444
rect 1820 13404 1826 13416
rect 2869 13413 2881 13416
rect 2915 13444 2927 13447
rect 4246 13444 4252 13456
rect 2915 13416 4252 13444
rect 2915 13413 2927 13416
rect 2869 13407 2927 13413
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 5166 13453 5172 13456
rect 5160 13444 5172 13453
rect 5127 13416 5172 13444
rect 5160 13407 5172 13416
rect 5166 13404 5172 13407
rect 5224 13404 5230 13456
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 8202 13444 8208 13456
rect 7607 13416 8208 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13376 2835 13379
rect 3050 13376 3056 13388
rect 2823 13348 3056 13376
rect 2823 13345 2835 13348
rect 2777 13339 2835 13345
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 8018 13376 8024 13388
rect 6972 13348 8024 13376
rect 6972 13336 6978 13348
rect 8018 13336 8024 13348
rect 8076 13376 8082 13388
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 8076 13348 8401 13376
rect 8076 13336 8082 13348
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 10284 13348 10517 13376
rect 10284 13336 10290 13348
rect 10505 13345 10517 13348
rect 10551 13376 10563 13379
rect 10778 13376 10784 13388
rect 10551 13348 10784 13376
rect 10551 13345 10563 13348
rect 10505 13339 10563 13345
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 2590 13268 2596 13320
rect 2648 13308 2654 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2648 13280 2973 13308
rect 2648 13268 2654 13280
rect 2961 13277 2973 13280
rect 3007 13308 3019 13311
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 3007 13280 4261 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 4249 13277 4261 13280
rect 4295 13308 4307 13311
rect 4706 13308 4712 13320
rect 4295 13280 4712 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4890 13308 4896 13320
rect 4851 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 8478 13308 8484 13320
rect 8439 13280 8484 13308
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 4724 13172 4752 13268
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 8588 13240 8616 13271
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 10376 13280 10609 13308
rect 10376 13268 10382 13280
rect 10597 13277 10609 13280
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 8444 13212 8616 13240
rect 10045 13243 10103 13249
rect 8444 13200 8450 13212
rect 10045 13209 10057 13243
rect 10091 13240 10103 13243
rect 10502 13240 10508 13252
rect 10091 13212 10508 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 10502 13200 10508 13212
rect 10560 13240 10566 13252
rect 10704 13240 10732 13271
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11882 13308 11888 13320
rect 11572 13280 11888 13308
rect 11572 13268 11578 13280
rect 11882 13268 11888 13280
rect 11940 13308 11946 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 11940 13280 12173 13308
rect 11940 13268 11946 13280
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13308 12403 13311
rect 12434 13308 12440 13320
rect 12391 13280 12440 13308
rect 12391 13277 12403 13280
rect 12345 13271 12403 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 10560 13212 10732 13240
rect 10560 13200 10566 13212
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 11701 13243 11759 13249
rect 11701 13240 11713 13243
rect 11112 13212 11713 13240
rect 11112 13200 11118 13212
rect 11701 13209 11713 13212
rect 11747 13209 11759 13243
rect 11701 13203 11759 13209
rect 6273 13175 6331 13181
rect 6273 13172 6285 13175
rect 4724 13144 6285 13172
rect 6273 13141 6285 13144
rect 6319 13141 6331 13175
rect 6914 13172 6920 13184
rect 6875 13144 6920 13172
rect 6273 13135 6331 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 1762 12968 1768 12980
rect 1723 12940 1768 12968
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 4338 12928 4344 12980
rect 4396 12968 4402 12980
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 4396 12940 4629 12968
rect 4396 12928 4402 12940
rect 4617 12937 4629 12940
rect 4663 12968 4675 12971
rect 5166 12968 5172 12980
rect 4663 12940 5172 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 7374 12968 7380 12980
rect 6319 12940 7380 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 8478 12968 8484 12980
rect 8391 12940 8484 12968
rect 8478 12928 8484 12940
rect 8536 12968 8542 12980
rect 9858 12968 9864 12980
rect 8536 12940 9864 12968
rect 8536 12928 8542 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10502 12968 10508 12980
rect 10463 12940 10508 12968
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11572 12940 11805 12968
rect 11572 12928 11578 12940
rect 11793 12937 11805 12940
rect 11839 12968 11851 12971
rect 12066 12968 12072 12980
rect 11839 12940 12072 12968
rect 11839 12937 11851 12940
rect 11793 12931 11851 12937
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 12492 12940 12633 12968
rect 12492 12928 12498 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 12621 12931 12679 12937
rect 6822 12900 6828 12912
rect 6783 12872 6828 12900
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 5626 12832 5632 12844
rect 4295 12804 5632 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5810 12832 5816 12844
rect 5771 12804 5816 12832
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 7392 12841 7420 12928
rect 8036 12900 8064 12928
rect 8386 12900 8392 12912
rect 8036 12872 8392 12900
rect 8386 12860 8392 12872
rect 8444 12860 8450 12912
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 11882 12832 11888 12844
rect 10744 12804 11888 12832
rect 10744 12792 10750 12804
rect 11882 12792 11888 12804
rect 11940 12832 11946 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 11940 12804 12081 12832
rect 11940 12792 11946 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 2133 12767 2191 12773
rect 2133 12733 2145 12767
rect 2179 12764 2191 12767
rect 2225 12767 2283 12773
rect 2225 12764 2237 12767
rect 2179 12736 2237 12764
rect 2179 12733 2191 12736
rect 2133 12727 2191 12733
rect 2225 12733 2237 12736
rect 2271 12764 2283 12767
rect 2314 12764 2320 12776
rect 2271 12736 2320 12764
rect 2271 12733 2283 12736
rect 2225 12727 2283 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 5534 12764 5540 12776
rect 5495 12736 5540 12764
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7190 12764 7196 12776
rect 6972 12736 7196 12764
rect 6972 12724 6978 12736
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12764 9091 12767
rect 9125 12767 9183 12773
rect 9125 12764 9137 12767
rect 9079 12736 9137 12764
rect 9079 12733 9091 12736
rect 9033 12727 9091 12733
rect 9125 12733 9137 12736
rect 9171 12733 9183 12767
rect 9125 12727 9183 12733
rect 2498 12705 2504 12708
rect 2492 12696 2504 12705
rect 2459 12668 2504 12696
rect 2492 12659 2504 12668
rect 2498 12656 2504 12659
rect 2556 12656 2562 12708
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 4985 12699 5043 12705
rect 4985 12696 4997 12699
rect 4948 12668 4997 12696
rect 4948 12656 4954 12668
rect 4985 12665 4997 12668
rect 5031 12696 5043 12699
rect 5031 12668 5304 12696
rect 5031 12665 5043 12668
rect 4985 12659 5043 12665
rect 2866 12588 2872 12640
rect 2924 12628 2930 12640
rect 3326 12628 3332 12640
rect 2924 12600 3332 12628
rect 2924 12588 2930 12600
rect 3326 12588 3332 12600
rect 3384 12628 3390 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3384 12600 3617 12628
rect 3384 12588 3390 12600
rect 3605 12597 3617 12600
rect 3651 12597 3663 12631
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 3605 12591 3663 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 5276 12628 5304 12668
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 6086 12696 6092 12708
rect 5684 12668 6092 12696
rect 5684 12656 5690 12668
rect 6086 12656 6092 12668
rect 6144 12696 6150 12708
rect 6549 12699 6607 12705
rect 6549 12696 6561 12699
rect 6144 12668 6561 12696
rect 6144 12656 6150 12668
rect 6549 12665 6561 12668
rect 6595 12696 6607 12699
rect 7285 12699 7343 12705
rect 7285 12696 7297 12699
rect 6595 12668 7297 12696
rect 6595 12665 6607 12668
rect 6549 12659 6607 12665
rect 7285 12665 7297 12668
rect 7331 12665 7343 12699
rect 7285 12659 7343 12665
rect 7098 12628 7104 12640
rect 5276 12600 7104 12628
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 9140 12628 9168 12727
rect 9306 12656 9312 12708
rect 9364 12705 9370 12708
rect 9364 12699 9428 12705
rect 9364 12665 9382 12699
rect 9416 12665 9428 12699
rect 9364 12659 9428 12665
rect 9364 12656 9370 12659
rect 9674 12628 9680 12640
rect 9140 12600 9680 12628
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 10778 12588 10784 12640
rect 10836 12628 10842 12640
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 10836 12600 11161 12628
rect 10836 12588 10842 12600
rect 11149 12597 11161 12600
rect 11195 12628 11207 12631
rect 12066 12628 12072 12640
rect 11195 12600 12072 12628
rect 11195 12597 11207 12600
rect 11149 12591 11207 12597
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 1670 12424 1676 12436
rect 1631 12396 1676 12424
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 2590 12424 2596 12436
rect 2551 12396 2596 12424
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 5534 12424 5540 12436
rect 5495 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 5994 12424 6000 12436
rect 5868 12396 6000 12424
rect 5868 12384 5874 12396
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 6914 12424 6920 12436
rect 6827 12396 6920 12424
rect 6914 12384 6920 12396
rect 6972 12424 6978 12436
rect 7098 12424 7104 12436
rect 6972 12396 7104 12424
rect 6972 12384 6978 12396
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 8478 12424 8484 12436
rect 8391 12396 8484 12424
rect 8478 12384 8484 12396
rect 8536 12424 8542 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 8536 12396 9229 12424
rect 8536 12384 8542 12396
rect 9217 12393 9229 12396
rect 9263 12424 9275 12427
rect 9306 12424 9312 12436
rect 9263 12396 9312 12424
rect 9263 12393 9275 12396
rect 9217 12387 9275 12393
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 10318 12424 10324 12436
rect 10275 12396 10324 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 10962 12424 10968 12436
rect 10428 12396 10968 12424
rect 5261 12359 5319 12365
rect 5261 12325 5273 12359
rect 5307 12356 5319 12359
rect 5442 12356 5448 12368
rect 5307 12328 5448 12356
rect 5307 12325 5319 12328
rect 5261 12319 5319 12325
rect 5442 12316 5448 12328
rect 5500 12316 5506 12368
rect 5905 12359 5963 12365
rect 5905 12325 5917 12359
rect 5951 12356 5963 12359
rect 6178 12356 6184 12368
rect 5951 12328 6184 12356
rect 5951 12325 5963 12328
rect 5905 12319 5963 12325
rect 6178 12316 6184 12328
rect 6236 12356 6242 12368
rect 6822 12356 6828 12368
rect 6236 12328 6828 12356
rect 6236 12316 6242 12328
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 5166 12288 5172 12300
rect 4939 12260 5172 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 5166 12248 5172 12260
rect 5224 12288 5230 12300
rect 5350 12288 5356 12300
rect 5224 12260 5356 12288
rect 5224 12248 5230 12260
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 7116 12297 7144 12384
rect 7368 12359 7426 12365
rect 7368 12356 7380 12359
rect 7208 12328 7380 12356
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12257 7159 12291
rect 7101 12251 7159 12257
rect 5994 12220 6000 12232
rect 5955 12192 6000 12220
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 6144 12192 6193 12220
rect 6144 12180 6150 12192
rect 6181 12189 6193 12192
rect 6227 12220 6239 12223
rect 6730 12220 6736 12232
rect 6227 12192 6736 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6730 12180 6736 12192
rect 6788 12220 6794 12232
rect 7208 12220 7236 12328
rect 7368 12325 7380 12328
rect 7414 12356 7426 12359
rect 7466 12356 7472 12368
rect 7414 12328 7472 12356
rect 7414 12325 7426 12328
rect 7368 12319 7426 12325
rect 7466 12316 7472 12328
rect 7524 12316 7530 12368
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10428 12356 10456 12396
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 12434 12424 12440 12436
rect 11931 12396 12440 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 9732 12328 10456 12356
rect 9732 12316 9738 12328
rect 9766 12248 9772 12300
rect 9824 12288 9830 12300
rect 10134 12288 10140 12300
rect 9824 12260 10140 12288
rect 9824 12248 9830 12260
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10428 12220 10456 12328
rect 10502 12316 10508 12368
rect 10560 12316 10566 12368
rect 10520 12288 10548 12316
rect 10778 12297 10784 12300
rect 10772 12288 10784 12297
rect 10520 12260 10784 12288
rect 10772 12251 10784 12260
rect 10778 12248 10784 12251
rect 10836 12248 10842 12300
rect 10502 12220 10508 12232
rect 6788 12192 7236 12220
rect 10415 12192 10508 12220
rect 6788 12180 6794 12192
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 2317 12155 2375 12161
rect 2317 12121 2329 12155
rect 2363 12152 2375 12155
rect 2498 12152 2504 12164
rect 2363 12124 2504 12152
rect 2363 12121 2375 12124
rect 2317 12115 2375 12121
rect 2498 12112 2504 12124
rect 2556 12152 2562 12164
rect 3510 12152 3516 12164
rect 2556 12124 3516 12152
rect 2556 12112 2562 12124
rect 3510 12112 3516 12124
rect 3568 12112 3574 12164
rect 3050 12084 3056 12096
rect 3011 12056 3056 12084
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 10410 12084 10416 12096
rect 5316 12056 10416 12084
rect 5316 12044 5322 12056
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3697 11883 3755 11889
rect 3697 11880 3709 11883
rect 3568 11852 3709 11880
rect 3568 11840 3574 11852
rect 3697 11849 3709 11852
rect 3743 11849 3755 11883
rect 3697 11843 3755 11849
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 4304 11852 4813 11880
rect 4304 11840 4310 11852
rect 4801 11849 4813 11852
rect 4847 11849 4859 11883
rect 4801 11843 4859 11849
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6086 11880 6092 11892
rect 5951 11852 6092 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 10502 11880 10508 11892
rect 10463 11852 10508 11880
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 10836 11852 10885 11880
rect 10836 11840 10842 11852
rect 10873 11849 10885 11852
rect 10919 11849 10931 11883
rect 10873 11843 10931 11849
rect 4338 11812 4344 11824
rect 4299 11784 4344 11812
rect 4338 11772 4344 11784
rect 4396 11812 4402 11824
rect 4396 11784 5396 11812
rect 4396 11772 4402 11784
rect 5368 11756 5396 11784
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2314 11744 2320 11756
rect 2271 11716 2320 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 5350 11744 5356 11756
rect 5263 11716 5356 11744
rect 5350 11704 5356 11716
rect 5408 11704 5414 11756
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 6822 11744 6828 11756
rect 6687 11716 6828 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 5166 11676 5172 11688
rect 5127 11648 5172 11676
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11676 5319 11679
rect 5442 11676 5448 11688
rect 5307 11648 5448 11676
rect 5307 11645 5319 11648
rect 5261 11639 5319 11645
rect 2038 11568 2044 11620
rect 2096 11608 2102 11620
rect 2562 11611 2620 11617
rect 2562 11608 2574 11611
rect 2096 11580 2574 11608
rect 2096 11568 2102 11580
rect 2562 11577 2574 11580
rect 2608 11577 2620 11611
rect 2562 11571 2620 11577
rect 4709 11611 4767 11617
rect 4709 11577 4721 11611
rect 4755 11608 4767 11611
rect 5074 11608 5080 11620
rect 4755 11580 5080 11608
rect 4755 11577 4767 11580
rect 4709 11571 4767 11577
rect 5074 11568 5080 11580
rect 5132 11608 5138 11620
rect 5276 11608 5304 11639
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6273 11679 6331 11685
rect 6273 11676 6285 11679
rect 6144 11648 6285 11676
rect 6144 11636 6150 11648
rect 6273 11645 6285 11648
rect 6319 11676 6331 11679
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6319 11648 7093 11676
rect 6319 11645 6331 11648
rect 6273 11639 6331 11645
rect 7081 11645 7093 11648
rect 7127 11676 7139 11679
rect 7374 11676 7380 11688
rect 7127 11648 7380 11676
rect 7127 11645 7139 11648
rect 7081 11639 7139 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 10686 11608 10692 11620
rect 5132 11580 5304 11608
rect 7208 11580 10692 11608
rect 5132 11568 5138 11580
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 7208 11540 7236 11580
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 5500 11512 7236 11540
rect 5500 11500 5506 11512
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7524 11512 8217 11540
rect 7524 11500 7530 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 4801 11339 4859 11345
rect 4801 11336 4813 11339
rect 3108 11308 4813 11336
rect 3108 11296 3114 11308
rect 4801 11305 4813 11308
rect 4847 11305 4859 11339
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 4801 11299 4859 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 5905 11339 5963 11345
rect 5905 11305 5917 11339
rect 5951 11336 5963 11339
rect 5994 11336 6000 11348
rect 5951 11308 6000 11336
rect 5951 11305 5963 11308
rect 5905 11299 5963 11305
rect 5994 11296 6000 11308
rect 6052 11336 6058 11348
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 6052 11308 6377 11336
rect 6052 11296 6058 11308
rect 6365 11305 6377 11308
rect 6411 11305 6423 11339
rect 6365 11299 6423 11305
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7248 11308 7941 11336
rect 7248 11296 7254 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 4982 11228 4988 11280
rect 5040 11268 5046 11280
rect 5169 11271 5227 11277
rect 5169 11268 5181 11271
rect 5040 11240 5181 11268
rect 5040 11228 5046 11240
rect 5169 11237 5181 11240
rect 5215 11268 5227 11271
rect 5442 11268 5448 11280
rect 5215 11240 5448 11268
rect 5215 11237 5227 11240
rect 5169 11231 5227 11237
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 6178 11268 6184 11280
rect 6139 11240 6184 11268
rect 6178 11228 6184 11240
rect 6236 11228 6242 11280
rect 7466 11268 7472 11280
rect 7427 11240 7472 11268
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 6454 11200 6460 11212
rect 5868 11172 6460 11200
rect 5868 11160 5874 11172
rect 6454 11160 6460 11172
rect 6512 11200 6518 11212
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 6512 11172 6745 11200
rect 6512 11160 6518 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 6733 11163 6791 11169
rect 5350 11132 5356 11144
rect 5311 11104 5356 11132
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7374 11132 7380 11144
rect 7055 11104 7380 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 1854 10996 1860 11008
rect 1815 10968 1860 10996
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 2038 10956 2044 11008
rect 2096 10996 2102 11008
rect 2317 10999 2375 11005
rect 2317 10996 2329 10999
rect 2096 10968 2329 10996
rect 2096 10956 2102 10968
rect 2317 10965 2329 10968
rect 2363 10965 2375 10999
rect 3418 10996 3424 11008
rect 3379 10968 3424 10996
rect 2317 10959 2375 10965
rect 3418 10956 3424 10968
rect 3476 10956 3482 11008
rect 6840 10996 6868 11095
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7006 10996 7012 11008
rect 6840 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10996 7070 11008
rect 8110 10996 8116 11008
rect 7064 10968 8116 10996
rect 7064 10956 7070 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 12526 10996 12532 11008
rect 12487 10968 12532 10996
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 3237 10795 3295 10801
rect 3237 10761 3249 10795
rect 3283 10792 3295 10795
rect 3510 10792 3516 10804
rect 3283 10764 3516 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 3510 10752 3516 10764
rect 3568 10752 3574 10804
rect 4893 10795 4951 10801
rect 4893 10761 4905 10795
rect 4939 10792 4951 10795
rect 5258 10792 5264 10804
rect 4939 10764 5264 10792
rect 4939 10761 4951 10764
rect 4893 10755 4951 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 6086 10792 6092 10804
rect 6047 10764 6092 10792
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 3329 10727 3387 10733
rect 3329 10693 3341 10727
rect 3375 10693 3387 10727
rect 3528 10724 3556 10752
rect 3528 10696 3924 10724
rect 3329 10687 3387 10693
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2317 10659 2375 10665
rect 2317 10656 2329 10659
rect 1719 10628 2329 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2317 10625 2329 10628
rect 2363 10656 2375 10659
rect 2866 10656 2872 10668
rect 2363 10628 2872 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 1854 10548 1860 10600
rect 1912 10588 1918 10600
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1912 10560 2145 10588
rect 1912 10548 1918 10560
rect 2133 10557 2145 10560
rect 2179 10588 2191 10591
rect 3344 10588 3372 10687
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 3896 10665 3924 10696
rect 4982 10684 4988 10736
rect 5040 10724 5046 10736
rect 5169 10727 5227 10733
rect 5169 10724 5181 10727
rect 5040 10696 5181 10724
rect 5040 10684 5046 10696
rect 5169 10693 5181 10696
rect 5215 10693 5227 10727
rect 5169 10687 5227 10693
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3476 10628 3801 10656
rect 3476 10616 3482 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10625 3939 10659
rect 3881 10619 3939 10625
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12986 10656 12992 10668
rect 12584 10628 12992 10656
rect 12584 10616 12590 10628
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 2179 10560 3372 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 3694 10520 3700 10532
rect 2915 10492 3700 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3694 10480 3700 10492
rect 3752 10480 3758 10532
rect 6454 10520 6460 10532
rect 6415 10492 6460 10520
rect 6454 10480 6460 10492
rect 6512 10480 6518 10532
rect 12250 10520 12256 10532
rect 12163 10492 12256 10520
rect 12250 10480 12256 10492
rect 12308 10520 12314 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12308 10492 12817 10520
rect 12308 10480 12314 10492
rect 12805 10489 12817 10492
rect 12851 10520 12863 10523
rect 14090 10520 14096 10532
rect 12851 10492 14096 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 2225 10455 2283 10461
rect 2225 10421 2237 10455
rect 2271 10452 2283 10455
rect 2406 10452 2412 10464
rect 2271 10424 2412 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 4430 10452 4436 10464
rect 4391 10424 4436 10452
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 7006 10452 7012 10464
rect 6967 10424 7012 10452
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7745 10455 7803 10461
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 8018 10452 8024 10464
rect 7791 10424 8024 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12526 10452 12532 10464
rect 12483 10424 12532 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12894 10452 12900 10464
rect 12855 10424 12900 10452
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2406 10248 2412 10260
rect 1903 10220 2412 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 3752 10220 4353 10248
rect 3752 10208 3758 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 8110 10248 8116 10260
rect 8071 10220 8116 10248
rect 4341 10211 4399 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12894 10248 12900 10260
rect 12575 10220 12900 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 2777 10183 2835 10189
rect 2777 10149 2789 10183
rect 2823 10180 2835 10183
rect 2866 10180 2872 10192
rect 2823 10152 2872 10180
rect 2823 10149 2835 10152
rect 2777 10143 2835 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 4706 10112 4712 10124
rect 4667 10084 4712 10112
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5626 10112 5632 10124
rect 4816 10084 5632 10112
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2406 10044 2412 10056
rect 2363 10016 2412 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2406 10004 2412 10016
rect 2464 10044 2470 10056
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2464 10016 2881 10044
rect 2464 10004 2470 10016
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3510 10044 3516 10056
rect 3099 10016 3516 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 3068 9976 3096 10007
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4246 10004 4252 10056
rect 4304 10044 4310 10056
rect 4816 10053 4844 10084
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7926 10112 7932 10124
rect 7340 10084 7932 10112
rect 7340 10072 7346 10084
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8478 10112 8484 10124
rect 8067 10084 8484 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 10413 10115 10471 10121
rect 10413 10081 10425 10115
rect 10459 10112 10471 10115
rect 10502 10112 10508 10124
rect 10459 10084 10508 10112
rect 10459 10081 10471 10084
rect 10413 10075 10471 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10686 10121 10692 10124
rect 10680 10112 10692 10121
rect 10647 10084 10692 10112
rect 10680 10075 10692 10084
rect 10686 10072 10692 10075
rect 10744 10072 10750 10124
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10112 13415 10115
rect 13630 10112 13636 10124
rect 13403 10084 13636 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 4801 10047 4859 10053
rect 4801 10044 4813 10047
rect 4304 10016 4813 10044
rect 4304 10004 4310 10016
rect 4801 10013 4813 10016
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 13446 10044 13452 10056
rect 13407 10016 13452 10044
rect 8205 10007 8263 10013
rect 2832 9948 3096 9976
rect 2832 9936 2838 9948
rect 4430 9936 4436 9988
rect 4488 9976 4494 9988
rect 4908 9976 4936 10007
rect 4488 9948 4936 9976
rect 4488 9936 4494 9948
rect 8018 9936 8024 9988
rect 8076 9976 8082 9988
rect 8220 9976 8248 10007
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 8076 9948 8248 9976
rect 12897 9979 12955 9985
rect 8076 9936 8082 9948
rect 12897 9945 12909 9979
rect 12943 9976 12955 9979
rect 13538 9976 13544 9988
rect 12943 9948 13544 9976
rect 12943 9945 12955 9948
rect 12897 9939 12955 9945
rect 13538 9936 13544 9948
rect 13596 9936 13602 9988
rect 7374 9908 7380 9920
rect 7335 9880 7380 9908
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 7524 9880 7665 9908
rect 7524 9868 7530 9880
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 8941 9911 8999 9917
rect 8941 9877 8953 9911
rect 8987 9908 8999 9911
rect 9306 9908 9312 9920
rect 8987 9880 9312 9908
rect 8987 9877 8999 9880
rect 8941 9871 8999 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 11793 9911 11851 9917
rect 11793 9877 11805 9911
rect 11839 9908 11851 9911
rect 11974 9908 11980 9920
rect 11839 9880 11980 9908
rect 11839 9877 11851 9880
rect 11793 9871 11851 9877
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 3476 9676 4108 9704
rect 3476 9664 3482 9676
rect 1578 9636 1584 9648
rect 1539 9608 1584 9636
rect 1578 9596 1584 9608
rect 1636 9596 1642 9648
rect 4080 9636 4108 9676
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4580 9676 4936 9704
rect 4580 9664 4586 9676
rect 4433 9639 4491 9645
rect 4433 9636 4445 9639
rect 4080 9608 4445 9636
rect 4433 9605 4445 9608
rect 4479 9605 4491 9639
rect 4433 9599 4491 9605
rect 4908 9636 4936 9676
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10778 9704 10784 9716
rect 10560 9676 10784 9704
rect 10560 9664 10566 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 13262 9704 13268 9716
rect 12483 9676 13268 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 5261 9639 5319 9645
rect 4908 9608 5120 9636
rect 2038 9568 2044 9580
rect 1951 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9568 2102 9580
rect 3050 9568 3056 9580
rect 2096 9540 3056 9568
rect 2096 9528 2102 9540
rect 3050 9528 3056 9540
rect 3108 9568 3114 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 3108 9540 3525 9568
rect 3108 9528 3114 9540
rect 3513 9537 3525 9540
rect 3559 9568 3571 9571
rect 4908 9568 4936 9608
rect 5092 9577 5120 9608
rect 5261 9605 5273 9639
rect 5307 9636 5319 9639
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5307 9608 5825 9636
rect 5307 9605 5319 9608
rect 5261 9599 5319 9605
rect 5813 9605 5825 9608
rect 5859 9605 5871 9639
rect 5813 9599 5871 9605
rect 11885 9639 11943 9645
rect 11885 9605 11897 9639
rect 11931 9636 11943 9639
rect 12526 9636 12532 9648
rect 11931 9608 12532 9636
rect 11931 9605 11943 9608
rect 11885 9599 11943 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 3559 9540 4936 9568
rect 5077 9571 5135 9577
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 5077 9537 5089 9571
rect 5123 9568 5135 9571
rect 5534 9568 5540 9580
rect 5123 9540 5540 9568
rect 5123 9537 5135 9540
rect 5077 9531 5135 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 7929 9571 7987 9577
rect 7929 9537 7941 9571
rect 7975 9568 7987 9571
rect 8018 9568 8024 9580
rect 7975 9540 8024 9568
rect 7975 9537 7987 9540
rect 7929 9531 7987 9537
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 12032 9540 12265 9568
rect 12032 9528 12038 9540
rect 12253 9537 12265 9540
rect 12299 9568 12311 9571
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12299 9540 13001 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13320 9540 14197 9568
rect 13320 9528 13326 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1762 9500 1768 9512
rect 1443 9472 1768 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 2372 9472 2421 9500
rect 2372 9460 2378 9472
rect 2409 9469 2421 9472
rect 2455 9500 2467 9503
rect 2455 9472 3372 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 3344 9444 3372 9472
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3476 9472 3985 9500
rect 3476 9460 3482 9472
rect 3973 9469 3985 9472
rect 4019 9500 4031 9503
rect 4246 9500 4252 9512
rect 4019 9472 4252 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4387 9472 4813 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 4801 9469 4813 9472
rect 4847 9500 4859 9503
rect 5810 9500 5816 9512
rect 4847 9472 5816 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 7432 9472 7665 9500
rect 7432 9460 7438 9472
rect 7653 9469 7665 9472
rect 7699 9469 7711 9503
rect 8754 9500 8760 9512
rect 8667 9472 8760 9500
rect 7653 9463 7711 9469
rect 8754 9460 8760 9472
rect 8812 9500 8818 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8812 9472 8861 9500
rect 8812 9460 8818 9472
rect 8849 9469 8861 9472
rect 8895 9500 8907 9503
rect 10502 9500 10508 9512
rect 8895 9472 10508 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 10502 9460 10508 9472
rect 10560 9460 10566 9512
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9500 11391 9503
rect 12434 9500 12440 9512
rect 11379 9472 12440 9500
rect 11379 9469 11391 9472
rect 11333 9463 11391 9469
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 12802 9500 12808 9512
rect 12715 9472 12808 9500
rect 12802 9460 12808 9472
rect 12860 9500 12866 9512
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 12860 9472 13829 9500
rect 12860 9460 12866 9472
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 3326 9432 3332 9444
rect 3287 9404 3332 9432
rect 3326 9392 3332 9404
rect 3384 9392 3390 9444
rect 4430 9392 4436 9444
rect 4488 9432 4494 9444
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4488 9404 4905 9432
rect 4488 9392 4494 9404
rect 4893 9401 4905 9404
rect 4939 9432 4951 9435
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 4939 9404 5457 9432
rect 4939 9401 4951 9404
rect 4893 9395 4951 9401
rect 5445 9401 5457 9404
rect 5491 9432 5503 9435
rect 5718 9432 5724 9444
rect 5491 9404 5724 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 7193 9435 7251 9441
rect 7193 9401 7205 9435
rect 7239 9432 7251 9435
rect 8389 9435 8447 9441
rect 7239 9404 7788 9432
rect 7239 9401 7251 9404
rect 7193 9395 7251 9401
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 2823 9336 3249 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3237 9333 3249 9336
rect 3283 9364 3295 9367
rect 3510 9364 3516 9376
rect 3283 9336 3516 9364
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 4764 9336 5273 9364
rect 4764 9324 4770 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 5261 9327 5319 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5592 9336 6193 9364
rect 5592 9324 5598 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6638 9364 6644 9376
rect 6599 9336 6644 9364
rect 6181 9327 6239 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7760 9373 7788 9404
rect 8389 9401 8401 9435
rect 8435 9432 8447 9435
rect 8478 9432 8484 9444
rect 8435 9404 8484 9432
rect 8435 9401 8447 9404
rect 8389 9395 8447 9401
rect 8478 9392 8484 9404
rect 8536 9432 8542 9444
rect 9116 9435 9174 9441
rect 8536 9404 9076 9432
rect 8536 9392 8542 9404
rect 7745 9367 7803 9373
rect 7745 9333 7757 9367
rect 7791 9364 7803 9367
rect 8294 9364 8300 9376
rect 7791 9336 8300 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 8294 9324 8300 9336
rect 8352 9364 8358 9376
rect 8570 9364 8576 9376
rect 8352 9336 8576 9364
rect 8352 9324 8358 9336
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 9048 9364 9076 9404
rect 9116 9401 9128 9435
rect 9162 9432 9174 9435
rect 9306 9432 9312 9444
rect 9162 9404 9312 9432
rect 9162 9401 9174 9404
rect 9116 9395 9174 9401
rect 9306 9392 9312 9404
rect 9364 9432 9370 9444
rect 10042 9432 10048 9444
rect 9364 9404 10048 9432
rect 9364 9392 9370 9404
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10686 9432 10692 9444
rect 10244 9404 10692 9432
rect 10244 9376 10272 9404
rect 10686 9392 10692 9404
rect 10744 9432 10750 9444
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 10744 9404 11161 9432
rect 10744 9392 10750 9404
rect 11149 9401 11161 9404
rect 11195 9401 11207 9435
rect 11149 9395 11207 9401
rect 9490 9364 9496 9376
rect 9048 9336 9496 9364
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10226 9364 10232 9376
rect 10187 9336 10232 9364
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12584 9336 12909 9364
rect 12584 9324 12590 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 12897 9327 12955 9333
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 5534 9160 5540 9172
rect 5491 9132 5540 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7374 9160 7380 9172
rect 7055 9132 7380 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 8067 9132 10609 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 10597 9129 10609 9132
rect 10643 9160 10655 9163
rect 10962 9160 10968 9172
rect 10643 9132 10968 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12676 9132 13093 9160
rect 12676 9120 12682 9132
rect 13081 9129 13093 9132
rect 13127 9160 13139 9163
rect 13446 9160 13452 9172
rect 13127 9132 13452 9160
rect 13127 9129 13139 9132
rect 13081 9123 13139 9129
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 13630 9160 13636 9172
rect 13591 9132 13636 9160
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 2866 9092 2872 9104
rect 1995 9064 2872 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 4522 9092 4528 9104
rect 4080 9064 4528 9092
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 9024 2375 9027
rect 2682 9024 2688 9036
rect 2363 8996 2688 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 4080 9033 4108 9064
rect 4522 9052 4528 9064
rect 4580 9052 4586 9104
rect 5994 9052 6000 9104
rect 6052 9092 6058 9104
rect 7745 9095 7803 9101
rect 7745 9092 7757 9095
rect 6052 9064 7757 9092
rect 6052 9052 6058 9064
rect 7745 9061 7757 9064
rect 7791 9092 7803 9095
rect 8110 9092 8116 9104
rect 7791 9064 8116 9092
rect 7791 9061 7803 9064
rect 7745 9055 7803 9061
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 11974 9101 11980 9104
rect 11968 9055 11980 9101
rect 12032 9092 12038 9104
rect 12032 9064 12068 9092
rect 11974 9052 11980 9055
rect 12032 9052 12038 9064
rect 4338 9033 4344 9036
rect 4065 9027 4123 9033
rect 2832 8996 2877 9024
rect 2832 8984 2838 8996
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4332 9024 4344 9033
rect 4299 8996 4344 9024
rect 4065 8987 4123 8993
rect 4332 8987 4344 8996
rect 4338 8984 4344 8987
rect 4396 8984 4402 9036
rect 8386 9024 8392 9036
rect 8347 8996 8392 9024
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 10502 9024 10508 9036
rect 10463 8996 10508 9024
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8352 8928 8493 8956
rect 8352 8916 8358 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 10226 8956 10232 8968
rect 8619 8928 10232 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 8588 8888 8616 8919
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10686 8956 10692 8968
rect 10647 8928 10692 8956
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 11698 8956 11704 8968
rect 10836 8928 11704 8956
rect 10836 8916 10842 8928
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 13630 8888 13636 8900
rect 8260 8860 8616 8888
rect 13004 8860 13636 8888
rect 8260 8848 8266 8860
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 9582 8820 9588 8832
rect 3568 8792 9588 8820
rect 3568 8780 3574 8792
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 10137 8823 10195 8829
rect 10137 8789 10149 8823
rect 10183 8820 10195 8823
rect 13004 8820 13032 8860
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 10183 8792 13032 8820
rect 10183 8789 10195 8792
rect 10137 8783 10195 8789
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8616 1731 8619
rect 1762 8616 1768 8628
rect 1719 8588 1768 8616
rect 1719 8585 1731 8588
rect 1673 8579 1731 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2501 8619 2559 8625
rect 2501 8585 2513 8619
rect 2547 8616 2559 8619
rect 2774 8616 2780 8628
rect 2547 8588 2780 8616
rect 2547 8585 2559 8588
rect 2501 8579 2559 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 2924 8588 3341 8616
rect 2924 8576 2930 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3329 8579 3387 8585
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 7282 8616 7288 8628
rect 6319 8588 7288 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8904 8588 9045 8616
rect 8904 8576 8910 8588
rect 9033 8585 9045 8588
rect 9079 8616 9091 8619
rect 10962 8616 10968 8628
rect 9079 8588 9996 8616
rect 10923 8588 10968 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 9585 8551 9643 8557
rect 9585 8548 9597 8551
rect 8352 8520 9597 8548
rect 8352 8508 8358 8520
rect 9585 8517 9597 8520
rect 9631 8517 9643 8551
rect 9585 8511 9643 8517
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3988 8412 4016 8443
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4764 8452 4905 8480
rect 4764 8440 4770 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 4338 8412 4344 8424
rect 2915 8384 4344 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 4338 8372 4344 8384
rect 4396 8412 4402 8424
rect 4396 8384 4752 8412
rect 4396 8372 4402 8384
rect 4724 8356 4752 8384
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6972 8384 7113 8412
rect 6972 8372 6978 8384
rect 7101 8381 7113 8384
rect 7147 8412 7159 8415
rect 8754 8412 8760 8424
rect 7147 8384 8760 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 9968 8421 9996 8588
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 11974 8576 11980 8628
rect 12032 8616 12038 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12032 8588 12173 8616
rect 12032 8576 12038 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 12437 8619 12495 8625
rect 12437 8585 12449 8619
rect 12483 8616 12495 8619
rect 12802 8616 12808 8628
rect 12483 8588 12808 8616
rect 12483 8585 12495 8588
rect 12437 8579 12495 8585
rect 10686 8548 10692 8560
rect 10599 8520 10692 8548
rect 10686 8508 10692 8520
rect 10744 8548 10750 8560
rect 11425 8551 11483 8557
rect 11425 8548 11437 8551
rect 10744 8520 11437 8548
rect 10744 8508 10750 8520
rect 11425 8517 11437 8520
rect 11471 8548 11483 8551
rect 11882 8548 11888 8560
rect 11471 8520 11888 8548
rect 11471 8517 11483 8520
rect 11425 8511 11483 8517
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10137 8483 10195 8489
rect 10137 8480 10149 8483
rect 10100 8452 10149 8480
rect 10100 8440 10106 8452
rect 10137 8449 10149 8452
rect 10183 8449 10195 8483
rect 12176 8480 12204 8579
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12176 8452 12909 8480
rect 10137 8443 10195 8449
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13044 8452 13089 8480
rect 13044 8440 13050 8452
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8381 10011 8415
rect 9953 8375 10011 8381
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12492 8384 12817 8412
rect 12492 8372 12498 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 3697 8347 3755 8353
rect 3697 8313 3709 8347
rect 3743 8344 3755 8347
rect 4062 8344 4068 8356
rect 3743 8316 4068 8344
rect 3743 8313 3755 8316
rect 3697 8307 3755 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4706 8344 4712 8356
rect 4667 8316 4712 8344
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 6638 8344 6644 8356
rect 6551 8316 6644 8344
rect 6638 8304 6644 8316
rect 6696 8344 6702 8356
rect 7368 8347 7426 8353
rect 7368 8344 7380 8347
rect 6696 8316 7380 8344
rect 6696 8304 6702 8316
rect 7368 8313 7380 8316
rect 7414 8344 7426 8347
rect 8018 8344 8024 8356
rect 7414 8316 8024 8344
rect 7414 8313 7426 8316
rect 7368 8307 7426 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 9401 8347 9459 8353
rect 9401 8344 9413 8347
rect 9364 8316 9413 8344
rect 9364 8304 9370 8316
rect 9401 8313 9413 8316
rect 9447 8344 9459 8347
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 9447 8316 10057 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 10045 8313 10057 8316
rect 10091 8344 10103 8347
rect 10134 8344 10140 8356
rect 10091 8316 10140 8344
rect 10091 8313 10103 8316
rect 10045 8307 10103 8313
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 3237 8279 3295 8285
rect 3237 8245 3249 8279
rect 3283 8276 3295 8279
rect 3786 8276 3792 8288
rect 3283 8248 3792 8276
rect 3283 8245 3295 8248
rect 3237 8239 3295 8245
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4522 8276 4528 8288
rect 4479 8248 4528 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 8481 8279 8539 8285
rect 8481 8276 8493 8279
rect 7708 8248 8493 8276
rect 7708 8236 7714 8248
rect 8481 8245 8493 8248
rect 8527 8245 8539 8279
rect 8481 8239 8539 8245
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2866 8072 2872 8084
rect 2547 8044 2872 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 6972 8044 7113 8072
rect 6972 8032 6978 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 7101 8035 7159 8041
rect 8021 8075 8079 8081
rect 8021 8041 8033 8075
rect 8067 8072 8079 8075
rect 8386 8072 8392 8084
rect 8067 8044 8392 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 8386 8032 8392 8044
rect 8444 8072 8450 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8444 8044 9045 8072
rect 8444 8032 8450 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 10321 8075 10379 8081
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 10413 8075 10471 8081
rect 10413 8072 10425 8075
rect 10367 8044 10425 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10413 8041 10425 8044
rect 10459 8072 10471 8075
rect 10502 8072 10508 8084
rect 10459 8044 10508 8072
rect 10459 8041 10471 8044
rect 10413 8035 10471 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12897 8075 12955 8081
rect 12492 8044 12537 8072
rect 12492 8032 12498 8044
rect 12897 8041 12909 8075
rect 12943 8072 12955 8075
rect 12986 8072 12992 8084
rect 12943 8044 12992 8072
rect 12943 8041 12955 8044
rect 12897 8035 12955 8041
rect 7561 8007 7619 8013
rect 7561 7973 7573 8007
rect 7607 8004 7619 8007
rect 8294 8004 8300 8016
rect 7607 7976 8300 8004
rect 7607 7973 7619 7976
rect 7561 7967 7619 7973
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 10226 7964 10232 8016
rect 10284 8004 10290 8016
rect 12912 8004 12940 8035
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 10284 7976 12940 8004
rect 10284 7964 10290 7976
rect 5436 7939 5494 7945
rect 5436 7905 5448 7939
rect 5482 7936 5494 7939
rect 5810 7936 5816 7948
rect 5482 7908 5816 7936
rect 5482 7905 5494 7908
rect 5436 7899 5494 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 8202 7936 8208 7948
rect 7975 7908 8208 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8386 7936 8392 7948
rect 8347 7908 8392 7936
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10244 7908 10793 7936
rect 10244 7880 10272 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 10980 7880 11008 7976
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 4062 7868 4068 7880
rect 3467 7840 4068 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4580 7840 5181 7868
rect 4580 7828 4586 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5184 7732 5212 7831
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 8168 7840 8493 7868
rect 8168 7828 8174 7840
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 8754 7868 8760 7880
rect 8711 7840 8760 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8754 7828 8760 7840
rect 8812 7868 8818 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 8812 7840 9413 7868
rect 8812 7828 8818 7840
rect 9401 7837 9413 7840
rect 9447 7868 9459 7871
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 9447 7840 9873 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9861 7837 9873 7840
rect 9907 7868 9919 7871
rect 10042 7868 10048 7880
rect 9907 7840 10048 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 10870 7868 10876 7880
rect 10831 7840 10876 7868
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11020 7840 11113 7868
rect 11020 7828 11026 7840
rect 6178 7760 6184 7812
rect 6236 7800 6242 7812
rect 8294 7800 8300 7812
rect 6236 7772 8300 7800
rect 6236 7760 6242 7772
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 5442 7732 5448 7744
rect 5184 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6086 7692 6092 7744
rect 6144 7732 6150 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 6144 7704 6561 7732
rect 6144 7692 6150 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6549 7695 6607 7701
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 9674 7732 9680 7744
rect 9456 7704 9680 7732
rect 9456 7692 9462 7704
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 5074 7488 5080 7500
rect 5132 7528 5138 7540
rect 5626 7528 5632 7540
rect 5132 7500 5632 7528
rect 5132 7488 5138 7500
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 8110 7488 8116 7500
rect 8168 7528 8174 7540
rect 8386 7528 8392 7540
rect 8168 7500 8248 7528
rect 8347 7500 8392 7528
rect 8168 7488 8174 7500
rect 2038 7420 2044 7472
rect 2096 7460 2102 7472
rect 6178 7460 6184 7472
rect 2096 7432 6184 7460
rect 2096 7420 2102 7432
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 6730 7460 6736 7472
rect 6687 7432 6736 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 6730 7420 6736 7432
rect 6788 7460 6794 7472
rect 8220 7460 8248 7500
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 9309 7531 9367 7537
rect 9309 7497 9321 7531
rect 9355 7528 9367 7531
rect 9674 7528 9680 7540
rect 9355 7500 9680 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 10781 7531 10839 7537
rect 10781 7497 10793 7531
rect 10827 7528 10839 7531
rect 10962 7528 10968 7540
rect 10827 7500 10968 7528
rect 10827 7497 10839 7500
rect 10781 7491 10839 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 15746 7528 15752 7540
rect 13872 7500 15752 7528
rect 13872 7488 13878 7500
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 8662 7460 8668 7472
rect 6788 7432 7696 7460
rect 8220 7432 8668 7460
rect 6788 7420 6794 7432
rect 7668 7404 7696 7432
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 9401 7463 9459 7469
rect 9401 7429 9413 7463
rect 9447 7460 9459 7463
rect 10870 7460 10876 7472
rect 9447 7432 10876 7460
rect 9447 7429 9459 7432
rect 9401 7423 9459 7429
rect 10870 7420 10876 7432
rect 10928 7460 10934 7472
rect 11149 7463 11207 7469
rect 11149 7460 11161 7463
rect 10928 7432 11161 7460
rect 10928 7420 10934 7432
rect 11149 7429 11161 7432
rect 11195 7429 11207 7463
rect 11149 7423 11207 7429
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 5810 7392 5816 7404
rect 4387 7364 5816 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 5810 7352 5816 7364
rect 5868 7392 5874 7404
rect 5868 7364 6316 7392
rect 5868 7352 5874 7364
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1443 7296 1992 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1964 7200 1992 7296
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 5224 7296 5549 7324
rect 5224 7284 5230 7296
rect 5537 7293 5549 7296
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 5684 7296 5729 7324
rect 5684 7284 5690 7296
rect 4709 7259 4767 7265
rect 4709 7225 4721 7259
rect 4755 7256 4767 7259
rect 5442 7256 5448 7268
rect 4755 7228 5448 7256
rect 4755 7225 4767 7228
rect 4709 7219 4767 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 6288 7265 6316 7364
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7466 7392 7472 7404
rect 6880 7364 7472 7392
rect 6880 7352 6886 7364
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 10042 7392 10048 7404
rect 10003 7364 10048 7392
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 7282 7284 7288 7336
rect 7340 7324 7346 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 7340 7296 7389 7324
rect 7340 7284 7346 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 8754 7324 8760 7336
rect 8715 7296 8760 7324
rect 7377 7287 7435 7293
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 6273 7259 6331 7265
rect 6273 7225 6285 7259
rect 6319 7256 6331 7259
rect 6638 7256 6644 7268
rect 6319 7228 6644 7256
rect 6319 7225 6331 7228
rect 6273 7219 6331 7225
rect 6638 7216 6644 7228
rect 6696 7216 6702 7268
rect 9769 7259 9827 7265
rect 9769 7225 9781 7259
rect 9815 7256 9827 7259
rect 9950 7256 9956 7268
rect 9815 7228 9956 7256
rect 9815 7225 9827 7228
rect 9769 7219 9827 7225
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7009 7191 7067 7197
rect 7009 7188 7021 7191
rect 6972 7160 7021 7188
rect 6972 7148 6978 7160
rect 7009 7157 7021 7160
rect 7055 7157 7067 7191
rect 7009 7151 7067 7157
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 9861 7191 9919 7197
rect 9861 7188 9873 7191
rect 9732 7160 9873 7188
rect 9732 7148 9738 7160
rect 9861 7157 9873 7160
rect 9907 7188 9919 7191
rect 10042 7188 10048 7200
rect 9907 7160 10048 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10226 7148 10232 7200
rect 10284 7188 10290 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10284 7160 10425 7188
rect 10284 7148 10290 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 5132 6956 5181 6984
rect 5132 6944 5138 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 5169 6947 5227 6953
rect 6638 6944 6644 6996
rect 6696 6984 6702 6996
rect 7009 6987 7067 6993
rect 7009 6984 7021 6987
rect 6696 6956 7021 6984
rect 6696 6944 6702 6956
rect 7009 6953 7021 6956
rect 7055 6953 7067 6987
rect 7009 6947 7067 6953
rect 6086 6916 6092 6928
rect 5460 6888 6092 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6817 1455 6851
rect 2406 6848 2412 6860
rect 2367 6820 2412 6848
rect 1397 6811 1455 6817
rect 1412 6780 1440 6811
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 5350 6848 5356 6860
rect 4939 6820 5356 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5350 6808 5356 6820
rect 5408 6848 5414 6860
rect 5460 6848 5488 6888
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 9950 6916 9956 6928
rect 9600 6888 9956 6916
rect 5408 6820 5488 6848
rect 5629 6851 5687 6857
rect 5408 6808 5414 6820
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 5718 6848 5724 6860
rect 5675 6820 5724 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 1412 6752 2360 6780
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1544 6616 1593 6644
rect 1544 6604 1550 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1581 6607 1639 6613
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2332 6653 2360 6752
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 5644 6780 5672 6811
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5896 6851 5954 6857
rect 5896 6817 5908 6851
rect 5942 6848 5954 6851
rect 6178 6848 6184 6860
rect 5942 6820 6184 6848
rect 5942 6817 5954 6820
rect 5896 6811 5954 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8202 6848 8208 6860
rect 8159 6820 8208 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8202 6808 8208 6820
rect 8260 6848 8266 6860
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 8260 6820 9505 6848
rect 8260 6808 8266 6820
rect 9493 6817 9505 6820
rect 9539 6848 9551 6851
rect 9600 6848 9628 6888
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 9539 6820 9628 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 12032 6820 12081 6848
rect 12032 6808 12038 6820
rect 12069 6817 12081 6820
rect 12115 6817 12127 6851
rect 12069 6811 12127 6817
rect 12336 6851 12394 6857
rect 12336 6817 12348 6851
rect 12382 6848 12394 6851
rect 12618 6848 12624 6860
rect 12382 6820 12624 6848
rect 12382 6817 12394 6820
rect 12336 6811 12394 6817
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 5500 6752 5672 6780
rect 5500 6740 5506 6752
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 2682 6712 2688 6724
rect 2639 6684 2688 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 9033 6715 9091 6721
rect 9033 6712 9045 6715
rect 7984 6684 9045 6712
rect 7984 6672 7990 6684
rect 9033 6681 9045 6684
rect 9079 6681 9091 6715
rect 9033 6675 9091 6681
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 2498 6644 2504 6656
rect 2363 6616 2504 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 7834 6644 7840 6656
rect 7795 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 8386 6644 8392 6656
rect 8343 6616 8392 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8662 6644 8668 6656
rect 8623 6616 8668 6644
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 10042 6644 10048 6656
rect 10003 6616 10048 6644
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 13446 6644 13452 6656
rect 13407 6616 13452 6644
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 3050 6440 3056 6452
rect 3011 6412 3056 6440
rect 3050 6400 3056 6412
rect 3108 6400 3114 6452
rect 6178 6440 6184 6452
rect 6139 6412 6184 6440
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6822 6440 6828 6452
rect 6687 6412 6828 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7098 6440 7104 6452
rect 7059 6412 7104 6440
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 12032 6412 12081 6440
rect 12032 6400 12038 6412
rect 12069 6409 12081 6412
rect 12115 6409 12127 6443
rect 12618 6440 12624 6452
rect 12579 6412 12624 6440
rect 12069 6403 12127 6409
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 9674 6332 9680 6384
rect 9732 6372 9738 6384
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 9732 6344 10057 6372
rect 9732 6332 9738 6344
rect 10045 6341 10057 6344
rect 10091 6341 10103 6375
rect 10045 6335 10103 6341
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 5166 6304 5172 6316
rect 4387 6276 5172 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 5350 6304 5356 6316
rect 5311 6276 5356 6304
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8720 6276 8861 6304
rect 8720 6264 8726 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 10594 6304 10600 6316
rect 9640 6276 10600 6304
rect 9640 6264 9646 6276
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 5184 6236 5212 6264
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5184 6208 5273 6236
rect 5261 6205 5273 6208
rect 5307 6205 5319 6239
rect 5261 6199 5319 6205
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 7156 6208 7205 6236
rect 7156 6196 7162 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 8168 6208 8769 6236
rect 8168 6196 8174 6208
rect 8757 6205 8769 6208
rect 8803 6236 8815 6239
rect 9306 6236 9312 6248
rect 8803 6208 9312 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9824 6208 9873 6236
rect 9824 6196 9830 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 1854 6128 1860 6180
rect 1912 6177 1918 6180
rect 1912 6171 1976 6177
rect 1912 6137 1930 6171
rect 1964 6137 1976 6171
rect 1912 6131 1976 6137
rect 4709 6171 4767 6177
rect 4709 6137 4721 6171
rect 4755 6168 4767 6171
rect 7837 6171 7895 6177
rect 4755 6140 5212 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 1912 6128 1918 6131
rect 4798 6100 4804 6112
rect 4759 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5184 6109 5212 6140
rect 7837 6137 7849 6171
rect 7883 6168 7895 6171
rect 8665 6171 8723 6177
rect 8665 6168 8677 6171
rect 7883 6140 8677 6168
rect 7883 6137 7895 6140
rect 7837 6131 7895 6137
rect 8665 6137 8677 6140
rect 8711 6168 8723 6171
rect 8846 6168 8852 6180
rect 8711 6140 8852 6168
rect 8711 6137 8723 6140
rect 8665 6131 8723 6137
rect 8846 6128 8852 6140
rect 8904 6128 8910 6180
rect 9876 6168 9904 6199
rect 10042 6196 10048 6248
rect 10100 6236 10106 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 10100 6208 10425 6236
rect 10100 6196 10106 6208
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 10134 6168 10140 6180
rect 9876 6140 10140 6168
rect 10134 6128 10140 6140
rect 10192 6168 10198 6180
rect 10505 6171 10563 6177
rect 10505 6168 10517 6171
rect 10192 6140 10517 6168
rect 10192 6128 10198 6140
rect 10505 6137 10517 6140
rect 10551 6137 10563 6171
rect 10505 6131 10563 6137
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5258 6100 5264 6112
rect 5215 6072 5264 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5810 6100 5816 6112
rect 5771 6072 5816 6100
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6100 7435 6103
rect 7650 6100 7656 6112
rect 7423 6072 7656 6100
rect 7423 6069 7435 6072
rect 7377 6063 7435 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 8110 6100 8116 6112
rect 8071 6072 8116 6100
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8294 6100 8300 6112
rect 8255 6072 8300 6100
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9582 6100 9588 6112
rect 9543 6072 9588 6100
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 1670 5856 1676 5908
rect 1728 5896 1734 5908
rect 1949 5899 2007 5905
rect 1949 5896 1961 5899
rect 1728 5868 1961 5896
rect 1728 5856 1734 5868
rect 1949 5865 1961 5868
rect 1995 5865 2007 5899
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 1949 5859 2007 5865
rect 1964 5828 1992 5859
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5258 5896 5264 5908
rect 4948 5868 5264 5896
rect 4948 5856 4954 5868
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 6178 5856 6184 5908
rect 6236 5896 6242 5908
rect 6730 5896 6736 5908
rect 6236 5868 6736 5896
rect 6236 5856 6242 5868
rect 6730 5856 6736 5868
rect 6788 5896 6794 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6788 5868 7297 5896
rect 6788 5856 6794 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 8202 5896 8208 5908
rect 8163 5868 8208 5896
rect 7285 5859 7343 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 8846 5896 8852 5908
rect 8352 5868 8852 5896
rect 8352 5856 8358 5868
rect 8846 5856 8852 5868
rect 8904 5896 8910 5908
rect 9309 5899 9367 5905
rect 9309 5896 9321 5899
rect 8904 5868 9321 5896
rect 8904 5856 8910 5868
rect 9309 5865 9321 5868
rect 9355 5865 9367 5899
rect 9309 5859 9367 5865
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 9640 5868 9873 5896
rect 9640 5856 9646 5868
rect 9861 5865 9873 5868
rect 9907 5865 9919 5899
rect 9861 5859 9919 5865
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 10505 5899 10563 5905
rect 10505 5896 10517 5899
rect 10468 5868 10517 5896
rect 10468 5856 10474 5868
rect 10505 5865 10517 5868
rect 10551 5865 10563 5899
rect 11054 5896 11060 5908
rect 11015 5868 11060 5896
rect 10505 5859 10563 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11974 5896 11980 5908
rect 11624 5868 11980 5896
rect 2590 5828 2596 5840
rect 1964 5800 2596 5828
rect 2590 5788 2596 5800
rect 2648 5788 2654 5840
rect 5074 5828 5080 5840
rect 2884 5800 5080 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 2682 5760 2688 5772
rect 1443 5732 2688 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 2884 5769 2912 5800
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5810 5788 5816 5840
rect 5868 5828 5874 5840
rect 6270 5828 6276 5840
rect 5868 5800 6276 5828
rect 5868 5788 5874 5800
rect 2869 5763 2927 5769
rect 2869 5760 2881 5763
rect 2832 5732 2881 5760
rect 2832 5720 2838 5732
rect 2869 5729 2881 5732
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 3881 5763 3939 5769
rect 3881 5729 3893 5763
rect 3927 5760 3939 5763
rect 4430 5760 4436 5772
rect 3927 5732 4436 5760
rect 3927 5729 3939 5732
rect 3881 5723 3939 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 4798 5760 4804 5772
rect 4540 5732 4804 5760
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3200 5664 3556 5692
rect 3200 5652 3206 5664
rect 2958 5584 2964 5636
rect 3016 5624 3022 5636
rect 3421 5627 3479 5633
rect 3421 5624 3433 5627
rect 3016 5596 3433 5624
rect 3016 5584 3022 5596
rect 3421 5593 3433 5596
rect 3467 5593 3479 5627
rect 3528 5624 3556 5664
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4540 5701 4568 5732
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 5920 5769 5948 5800
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 11624 5772 11652 5868
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 13446 5828 13452 5840
rect 11900 5800 13452 5828
rect 11900 5772 11928 5800
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5729 5963 5763
rect 5905 5723 5963 5729
rect 6172 5763 6230 5769
rect 6172 5729 6184 5763
rect 6218 5760 6230 5763
rect 6638 5760 6644 5772
rect 6218 5732 6644 5760
rect 6218 5729 6230 5732
rect 6172 5723 6230 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 8202 5720 8208 5772
rect 8260 5760 8266 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8260 5732 8401 5760
rect 8260 5720 8266 5732
rect 8389 5729 8401 5732
rect 8435 5760 8447 5763
rect 8570 5760 8576 5772
rect 8435 5732 8576 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10502 5760 10508 5772
rect 10459 5732 10508 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 11606 5760 11612 5772
rect 11519 5732 11612 5760
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 11882 5769 11888 5772
rect 11876 5760 11888 5769
rect 11843 5732 11888 5760
rect 11876 5723 11888 5732
rect 11882 5720 11888 5723
rect 11940 5720 11946 5772
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4212 5664 4537 5692
rect 4212 5652 4218 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4890 5692 4896 5704
rect 4755 5664 4896 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 5442 5692 5448 5704
rect 5403 5664 5448 5692
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 10652 5664 10697 5692
rect 10652 5652 10658 5664
rect 4798 5624 4804 5636
rect 3528 5596 4804 5624
rect 3421 5587 3479 5593
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 1302 5516 1308 5568
rect 1360 5556 1366 5568
rect 1581 5559 1639 5565
rect 1581 5556 1593 5559
rect 1360 5528 1593 5556
rect 1360 5516 1366 5528
rect 1581 5525 1593 5528
rect 1627 5525 1639 5559
rect 3050 5556 3056 5568
rect 3011 5528 3056 5556
rect 1581 5519 1639 5525
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 4065 5559 4123 5565
rect 4065 5556 4077 5559
rect 3200 5528 4077 5556
rect 3200 5516 3206 5528
rect 4065 5525 4077 5528
rect 4111 5525 4123 5559
rect 4065 5519 4123 5525
rect 5813 5559 5871 5565
rect 5813 5525 5825 5559
rect 5859 5556 5871 5559
rect 6638 5556 6644 5568
rect 5859 5528 6644 5556
rect 5859 5525 5871 5528
rect 5813 5519 5871 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8573 5559 8631 5565
rect 8573 5556 8585 5559
rect 8352 5528 8585 5556
rect 8352 5516 8358 5528
rect 8573 5525 8585 5528
rect 8619 5525 8631 5559
rect 8573 5519 8631 5525
rect 8662 5516 8668 5568
rect 8720 5556 8726 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 8720 5528 8953 5556
rect 8720 5516 8726 5528
rect 8941 5525 8953 5528
rect 8987 5525 8999 5559
rect 10042 5556 10048 5568
rect 10003 5528 10048 5556
rect 8941 5519 8999 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 12986 5556 12992 5568
rect 12947 5528 12992 5556
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 2314 5352 2320 5364
rect 2275 5324 2320 5352
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 2774 5352 2780 5364
rect 2735 5324 2780 5352
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4706 5352 4712 5364
rect 4295 5324 4712 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5960 5324 6193 5352
rect 5960 5312 5966 5324
rect 6181 5321 6193 5324
rect 6227 5321 6239 5355
rect 6181 5315 6239 5321
rect 7469 5355 7527 5361
rect 7469 5321 7481 5355
rect 7515 5352 7527 5355
rect 7742 5352 7748 5364
rect 7515 5324 7748 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 2041 5287 2099 5293
rect 2041 5253 2053 5287
rect 2087 5284 2099 5287
rect 2682 5284 2688 5296
rect 2087 5256 2688 5284
rect 2087 5253 2099 5256
rect 2041 5247 2099 5253
rect 2682 5244 2688 5256
rect 2740 5244 2746 5296
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2648 5188 2881 5216
rect 2648 5176 2654 5188
rect 2869 5185 2881 5188
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 6546 5216 6552 5228
rect 5583 5188 6552 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 6546 5176 6552 5188
rect 6604 5216 6610 5228
rect 7374 5216 7380 5228
rect 6604 5188 7380 5216
rect 6604 5176 6610 5188
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2314 5148 2320 5160
rect 1443 5120 2320 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5902 5148 5908 5160
rect 5675 5120 5908 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7484 5148 7512 5315
rect 7742 5312 7748 5324
rect 7800 5312 7806 5364
rect 10137 5355 10195 5361
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 10410 5352 10416 5364
rect 10183 5324 10416 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 7742 5176 7748 5228
rect 7800 5216 7806 5228
rect 7929 5219 7987 5225
rect 7929 5216 7941 5219
rect 7800 5188 7941 5216
rect 7800 5176 7806 5188
rect 7929 5185 7941 5188
rect 7975 5185 7987 5219
rect 7929 5179 7987 5185
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 10152 5216 10180 5315
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 11606 5352 11612 5364
rect 11567 5324 11612 5352
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 9364 5188 10180 5216
rect 9364 5176 9370 5188
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10376 5188 10425 5216
rect 10376 5176 10382 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 6871 5120 7512 5148
rect 8113 5151 8171 5157
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 8202 5148 8208 5160
rect 8159 5120 8208 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 2958 5040 2964 5092
rect 3016 5080 3022 5092
rect 3114 5083 3172 5089
rect 3114 5080 3126 5083
rect 3016 5052 3126 5080
rect 3016 5040 3022 5052
rect 3114 5049 3126 5052
rect 3160 5049 3172 5083
rect 3114 5043 3172 5049
rect 3602 5040 3608 5092
rect 3660 5080 3666 5092
rect 4154 5080 4160 5092
rect 3660 5052 4160 5080
rect 3660 5040 3666 5052
rect 4154 5040 4160 5052
rect 4212 5080 4218 5092
rect 6270 5080 6276 5092
rect 4212 5052 6276 5080
rect 4212 5040 4218 5052
rect 6270 5040 6276 5052
rect 6328 5080 6334 5092
rect 6641 5083 6699 5089
rect 6641 5080 6653 5083
rect 6328 5052 6653 5080
rect 6328 5040 6334 5052
rect 6641 5049 6653 5052
rect 6687 5080 6699 5083
rect 8128 5080 8156 5111
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8358 5083 8416 5089
rect 8358 5080 8370 5083
rect 6687 5052 8156 5080
rect 8220 5052 8370 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 992 4984 1593 5012
rect 992 4972 998 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 4890 5012 4896 5024
rect 4803 4984 4896 5012
rect 1581 4975 1639 4981
rect 4890 4972 4896 4984
rect 4948 5012 4954 5024
rect 5442 5012 5448 5024
rect 4948 4984 5448 5012
rect 4948 4972 4954 4984
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 5810 5012 5816 5024
rect 5771 4984 5816 5012
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7009 5015 7067 5021
rect 7009 5012 7021 5015
rect 6972 4984 7021 5012
rect 6972 4972 6978 4984
rect 7009 4981 7021 4984
rect 7055 4981 7067 5015
rect 7009 4975 7067 4981
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8220 5012 8248 5052
rect 8358 5049 8370 5052
rect 8404 5080 8416 5083
rect 8570 5080 8576 5092
rect 8404 5052 8576 5080
rect 8404 5049 8416 5052
rect 8358 5043 8416 5049
rect 8570 5040 8576 5052
rect 8628 5040 8634 5092
rect 10428 5080 10456 5179
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 10652 5188 11161 5216
rect 10652 5176 10658 5188
rect 11149 5185 11161 5188
rect 11195 5216 11207 5219
rect 11330 5216 11336 5228
rect 11195 5188 11336 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11330 5176 11336 5188
rect 11388 5216 11394 5228
rect 11882 5216 11888 5228
rect 11388 5188 11888 5216
rect 11388 5176 11394 5188
rect 11882 5176 11888 5188
rect 11940 5216 11946 5228
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 11940 5188 11989 5216
rect 11940 5176 11946 5188
rect 11977 5185 11989 5188
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 10962 5148 10968 5160
rect 10923 5120 10968 5148
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11057 5083 11115 5089
rect 11057 5080 11069 5083
rect 10428 5052 11069 5080
rect 11057 5049 11069 5052
rect 11103 5049 11115 5083
rect 11057 5043 11115 5049
rect 9490 5012 9496 5024
rect 7800 4984 8248 5012
rect 9451 4984 9496 5012
rect 7800 4972 7806 4984
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10870 5012 10876 5024
rect 10643 4984 10876 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 2832 4780 2877 4808
rect 2832 4768 2838 4780
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4488 4780 4629 4808
rect 4488 4768 4494 4780
rect 4617 4777 4629 4780
rect 4663 4777 4675 4811
rect 4617 4771 4675 4777
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 5040 4780 5089 4808
rect 5040 4768 5046 4780
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 5077 4771 5135 4777
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 5592 4780 6193 4808
rect 5592 4768 5598 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6638 4808 6644 4820
rect 6599 4780 6644 4808
rect 6181 4771 6239 4777
rect 6638 4768 6644 4780
rect 6696 4808 6702 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 6696 4780 7757 4808
rect 6696 4768 6702 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7892 4780 8125 4808
rect 7892 4768 7898 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 8113 4771 8171 4777
rect 8849 4811 8907 4817
rect 8849 4777 8861 4811
rect 8895 4808 8907 4811
rect 8938 4808 8944 4820
rect 8895 4780 8944 4808
rect 8895 4777 8907 4780
rect 8849 4771 8907 4777
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 9582 4808 9588 4820
rect 9539 4780 9588 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10502 4808 10508 4820
rect 10183 4780 10508 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10870 4808 10876 4820
rect 10831 4780 10876 4808
rect 10870 4768 10876 4780
rect 10928 4808 10934 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 10928 4780 11805 4808
rect 10928 4768 10934 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 12437 4811 12495 4817
rect 12437 4777 12449 4811
rect 12483 4808 12495 4811
rect 12618 4808 12624 4820
rect 12483 4780 12624 4808
rect 12483 4777 12495 4780
rect 12437 4771 12495 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 2869 4743 2927 4749
rect 2869 4740 2881 4743
rect 2792 4712 2881 4740
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 2792 4604 2820 4712
rect 2869 4709 2881 4712
rect 2915 4740 2927 4743
rect 3142 4740 3148 4752
rect 2915 4712 3148 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 3513 4743 3571 4749
rect 3513 4709 3525 4743
rect 3559 4740 3571 4743
rect 3602 4740 3608 4752
rect 3559 4712 3608 4740
rect 3559 4709 3571 4712
rect 3513 4703 3571 4709
rect 2958 4604 2964 4616
rect 1995 4576 2820 4604
rect 2919 4576 2964 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 2590 4496 2596 4548
rect 2648 4536 2654 4548
rect 3528 4536 3556 4703
rect 3602 4700 3608 4712
rect 3660 4700 3666 4752
rect 3881 4743 3939 4749
rect 3881 4709 3893 4743
rect 3927 4740 3939 4743
rect 3970 4740 3976 4752
rect 3927 4712 3976 4740
rect 3927 4709 3939 4712
rect 3881 4703 3939 4709
rect 3970 4700 3976 4712
rect 4028 4700 4034 4752
rect 5721 4743 5779 4749
rect 5721 4709 5733 4743
rect 5767 4740 5779 4743
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 5767 4712 8217 4740
rect 5767 4709 5779 4712
rect 5721 4703 5779 4709
rect 8205 4709 8217 4712
rect 8251 4740 8263 4743
rect 8294 4740 8300 4752
rect 8251 4712 8300 4740
rect 8251 4709 8263 4712
rect 8205 4703 8263 4709
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11425 4743 11483 4749
rect 11425 4740 11437 4743
rect 11388 4712 11437 4740
rect 11388 4700 11394 4712
rect 11425 4709 11437 4712
rect 11471 4709 11483 4743
rect 11425 4703 11483 4709
rect 4890 4632 4896 4684
rect 4948 4672 4954 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4948 4644 4997 4672
rect 4948 4632 4954 4644
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 6822 4672 6828 4684
rect 6595 4644 6828 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7561 4675 7619 4681
rect 7561 4672 7573 4675
rect 7432 4644 7573 4672
rect 7432 4632 7438 4644
rect 7561 4641 7573 4644
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5350 4604 5356 4616
rect 5307 4576 5356 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 2648 4508 3556 4536
rect 4525 4539 4583 4545
rect 2648 4496 2654 4508
rect 4525 4505 4537 4539
rect 4571 4536 4583 4539
rect 4706 4536 4712 4548
rect 4571 4508 4712 4536
rect 4571 4505 4583 4508
rect 4525 4499 4583 4505
rect 4706 4496 4712 4508
rect 4764 4536 4770 4548
rect 5276 4536 5304 4567
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6730 4604 6736 4616
rect 6691 4576 6736 4604
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7576 4604 7604 4635
rect 9674 4632 9680 4684
rect 9732 4672 9738 4684
rect 10042 4672 10048 4684
rect 9732 4644 10048 4672
rect 9732 4632 9738 4644
rect 10042 4632 10048 4644
rect 10100 4672 10106 4684
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 10100 4644 10793 4672
rect 10100 4632 10106 4644
rect 10781 4641 10793 4644
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 12434 4672 12440 4684
rect 12391 4644 12440 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 7576 4576 8309 4604
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 10962 4604 10968 4616
rect 10923 4576 10968 4604
rect 8297 4567 8355 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 12526 4604 12532 4616
rect 12487 4576 12532 4604
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 4764 4508 5304 4536
rect 6089 4539 6147 4545
rect 4764 4496 4770 4508
rect 6089 4505 6101 4539
rect 6135 4536 6147 4539
rect 6638 4536 6644 4548
rect 6135 4508 6644 4536
rect 6135 4505 6147 4508
rect 6089 4499 6147 4505
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 11238 4496 11244 4548
rect 11296 4536 11302 4548
rect 11977 4539 12035 4545
rect 11977 4536 11989 4539
rect 11296 4508 11989 4536
rect 11296 4496 11302 4508
rect 11977 4505 11989 4508
rect 12023 4505 12035 4539
rect 11977 4499 12035 4505
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 6822 4468 6828 4480
rect 2832 4440 6828 4468
rect 2832 4428 2838 4440
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 7374 4468 7380 4480
rect 7331 4440 7380 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 10410 4468 10416 4480
rect 10371 4440 10416 4468
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 12989 4471 13047 4477
rect 12989 4468 13001 4471
rect 12860 4440 13001 4468
rect 12860 4428 12866 4440
rect 12989 4437 13001 4440
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 4157 4267 4215 4273
rect 4157 4264 4169 4267
rect 3016 4236 4169 4264
rect 3016 4224 3022 4236
rect 4157 4233 4169 4236
rect 4203 4233 4215 4267
rect 4157 4227 4215 4233
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 5040 4236 5089 4264
rect 5040 4224 5046 4236
rect 5077 4233 5089 4236
rect 5123 4233 5135 4267
rect 5077 4227 5135 4233
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 5408 4236 5457 4264
rect 5408 4224 5414 4236
rect 5445 4233 5457 4236
rect 5491 4233 5503 4267
rect 5445 4227 5503 4233
rect 6641 4267 6699 4273
rect 6641 4233 6653 4267
rect 6687 4264 6699 4267
rect 6730 4264 6736 4276
rect 6687 4236 6736 4264
rect 6687 4233 6699 4236
rect 6641 4227 6699 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 6822 4224 6828 4276
rect 6880 4264 6886 4276
rect 6880 4236 6925 4264
rect 6880 4224 6886 4236
rect 2590 4128 2596 4140
rect 2551 4100 2596 4128
rect 2590 4088 2596 4100
rect 2648 4128 2654 4140
rect 2777 4131 2835 4137
rect 2777 4128 2789 4131
rect 2648 4100 2789 4128
rect 2648 4088 2654 4100
rect 2777 4097 2789 4100
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 1627 4032 2237 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 2225 4029 2237 4032
rect 2271 4060 2283 4063
rect 5000 4060 5028 4224
rect 7374 4196 7380 4208
rect 6840 4168 7380 4196
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 6840 4128 6868 4168
rect 7374 4156 7380 4168
rect 7432 4196 7438 4208
rect 11514 4196 11520 4208
rect 7432 4168 7512 4196
rect 7432 4156 7438 4168
rect 7282 4128 7288 4140
rect 5500 4100 6868 4128
rect 7243 4100 7288 4128
rect 5500 4088 5506 4100
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7484 4137 7512 4168
rect 8312 4168 8984 4196
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 8018 4088 8024 4140
rect 8076 4128 8082 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 8076 4100 8125 4128
rect 8076 4088 8082 4100
rect 8113 4097 8125 4100
rect 8159 4128 8171 4131
rect 8312 4128 8340 4168
rect 8956 4140 8984 4168
rect 10796 4168 11520 4196
rect 8846 4128 8852 4140
rect 8159 4100 8340 4128
rect 8807 4100 8852 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8996 4100 9045 4128
rect 8996 4088 9002 4100
rect 9033 4097 9045 4100
rect 9079 4128 9091 4131
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9079 4100 9413 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9401 4097 9413 4100
rect 9447 4128 9459 4131
rect 9490 4128 9496 4140
rect 9447 4100 9496 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 9824 4100 10701 4128
rect 9824 4088 9830 4100
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 5626 4060 5632 4072
rect 2271 4032 5028 4060
rect 5587 4032 5632 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 6822 4060 6828 4072
rect 5776 4032 6828 4060
rect 5776 4020 5782 4032
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 6972 4032 8769 4060
rect 6972 4020 6978 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10594 4060 10600 4072
rect 10183 4032 10600 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10594 4020 10600 4032
rect 10652 4060 10658 4072
rect 10796 4060 10824 4168
rect 11514 4156 11520 4168
rect 11572 4156 11578 4208
rect 12342 4196 12348 4208
rect 11992 4168 12348 4196
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 10962 4128 10968 4140
rect 10919 4100 10968 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 10962 4088 10968 4100
rect 11020 4128 11026 4140
rect 11330 4128 11336 4140
rect 11020 4100 11336 4128
rect 11020 4088 11026 4100
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 10652 4032 10824 4060
rect 10652 4020 10658 4032
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11992 4069 12020 4168
rect 12342 4156 12348 4168
rect 12400 4196 12406 4208
rect 12526 4196 12532 4208
rect 12400 4168 12532 4196
rect 12400 4156 12406 4168
rect 12526 4156 12532 4168
rect 12584 4196 12590 4208
rect 12584 4168 13032 4196
rect 12584 4156 12590 4168
rect 12894 4128 12900 4140
rect 12855 4100 12900 4128
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13004 4137 13032 4168
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11112 4032 11621 4060
rect 11112 4020 11118 4032
rect 11609 4029 11621 4032
rect 11655 4060 11667 4063
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11655 4032 11989 4060
rect 11655 4029 11667 4032
rect 11609 4023 11667 4029
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 11977 4023 12035 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12912 4060 12940 4088
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 12912 4032 13461 4060
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 3044 3995 3102 4001
rect 3044 3961 3056 3995
rect 3090 3992 3102 3995
rect 3602 3992 3608 4004
rect 3090 3964 3608 3992
rect 3090 3961 3102 3964
rect 3044 3955 3102 3961
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5040 3964 5856 3992
rect 5040 3952 5046 3964
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1765 3927 1823 3933
rect 1765 3924 1777 3927
rect 1452 3896 1777 3924
rect 1452 3884 1458 3896
rect 1765 3893 1777 3896
rect 1811 3893 1823 3927
rect 1765 3887 1823 3893
rect 4801 3927 4859 3933
rect 4801 3893 4813 3927
rect 4847 3924 4859 3927
rect 4890 3924 4896 3936
rect 4847 3896 4896 3924
rect 4847 3893 4859 3896
rect 4801 3887 4859 3893
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5828 3933 5856 3964
rect 5994 3952 6000 4004
rect 6052 3992 6058 4004
rect 6181 3995 6239 4001
rect 6181 3992 6193 3995
rect 6052 3964 6193 3992
rect 6052 3952 6058 3964
rect 6181 3961 6193 3964
rect 6227 3961 6239 3995
rect 6181 3955 6239 3961
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 8202 3992 8208 4004
rect 7432 3964 8208 3992
rect 7432 3952 7438 3964
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 12820 3992 12848 4020
rect 10244 3964 12848 3992
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3893 5871 3927
rect 7190 3924 7196 3936
rect 7103 3896 7196 3924
rect 5813 3887 5871 3893
rect 7190 3884 7196 3896
rect 7248 3924 7254 3936
rect 7926 3924 7932 3936
rect 7248 3896 7932 3924
rect 7248 3884 7254 3896
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 10244 3933 10272 3964
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8352 3896 8401 3924
rect 8352 3884 8358 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3893 10287 3927
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10229 3887 10287 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11330 3924 11336 3936
rect 11291 3896 11336 3924
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12526 3924 12532 3936
rect 12483 3896 12532 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 2682 3720 2688 3732
rect 1719 3692 2688 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 2958 3720 2964 3732
rect 2823 3692 2964 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 3602 3720 3608 3732
rect 3559 3692 3608 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 3881 3723 3939 3729
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 4706 3720 4712 3732
rect 3927 3692 4712 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 4856 3692 4905 3720
rect 4856 3680 4862 3692
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 4893 3683 4951 3689
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 5994 3720 6000 3732
rect 5684 3692 6000 3720
rect 5684 3680 5690 3692
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 6273 3723 6331 3729
rect 6273 3720 6285 3723
rect 6236 3692 6285 3720
rect 6236 3680 6242 3692
rect 6273 3689 6285 3692
rect 6319 3720 6331 3723
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 6319 3692 6837 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 7466 3720 7472 3732
rect 7427 3692 7472 3720
rect 6825 3683 6883 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 8021 3723 8079 3729
rect 8021 3720 8033 3723
rect 7892 3692 8033 3720
rect 7892 3680 7898 3692
rect 8021 3689 8033 3692
rect 8067 3689 8079 3723
rect 8021 3683 8079 3689
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 8478 3720 8484 3732
rect 8435 3692 8484 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9582 3720 9588 3732
rect 9539 3692 9588 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 12342 3720 12348 3732
rect 12303 3692 12348 3720
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 4246 3612 4252 3664
rect 4304 3652 4310 3664
rect 5353 3655 5411 3661
rect 5353 3652 5365 3655
rect 4304 3624 5365 3652
rect 4304 3612 4310 3624
rect 5353 3621 5365 3624
rect 5399 3621 5411 3655
rect 5353 3615 5411 3621
rect 5902 3612 5908 3664
rect 5960 3652 5966 3664
rect 6917 3655 6975 3661
rect 6917 3652 6929 3655
rect 5960 3624 6929 3652
rect 5960 3612 5966 3624
rect 6917 3621 6929 3624
rect 6963 3621 6975 3655
rect 6917 3615 6975 3621
rect 11232 3655 11290 3661
rect 11232 3621 11244 3655
rect 11278 3652 11290 3655
rect 11330 3652 11336 3664
rect 11278 3624 11336 3652
rect 11278 3621 11290 3624
rect 11232 3615 11290 3621
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3584 1823 3587
rect 2314 3584 2320 3596
rect 1811 3556 2320 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3584 2927 3587
rect 2958 3584 2964 3596
rect 2915 3556 2964 3584
rect 2915 3553 2927 3556
rect 2869 3547 2927 3553
rect 2958 3544 2964 3556
rect 3016 3584 3022 3596
rect 3418 3584 3424 3596
rect 3016 3556 3424 3584
rect 3016 3544 3022 3556
rect 3418 3544 3424 3556
rect 3476 3544 3482 3596
rect 4890 3544 4896 3596
rect 4948 3584 4954 3596
rect 7926 3584 7932 3596
rect 4948 3556 7932 3584
rect 4948 3544 4954 3556
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 8754 3584 8760 3596
rect 8527 3556 8760 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 10686 3584 10692 3596
rect 9723 3556 10692 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10870 3544 10876 3596
rect 10928 3584 10934 3596
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10928 3556 10977 3584
rect 10928 3544 10934 3556
rect 10965 3553 10977 3556
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 4212 3488 4261 3516
rect 4212 3476 4218 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 5445 3519 5503 3525
rect 5445 3516 5457 3519
rect 5408 3488 5457 3516
rect 5408 3476 5414 3488
rect 5445 3485 5457 3488
rect 5491 3516 5503 3519
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 5491 3488 7021 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 8938 3516 8944 3528
rect 8711 3488 8944 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 13446 3516 13452 3528
rect 13407 3488 13452 3516
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3448 2007 3451
rect 2590 3448 2596 3460
rect 1995 3420 2596 3448
rect 1995 3417 2007 3420
rect 1949 3411 2007 3417
rect 2590 3408 2596 3420
rect 2648 3408 2654 3460
rect 6457 3451 6515 3457
rect 6457 3417 6469 3451
rect 6503 3448 6515 3451
rect 7190 3448 7196 3460
rect 6503 3420 7196 3448
rect 6503 3417 6515 3420
rect 6457 3411 6515 3417
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13265 3451 13323 3457
rect 13265 3448 13277 3451
rect 12492 3420 13277 3448
rect 12492 3408 12498 3420
rect 13265 3417 13277 3420
rect 13311 3417 13323 3451
rect 13265 3411 13323 3417
rect 3050 3380 3056 3392
rect 3011 3352 3056 3380
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 5905 3383 5963 3389
rect 5905 3380 5917 3383
rect 5500 3352 5917 3380
rect 5500 3340 5506 3352
rect 5905 3349 5917 3352
rect 5951 3380 5963 3383
rect 7742 3380 7748 3392
rect 5951 3352 7748 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 7742 3340 7748 3352
rect 7800 3380 7806 3392
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 7800 3352 7849 3380
rect 7800 3340 7806 3352
rect 7837 3349 7849 3352
rect 7883 3349 7895 3383
rect 7837 3343 7895 3349
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8904 3352 9045 3380
rect 8904 3340 8910 3352
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9033 3343 9091 3349
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 9861 3383 9919 3389
rect 9861 3380 9873 3383
rect 9732 3352 9873 3380
rect 9732 3340 9738 3352
rect 9861 3349 9873 3352
rect 9907 3349 9919 3383
rect 9861 3343 9919 3349
rect 10321 3383 10379 3389
rect 10321 3349 10333 3383
rect 10367 3380 10379 3383
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10367 3352 10885 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 10873 3349 10885 3352
rect 10919 3380 10931 3383
rect 11330 3380 11336 3392
rect 10919 3352 11336 3380
rect 10919 3349 10931 3352
rect 10873 3343 10931 3349
rect 11330 3340 11336 3352
rect 11388 3380 11394 3392
rect 12986 3380 12992 3392
rect 11388 3352 12992 3380
rect 11388 3340 11394 3352
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 2038 3176 2044 3188
rect 1995 3148 2044 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3568 3148 3709 3176
rect 3568 3136 3574 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4246 3176 4252 3188
rect 4203 3148 4252 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5592 3148 5641 3176
rect 5592 3136 5598 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 5629 3139 5687 3145
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5960 3148 6193 3176
rect 5960 3136 5966 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6972 3148 7113 3176
rect 6972 3136 6978 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 8294 3176 8300 3188
rect 8251 3148 8300 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 8294 3136 8300 3148
rect 8352 3176 8358 3188
rect 8478 3176 8484 3188
rect 8352 3148 8484 3176
rect 8352 3136 8358 3148
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 8588 3148 10057 3176
rect 6641 3111 6699 3117
rect 6641 3077 6653 3111
rect 6687 3108 6699 3111
rect 7282 3108 7288 3120
rect 6687 3080 7288 3108
rect 6687 3077 6699 3080
rect 6641 3071 6699 3077
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 8588 3108 8616 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10686 3176 10692 3188
rect 10647 3148 10692 3176
rect 10045 3139 10103 3145
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 11057 3179 11115 3185
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 11146 3176 11152 3188
rect 11103 3148 11152 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 11146 3136 11152 3148
rect 11204 3176 11210 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11204 3148 11805 3176
rect 11204 3136 11210 3148
rect 11793 3145 11805 3148
rect 11839 3145 11851 3179
rect 11793 3139 11851 3145
rect 7760 3080 8616 3108
rect 7760 3052 7788 3080
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4212 3012 4261 3040
rect 4212 3000 4218 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 7742 3040 7748 3052
rect 7703 3012 7748 3040
rect 4249 3003 4307 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 8128 3012 8800 3040
rect 2038 2972 2044 2984
rect 1999 2944 2044 2972
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 3510 2972 3516 2984
rect 3191 2944 3516 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 7466 2972 7472 2984
rect 7427 2944 7472 2972
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 8128 2972 8156 3012
rect 7576 2944 8156 2972
rect 8665 2975 8723 2981
rect 4516 2907 4574 2913
rect 4516 2873 4528 2907
rect 4562 2904 4574 2907
rect 4706 2904 4712 2916
rect 4562 2876 4712 2904
rect 4562 2873 4574 2876
rect 4516 2867 4574 2873
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 7282 2864 7288 2916
rect 7340 2904 7346 2916
rect 7576 2913 7604 2944
rect 8665 2941 8677 2975
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 7561 2907 7619 2913
rect 7561 2904 7573 2907
rect 7340 2876 7573 2904
rect 7340 2864 7346 2876
rect 7561 2873 7573 2876
rect 7607 2873 7619 2907
rect 7561 2867 7619 2873
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 1302 2836 1308 2848
rect 256 2808 1308 2836
rect 256 2796 262 2808
rect 1302 2796 1308 2808
rect 1360 2796 1366 2848
rect 2130 2796 2136 2848
rect 2188 2836 2194 2848
rect 2225 2839 2283 2845
rect 2225 2836 2237 2839
rect 2188 2808 2237 2836
rect 2188 2796 2194 2808
rect 2225 2805 2237 2808
rect 2271 2805 2283 2839
rect 2225 2799 2283 2805
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 3510 2836 3516 2848
rect 3375 2808 3516 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 8680 2836 8708 2935
rect 8772 2904 8800 3012
rect 8938 2981 8944 2984
rect 8932 2972 8944 2981
rect 8899 2944 8944 2972
rect 8932 2935 8944 2944
rect 8938 2932 8944 2935
rect 8996 2932 9002 2984
rect 11164 2981 11192 3136
rect 11808 3040 11836 3139
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 12124 3148 12173 3176
rect 12124 3136 12130 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 12618 3176 12624 3188
rect 12483 3148 12624 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 11808 3012 12909 3040
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13262 3040 13268 3052
rect 13044 3012 13268 3040
rect 13044 3000 13050 3012
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 8846 2904 8852 2916
rect 8772 2876 8852 2904
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 9582 2836 9588 2848
rect 8619 2808 9588 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 11146 2796 11152 2848
rect 11204 2836 11210 2848
rect 11333 2839 11391 2845
rect 11333 2836 11345 2839
rect 11204 2808 11345 2836
rect 11204 2796 11210 2808
rect 11333 2805 11345 2808
rect 11379 2805 11391 2839
rect 11333 2799 11391 2805
rect 12066 2796 12072 2848
rect 12124 2836 12130 2848
rect 12802 2836 12808 2848
rect 12124 2808 12808 2836
rect 12124 2796 12130 2808
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 12894 2796 12900 2848
rect 12952 2836 12958 2848
rect 13449 2839 13507 2845
rect 13449 2836 13461 2839
rect 12952 2808 13461 2836
rect 12952 2796 12958 2808
rect 13449 2805 13461 2808
rect 13495 2805 13507 2839
rect 13449 2799 13507 2805
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 1946 2632 1952 2644
rect 1907 2604 1952 2632
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 4338 2632 4344 2644
rect 3559 2604 4344 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 2406 2496 2412 2508
rect 1811 2468 2412 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3528 2496 3556 2595
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4985 2635 5043 2641
rect 4985 2601 4997 2635
rect 5031 2632 5043 2635
rect 5258 2632 5264 2644
rect 5031 2604 5264 2632
rect 5031 2601 5043 2604
rect 4985 2595 5043 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5626 2632 5632 2644
rect 5539 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2632 5690 2644
rect 6730 2632 6736 2644
rect 5684 2604 6736 2632
rect 5684 2592 5690 2604
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 10928 2604 11713 2632
rect 10928 2592 10934 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12492 2604 12633 2632
rect 12492 2592 12498 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12621 2595 12679 2601
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 13446 2632 13452 2644
rect 13035 2604 13452 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13446 2592 13452 2604
rect 13504 2632 13510 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13504 2604 13645 2632
rect 13504 2592 13510 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 5721 2567 5779 2573
rect 5721 2533 5733 2567
rect 5767 2564 5779 2567
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 5767 2536 6377 2564
rect 5767 2533 5779 2536
rect 5721 2527 5779 2533
rect 6365 2533 6377 2536
rect 6411 2564 6423 2567
rect 7098 2564 7104 2576
rect 6411 2536 7104 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 10036 2567 10094 2573
rect 10036 2564 10048 2567
rect 9263 2536 10048 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 10036 2533 10048 2536
rect 10082 2564 10094 2567
rect 11054 2564 11060 2576
rect 10082 2536 11060 2564
rect 10082 2533 10094 2536
rect 10036 2527 10094 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 12710 2564 12716 2576
rect 12452 2536 12716 2564
rect 2915 2468 3556 2496
rect 3881 2499 3939 2505
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3927 2468 4077 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4065 2465 4077 2468
rect 4111 2496 4123 2499
rect 4246 2496 4252 2508
rect 4111 2468 4252 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7006 2496 7012 2508
rect 6963 2468 7012 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7006 2456 7012 2468
rect 7064 2496 7070 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 7064 2468 7481 2496
rect 7064 2456 7070 2468
rect 7469 2465 7481 2468
rect 7515 2465 7527 2499
rect 9582 2496 9588 2508
rect 9495 2468 9588 2496
rect 7469 2459 7527 2465
rect 9582 2456 9588 2468
rect 9640 2496 9646 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9640 2468 9781 2496
rect 9640 2456 9646 2468
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10870 2496 10876 2508
rect 9815 2468 10876 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 12452 2505 12480 2536
rect 12710 2524 12716 2536
rect 12768 2564 12774 2576
rect 13081 2567 13139 2573
rect 13081 2564 13093 2567
rect 12768 2536 13093 2564
rect 12768 2524 12774 2536
rect 13081 2533 13093 2536
rect 13127 2533 13139 2567
rect 13081 2527 13139 2533
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2465 12495 2499
rect 12437 2459 12495 2465
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 5500 2400 5825 2428
rect 5500 2388 5506 2400
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8536 2400 8585 2428
rect 8536 2388 8542 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 8938 2428 8944 2440
rect 8803 2400 8944 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 2774 2320 2780 2372
rect 2832 2360 2838 2372
rect 2832 2332 2877 2360
rect 2832 2320 2838 2332
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 3016 2332 4261 2360
rect 3016 2320 3022 2332
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 8021 2363 8079 2369
rect 8021 2329 8033 2363
rect 8067 2360 8079 2363
rect 8772 2360 8800 2391
rect 8938 2388 8944 2400
rect 8996 2428 9002 2440
rect 13262 2428 13268 2440
rect 8996 2400 9168 2428
rect 13175 2400 13268 2428
rect 8996 2388 9002 2400
rect 8067 2332 8800 2360
rect 8067 2329 8079 2332
rect 8021 2323 8079 2329
rect 2406 2292 2412 2304
rect 2367 2264 2412 2292
rect 2406 2252 2412 2264
rect 2464 2252 2470 2304
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 3326 2292 3332 2304
rect 3099 2264 3332 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 3326 2252 3332 2264
rect 3384 2252 3390 2304
rect 5258 2292 5264 2304
rect 5219 2264 5264 2292
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 9140 2292 9168 2400
rect 13262 2388 13268 2400
rect 13320 2428 13326 2440
rect 14001 2431 14059 2437
rect 14001 2428 14013 2431
rect 13320 2400 14013 2428
rect 13320 2388 13326 2400
rect 14001 2397 14013 2400
rect 14047 2397 14059 2431
rect 14001 2391 14059 2397
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 9140 2264 11161 2292
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11149 2255 11207 2261
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 14148 2264 14381 2292
rect 14148 2252 14154 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 10594 2048 10600 2100
rect 10652 2088 10658 2100
rect 12526 2088 12532 2100
rect 10652 2060 12532 2088
rect 10652 2048 10658 2060
rect 12526 2048 12532 2060
rect 12584 2048 12590 2100
rect 5810 552 5816 604
rect 5868 592 5874 604
rect 6178 592 6184 604
rect 5868 564 6184 592
rect 5868 552 5874 564
rect 6178 552 6184 564
rect 6236 552 6242 604
rect 9766 552 9772 604
rect 9824 592 9830 604
rect 9950 592 9956 604
rect 9824 564 9956 592
rect 9824 552 9830 564
rect 9950 552 9956 564
rect 10008 552 10014 604
rect 10226 552 10232 604
rect 10284 592 10290 604
rect 12158 592 12164 604
rect 10284 564 12164 592
rect 10284 552 10290 564
rect 12158 552 12164 564
rect 12216 552 12222 604
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 5356 36864 5408 36916
rect 5908 36567 5960 36576
rect 5908 36533 5917 36567
rect 5917 36533 5951 36567
rect 5951 36533 5960 36567
rect 5908 36524 5960 36533
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 6184 36320 6236 36372
rect 9864 36363 9916 36372
rect 9864 36329 9873 36363
rect 9873 36329 9907 36363
rect 9907 36329 9916 36363
rect 9864 36320 9916 36329
rect 5448 36227 5500 36236
rect 5448 36193 5457 36227
rect 5457 36193 5491 36227
rect 5491 36193 5500 36227
rect 5448 36184 5500 36193
rect 9680 36227 9732 36236
rect 9680 36193 9689 36227
rect 9689 36193 9723 36227
rect 9723 36193 9732 36227
rect 9680 36184 9732 36193
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 1584 35819 1636 35828
rect 1584 35785 1593 35819
rect 1593 35785 1627 35819
rect 1627 35785 1636 35819
rect 1584 35776 1636 35785
rect 3332 35776 3384 35828
rect 3976 35776 4028 35828
rect 6644 35776 6696 35828
rect 7380 35776 7432 35828
rect 9588 35819 9640 35828
rect 9588 35785 9597 35819
rect 9597 35785 9631 35819
rect 9631 35785 9640 35819
rect 9588 35776 9640 35785
rect 5724 35708 5776 35760
rect 9864 35751 9916 35760
rect 9864 35717 9873 35751
rect 9873 35717 9907 35751
rect 9907 35717 9916 35751
rect 9864 35708 9916 35717
rect 4436 35640 4488 35692
rect 5448 35683 5500 35692
rect 5448 35649 5457 35683
rect 5457 35649 5491 35683
rect 5491 35649 5500 35683
rect 5448 35640 5500 35649
rect 2780 35572 2832 35624
rect 1860 35479 1912 35488
rect 1860 35445 1869 35479
rect 1869 35445 1903 35479
rect 1903 35445 1912 35479
rect 1860 35436 1912 35445
rect 4620 35479 4672 35488
rect 4620 35445 4629 35479
rect 4629 35445 4663 35479
rect 4663 35445 4672 35479
rect 4620 35436 4672 35445
rect 6736 35436 6788 35488
rect 8116 35436 8168 35488
rect 8668 35436 8720 35488
rect 10416 35436 10468 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 940 35232 992 35284
rect 2136 35232 2188 35284
rect 4712 35275 4764 35284
rect 4712 35241 4721 35275
rect 4721 35241 4755 35275
rect 4755 35241 4764 35275
rect 4712 35232 4764 35241
rect 4988 35232 5040 35284
rect 7564 35275 7616 35284
rect 7564 35241 7573 35275
rect 7573 35241 7607 35275
rect 7607 35241 7616 35275
rect 7564 35232 7616 35241
rect 12532 35275 12584 35284
rect 12532 35241 12541 35275
rect 12541 35241 12575 35275
rect 12575 35241 12584 35275
rect 12532 35232 12584 35241
rect 1676 35096 1728 35148
rect 2504 35139 2556 35148
rect 2504 35105 2513 35139
rect 2513 35105 2547 35139
rect 2547 35105 2556 35139
rect 2504 35096 2556 35105
rect 4712 35096 4764 35148
rect 5632 35139 5684 35148
rect 5632 35105 5641 35139
rect 5641 35105 5675 35139
rect 5675 35105 5684 35139
rect 5632 35096 5684 35105
rect 7196 35096 7248 35148
rect 8484 35139 8536 35148
rect 8484 35105 8493 35139
rect 8493 35105 8527 35139
rect 8527 35105 8536 35139
rect 8484 35096 8536 35105
rect 9496 35096 9548 35148
rect 9680 35071 9732 35080
rect 9680 35037 9689 35071
rect 9689 35037 9723 35071
rect 9723 35037 9732 35071
rect 9680 35028 9732 35037
rect 6920 34960 6972 35012
rect 7656 34892 7708 34944
rect 11152 34892 11204 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 204 34688 256 34740
rect 12072 34688 12124 34740
rect 5632 34620 5684 34672
rect 7380 34620 7432 34672
rect 12256 34552 12308 34604
rect 2044 34527 2096 34536
rect 2044 34493 2053 34527
rect 2053 34493 2087 34527
rect 2087 34493 2096 34527
rect 2044 34484 2096 34493
rect 2136 34484 2188 34536
rect 2504 34527 2556 34536
rect 2504 34493 2513 34527
rect 2513 34493 2547 34527
rect 2547 34493 2556 34527
rect 2504 34484 2556 34493
rect 4068 34484 4120 34536
rect 7656 34527 7708 34536
rect 7656 34493 7690 34527
rect 7690 34493 7708 34527
rect 3516 34416 3568 34468
rect 7656 34484 7708 34493
rect 8208 34484 8260 34536
rect 8484 34484 8536 34536
rect 9680 34484 9732 34536
rect 7748 34416 7800 34468
rect 4804 34391 4856 34400
rect 4804 34357 4813 34391
rect 4813 34357 4847 34391
rect 4847 34357 4856 34391
rect 4804 34348 4856 34357
rect 7196 34391 7248 34400
rect 7196 34357 7205 34391
rect 7205 34357 7239 34391
rect 7239 34357 7248 34391
rect 7196 34348 7248 34357
rect 8576 34348 8628 34400
rect 9496 34348 9548 34400
rect 12072 34484 12124 34536
rect 11152 34416 11204 34468
rect 12532 34484 12584 34536
rect 9956 34348 10008 34400
rect 12072 34348 12124 34400
rect 12256 34348 12308 34400
rect 12440 34391 12492 34400
rect 12440 34357 12449 34391
rect 12449 34357 12483 34391
rect 12483 34357 12492 34391
rect 12808 34391 12860 34400
rect 12440 34348 12492 34357
rect 12808 34357 12817 34391
rect 12817 34357 12851 34391
rect 12851 34357 12860 34391
rect 12808 34348 12860 34357
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 1400 34144 1452 34196
rect 2964 34144 3016 34196
rect 4160 34144 4212 34196
rect 9496 34187 9548 34196
rect 9496 34153 9505 34187
rect 9505 34153 9539 34187
rect 9539 34153 9548 34187
rect 9496 34144 9548 34153
rect 9956 34187 10008 34196
rect 9956 34153 9965 34187
rect 9965 34153 9999 34187
rect 9999 34153 10008 34187
rect 9956 34144 10008 34153
rect 11244 34144 11296 34196
rect 1676 34119 1728 34128
rect 1676 34085 1685 34119
rect 1685 34085 1719 34119
rect 1719 34085 1728 34119
rect 1676 34076 1728 34085
rect 10876 34076 10928 34128
rect 12072 34076 12124 34128
rect 1952 34008 2004 34060
rect 3148 34008 3200 34060
rect 4160 34008 4212 34060
rect 4988 34008 5040 34060
rect 7012 34008 7064 34060
rect 10784 34051 10836 34060
rect 10784 34017 10793 34051
rect 10793 34017 10827 34051
rect 10827 34017 10836 34051
rect 10784 34008 10836 34017
rect 6276 33983 6328 33992
rect 6276 33949 6285 33983
rect 6285 33949 6319 33983
rect 6319 33949 6328 33983
rect 6276 33940 6328 33949
rect 10968 33983 11020 33992
rect 10968 33949 10977 33983
rect 10977 33949 11011 33983
rect 11011 33949 11020 33983
rect 10968 33940 11020 33949
rect 11888 33983 11940 33992
rect 11888 33949 11897 33983
rect 11897 33949 11931 33983
rect 11931 33949 11940 33983
rect 11888 33940 11940 33949
rect 4252 33915 4304 33924
rect 4252 33881 4261 33915
rect 4261 33881 4295 33915
rect 4295 33881 4304 33915
rect 4252 33872 4304 33881
rect 3516 33847 3568 33856
rect 3516 33813 3525 33847
rect 3525 33813 3559 33847
rect 3559 33813 3568 33847
rect 3516 33804 3568 33813
rect 4712 33847 4764 33856
rect 4712 33813 4721 33847
rect 4721 33813 4755 33847
rect 4755 33813 4764 33847
rect 4712 33804 4764 33813
rect 7656 33847 7708 33856
rect 7656 33813 7665 33847
rect 7665 33813 7699 33847
rect 7699 33813 7708 33847
rect 7656 33804 7708 33813
rect 11060 33804 11112 33856
rect 13084 33804 13136 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 1492 33600 1544 33652
rect 8300 33600 8352 33652
rect 8852 33600 8904 33652
rect 10784 33600 10836 33652
rect 2320 33507 2372 33516
rect 2320 33473 2329 33507
rect 2329 33473 2363 33507
rect 2363 33473 2372 33507
rect 2320 33464 2372 33473
rect 12072 33464 12124 33516
rect 12440 33464 12492 33516
rect 13084 33507 13136 33516
rect 13084 33473 13093 33507
rect 13093 33473 13127 33507
rect 13127 33473 13136 33507
rect 13084 33464 13136 33473
rect 1952 33439 2004 33448
rect 1952 33405 1961 33439
rect 1961 33405 1995 33439
rect 1995 33405 2004 33439
rect 1952 33396 2004 33405
rect 4068 33396 4120 33448
rect 4252 33439 4304 33448
rect 4252 33405 4261 33439
rect 4261 33405 4295 33439
rect 4295 33405 4304 33439
rect 4252 33396 4304 33405
rect 6276 33396 6328 33448
rect 7748 33396 7800 33448
rect 10140 33396 10192 33448
rect 11244 33396 11296 33448
rect 11888 33439 11940 33448
rect 11888 33405 11897 33439
rect 11897 33405 11931 33439
rect 11931 33405 11940 33439
rect 11888 33396 11940 33405
rect 3148 33260 3200 33312
rect 3424 33260 3476 33312
rect 4804 33328 4856 33380
rect 8208 33328 8260 33380
rect 10232 33328 10284 33380
rect 12348 33328 12400 33380
rect 4160 33303 4212 33312
rect 4160 33269 4169 33303
rect 4169 33269 4203 33303
rect 4203 33269 4212 33303
rect 4160 33260 4212 33269
rect 7012 33303 7064 33312
rect 7012 33269 7021 33303
rect 7021 33269 7055 33303
rect 7055 33269 7064 33303
rect 7012 33260 7064 33269
rect 12440 33303 12492 33312
rect 12440 33269 12449 33303
rect 12449 33269 12483 33303
rect 12483 33269 12492 33303
rect 12440 33260 12492 33269
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 1584 33099 1636 33108
rect 1584 33065 1593 33099
rect 1593 33065 1627 33099
rect 1627 33065 1636 33099
rect 1584 33056 1636 33065
rect 4252 33099 4304 33108
rect 4252 33065 4261 33099
rect 4261 33065 4295 33099
rect 4295 33065 4304 33099
rect 4252 33056 4304 33065
rect 6644 33056 6696 33108
rect 7564 33099 7616 33108
rect 7564 33065 7573 33099
rect 7573 33065 7607 33099
rect 7607 33065 7616 33099
rect 7564 33056 7616 33065
rect 10784 33099 10836 33108
rect 10784 33065 10793 33099
rect 10793 33065 10827 33099
rect 10827 33065 10836 33099
rect 10784 33056 10836 33065
rect 11060 33056 11112 33108
rect 12348 33099 12400 33108
rect 12348 33065 12357 33099
rect 12357 33065 12391 33099
rect 12391 33065 12400 33099
rect 12348 33056 12400 33065
rect 12900 33056 12952 33108
rect 15752 33056 15804 33108
rect 7288 32988 7340 33040
rect 7472 33031 7524 33040
rect 7472 32997 7481 33031
rect 7481 32997 7515 33031
rect 7515 32997 7524 33031
rect 7472 32988 7524 32997
rect 12072 32988 12124 33040
rect 1676 32920 1728 32972
rect 10048 32920 10100 32972
rect 12348 32920 12400 32972
rect 12716 32963 12768 32972
rect 12716 32929 12725 32963
rect 12725 32929 12759 32963
rect 12759 32929 12768 32963
rect 12716 32920 12768 32929
rect 6000 32895 6052 32904
rect 6000 32861 6009 32895
rect 6009 32861 6043 32895
rect 6043 32861 6052 32895
rect 6000 32852 6052 32861
rect 6184 32895 6236 32904
rect 6184 32861 6193 32895
rect 6193 32861 6227 32895
rect 6227 32861 6236 32895
rect 6184 32852 6236 32861
rect 6552 32852 6604 32904
rect 7012 32852 7064 32904
rect 9588 32852 9640 32904
rect 11428 32895 11480 32904
rect 11428 32861 11437 32895
rect 11437 32861 11471 32895
rect 11471 32861 11480 32895
rect 11428 32852 11480 32861
rect 9496 32784 9548 32836
rect 10784 32784 10836 32836
rect 11152 32784 11204 32836
rect 4988 32716 5040 32768
rect 5540 32759 5592 32768
rect 5540 32725 5549 32759
rect 5549 32725 5583 32759
rect 5583 32725 5592 32759
rect 5540 32716 5592 32725
rect 7012 32759 7064 32768
rect 7012 32725 7021 32759
rect 7021 32725 7055 32759
rect 7055 32725 7064 32759
rect 7012 32716 7064 32725
rect 8300 32716 8352 32768
rect 9404 32759 9456 32768
rect 9404 32725 9413 32759
rect 9413 32725 9447 32759
rect 9447 32725 9456 32759
rect 9404 32716 9456 32725
rect 10968 32716 11020 32768
rect 11520 32716 11572 32768
rect 12072 32716 12124 32768
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 7104 32512 7156 32564
rect 7564 32512 7616 32564
rect 8576 32555 8628 32564
rect 8576 32521 8585 32555
rect 8585 32521 8619 32555
rect 8619 32521 8628 32555
rect 8576 32512 8628 32521
rect 8852 32555 8904 32564
rect 8852 32521 8861 32555
rect 8861 32521 8895 32555
rect 8895 32521 8904 32555
rect 8852 32512 8904 32521
rect 1676 32487 1728 32496
rect 1676 32453 1685 32487
rect 1685 32453 1719 32487
rect 1719 32453 1728 32487
rect 1676 32444 1728 32453
rect 6000 32444 6052 32496
rect 7472 32487 7524 32496
rect 7472 32453 7481 32487
rect 7481 32453 7515 32487
rect 7515 32453 7524 32487
rect 7472 32444 7524 32453
rect 5816 32308 5868 32360
rect 9496 32419 9548 32428
rect 9496 32385 9505 32419
rect 9505 32385 9539 32419
rect 9539 32385 9548 32419
rect 9496 32376 9548 32385
rect 9680 32512 9732 32564
rect 10140 32512 10192 32564
rect 10876 32512 10928 32564
rect 12900 32555 12952 32564
rect 12900 32521 12909 32555
rect 12909 32521 12943 32555
rect 12943 32521 12952 32555
rect 12900 32512 12952 32521
rect 12072 32376 12124 32428
rect 12716 32376 12768 32428
rect 7012 32308 7064 32360
rect 9404 32351 9456 32360
rect 9404 32317 9413 32351
rect 9413 32317 9447 32351
rect 9447 32317 9456 32351
rect 9404 32308 9456 32317
rect 9680 32308 9732 32360
rect 4160 32240 4212 32292
rect 6092 32240 6144 32292
rect 6552 32283 6604 32292
rect 6552 32249 6561 32283
rect 6561 32249 6595 32283
rect 6595 32249 6604 32283
rect 6552 32240 6604 32249
rect 6828 32240 6880 32292
rect 5632 32215 5684 32224
rect 5632 32181 5641 32215
rect 5641 32181 5675 32215
rect 5675 32181 5684 32215
rect 6184 32215 6236 32224
rect 5632 32172 5684 32181
rect 6184 32181 6193 32215
rect 6193 32181 6227 32215
rect 6227 32181 6236 32215
rect 6184 32172 6236 32181
rect 10416 32172 10468 32224
rect 11152 32215 11204 32224
rect 11152 32181 11161 32215
rect 11161 32181 11195 32215
rect 11195 32181 11204 32215
rect 11152 32172 11204 32181
rect 12072 32172 12124 32224
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 6000 32011 6052 32020
rect 6000 31977 6009 32011
rect 6009 31977 6043 32011
rect 6043 31977 6052 32011
rect 6000 31968 6052 31977
rect 6644 31968 6696 32020
rect 6828 32011 6880 32020
rect 6828 31977 6837 32011
rect 6837 31977 6871 32011
rect 6871 31977 6880 32011
rect 6828 31968 6880 31977
rect 7012 31968 7064 32020
rect 10048 32011 10100 32020
rect 10048 31977 10057 32011
rect 10057 31977 10091 32011
rect 10091 31977 10100 32011
rect 10048 31968 10100 31977
rect 10232 31968 10284 32020
rect 10508 32011 10560 32020
rect 10508 31977 10517 32011
rect 10517 31977 10551 32011
rect 10551 31977 10560 32011
rect 10508 31968 10560 31977
rect 11060 31968 11112 32020
rect 12072 31968 12124 32020
rect 4252 31900 4304 31952
rect 7288 31900 7340 31952
rect 4068 31875 4120 31884
rect 4068 31841 4077 31875
rect 4077 31841 4111 31875
rect 4111 31841 4120 31875
rect 4068 31832 4120 31841
rect 5080 31832 5132 31884
rect 6184 31832 6236 31884
rect 7748 31875 7800 31884
rect 7748 31841 7757 31875
rect 7757 31841 7791 31875
rect 7791 31841 7800 31875
rect 7748 31832 7800 31841
rect 11428 31832 11480 31884
rect 12348 31832 12400 31884
rect 7564 31764 7616 31816
rect 8024 31807 8076 31816
rect 8024 31773 8033 31807
rect 8033 31773 8067 31807
rect 8067 31773 8076 31807
rect 8024 31764 8076 31773
rect 8852 31764 8904 31816
rect 10416 31764 10468 31816
rect 10784 31807 10836 31816
rect 10784 31773 10793 31807
rect 10793 31773 10827 31807
rect 10827 31773 10836 31807
rect 10784 31764 10836 31773
rect 11152 31764 11204 31816
rect 12072 31764 12124 31816
rect 7656 31696 7708 31748
rect 3056 31671 3108 31680
rect 3056 31637 3065 31671
rect 3065 31637 3099 31671
rect 3099 31637 3108 31671
rect 3056 31628 3108 31637
rect 5448 31671 5500 31680
rect 5448 31637 5457 31671
rect 5457 31637 5491 31671
rect 5491 31637 5500 31671
rect 5448 31628 5500 31637
rect 8300 31628 8352 31680
rect 9312 31628 9364 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 4068 31467 4120 31476
rect 4068 31433 4077 31467
rect 4077 31433 4111 31467
rect 4111 31433 4120 31467
rect 4068 31424 4120 31433
rect 4620 31424 4672 31476
rect 4896 31424 4948 31476
rect 4988 31424 5040 31476
rect 5356 31424 5408 31476
rect 7748 31424 7800 31476
rect 9404 31424 9456 31476
rect 10784 31424 10836 31476
rect 13728 31467 13780 31476
rect 13728 31433 13737 31467
rect 13737 31433 13771 31467
rect 13771 31433 13780 31467
rect 13728 31424 13780 31433
rect 8024 31356 8076 31408
rect 3516 31288 3568 31340
rect 4620 31288 4672 31340
rect 5080 31331 5132 31340
rect 5080 31297 5089 31331
rect 5089 31297 5123 31331
rect 5123 31297 5132 31331
rect 5080 31288 5132 31297
rect 8576 31288 8628 31340
rect 8760 31288 8812 31340
rect 9312 31288 9364 31340
rect 10232 31288 10284 31340
rect 12624 31288 12676 31340
rect 12900 31288 12952 31340
rect 4988 31263 5040 31272
rect 4988 31229 4997 31263
rect 4997 31229 5031 31263
rect 5031 31229 5040 31263
rect 4988 31220 5040 31229
rect 9588 31220 9640 31272
rect 13544 31263 13596 31272
rect 13544 31229 13553 31263
rect 13553 31229 13587 31263
rect 13587 31229 13596 31263
rect 13544 31220 13596 31229
rect 2412 31152 2464 31204
rect 4160 31152 4212 31204
rect 2964 31127 3016 31136
rect 2964 31093 2973 31127
rect 2973 31093 3007 31127
rect 3007 31093 3016 31127
rect 2964 31084 3016 31093
rect 3056 31084 3108 31136
rect 4436 31084 4488 31136
rect 7564 31084 7616 31136
rect 9312 31084 9364 31136
rect 9956 31084 10008 31136
rect 10416 31084 10468 31136
rect 10508 31084 10560 31136
rect 10968 31084 11020 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 2412 30923 2464 30932
rect 2412 30889 2421 30923
rect 2421 30889 2455 30923
rect 2455 30889 2464 30923
rect 2412 30880 2464 30889
rect 2780 30923 2832 30932
rect 2780 30889 2789 30923
rect 2789 30889 2823 30923
rect 2823 30889 2832 30923
rect 5540 30923 5592 30932
rect 2780 30880 2832 30889
rect 5540 30889 5549 30923
rect 5549 30889 5583 30923
rect 5583 30889 5592 30923
rect 5540 30880 5592 30889
rect 6828 30880 6880 30932
rect 7656 30880 7708 30932
rect 7748 30880 7800 30932
rect 8116 30880 8168 30932
rect 9680 30923 9732 30932
rect 9680 30889 9689 30923
rect 9689 30889 9723 30923
rect 9723 30889 9732 30923
rect 9680 30880 9732 30889
rect 12440 30880 12492 30932
rect 2228 30812 2280 30864
rect 8576 30812 8628 30864
rect 9588 30812 9640 30864
rect 11520 30812 11572 30864
rect 4344 30744 4396 30796
rect 10048 30787 10100 30796
rect 10048 30753 10057 30787
rect 10057 30753 10091 30787
rect 10091 30753 10100 30787
rect 10048 30744 10100 30753
rect 10692 30744 10744 30796
rect 2872 30676 2924 30728
rect 4528 30719 4580 30728
rect 3240 30608 3292 30660
rect 4528 30685 4537 30719
rect 4537 30685 4571 30719
rect 4571 30685 4580 30719
rect 4528 30676 4580 30685
rect 4620 30676 4672 30728
rect 5448 30676 5500 30728
rect 6184 30676 6236 30728
rect 8392 30719 8444 30728
rect 4988 30608 5040 30660
rect 6092 30608 6144 30660
rect 6644 30608 6696 30660
rect 8392 30685 8401 30719
rect 8401 30685 8435 30719
rect 8435 30685 8444 30719
rect 8392 30676 8444 30685
rect 8300 30608 8352 30660
rect 10232 30719 10284 30728
rect 10232 30685 10241 30719
rect 10241 30685 10275 30719
rect 10275 30685 10284 30719
rect 10232 30676 10284 30685
rect 11244 30676 11296 30728
rect 11428 30676 11480 30728
rect 5816 30583 5868 30592
rect 5816 30549 5825 30583
rect 5825 30549 5859 30583
rect 5859 30549 5868 30583
rect 5816 30540 5868 30549
rect 6920 30540 6972 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 2228 30336 2280 30388
rect 4620 30336 4672 30388
rect 6184 30379 6236 30388
rect 6184 30345 6193 30379
rect 6193 30345 6227 30379
rect 6227 30345 6236 30379
rect 6184 30336 6236 30345
rect 10232 30336 10284 30388
rect 11520 30336 11572 30388
rect 7840 30268 7892 30320
rect 8116 30268 8168 30320
rect 9772 30268 9824 30320
rect 10048 30268 10100 30320
rect 2964 30200 3016 30252
rect 3424 30243 3476 30252
rect 3424 30209 3433 30243
rect 3433 30209 3467 30243
rect 3467 30209 3476 30243
rect 3424 30200 3476 30209
rect 5540 30200 5592 30252
rect 6000 30200 6052 30252
rect 6920 30200 6972 30252
rect 7288 30243 7340 30252
rect 7288 30209 7297 30243
rect 7297 30209 7331 30243
rect 7331 30209 7340 30243
rect 7288 30200 7340 30209
rect 7656 30200 7708 30252
rect 10508 30200 10560 30252
rect 3240 30175 3292 30184
rect 3240 30141 3249 30175
rect 3249 30141 3283 30175
rect 3283 30141 3292 30175
rect 3240 30132 3292 30141
rect 5908 30132 5960 30184
rect 5816 30064 5868 30116
rect 2504 30039 2556 30048
rect 2504 30005 2513 30039
rect 2513 30005 2547 30039
rect 2547 30005 2556 30039
rect 2504 29996 2556 30005
rect 2872 30039 2924 30048
rect 2872 30005 2881 30039
rect 2881 30005 2915 30039
rect 2915 30005 2924 30039
rect 2872 29996 2924 30005
rect 4528 30039 4580 30048
rect 4528 30005 4537 30039
rect 4537 30005 4571 30039
rect 4571 30005 4580 30039
rect 4528 29996 4580 30005
rect 4988 30039 5040 30048
rect 4988 30005 4997 30039
rect 4997 30005 5031 30039
rect 5031 30005 5040 30039
rect 4988 29996 5040 30005
rect 5172 30039 5224 30048
rect 5172 30005 5181 30039
rect 5181 30005 5215 30039
rect 5215 30005 5224 30039
rect 5172 29996 5224 30005
rect 7932 30132 7984 30184
rect 9772 30132 9824 30184
rect 9680 30064 9732 30116
rect 10232 30064 10284 30116
rect 11428 30064 11480 30116
rect 7196 30039 7248 30048
rect 7196 30005 7205 30039
rect 7205 30005 7239 30039
rect 7239 30005 7248 30039
rect 7196 29996 7248 30005
rect 8300 30039 8352 30048
rect 8300 30005 8309 30039
rect 8309 30005 8343 30039
rect 8343 30005 8352 30039
rect 8300 29996 8352 30005
rect 8760 29996 8812 30048
rect 9588 30039 9640 30048
rect 9588 30005 9597 30039
rect 9597 30005 9631 30039
rect 9631 30005 9640 30039
rect 9588 29996 9640 30005
rect 9772 29996 9824 30048
rect 10692 30039 10744 30048
rect 10692 30005 10701 30039
rect 10701 30005 10735 30039
rect 10735 30005 10744 30039
rect 10692 29996 10744 30005
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 2964 29792 3016 29844
rect 4344 29835 4396 29844
rect 4344 29801 4353 29835
rect 4353 29801 4387 29835
rect 4387 29801 4396 29835
rect 4344 29792 4396 29801
rect 6920 29835 6972 29844
rect 6920 29801 6929 29835
rect 6929 29801 6963 29835
rect 6963 29801 6972 29835
rect 6920 29792 6972 29801
rect 7288 29792 7340 29844
rect 6644 29724 6696 29776
rect 2320 29656 2372 29708
rect 3424 29656 3476 29708
rect 4988 29656 5040 29708
rect 6000 29656 6052 29708
rect 8024 29656 8076 29708
rect 8668 29656 8720 29708
rect 10508 29699 10560 29708
rect 10508 29665 10542 29699
rect 10542 29665 10560 29699
rect 10508 29656 10560 29665
rect 4804 29588 4856 29640
rect 7748 29588 7800 29640
rect 8576 29588 8628 29640
rect 10232 29631 10284 29640
rect 10232 29597 10241 29631
rect 10241 29597 10275 29631
rect 10275 29597 10284 29631
rect 10232 29588 10284 29597
rect 2780 29452 2832 29504
rect 6276 29495 6328 29504
rect 6276 29461 6285 29495
rect 6285 29461 6319 29495
rect 6319 29461 6328 29495
rect 6276 29452 6328 29461
rect 7932 29452 7984 29504
rect 8392 29452 8444 29504
rect 9404 29452 9456 29504
rect 9772 29452 9824 29504
rect 11612 29495 11664 29504
rect 11612 29461 11621 29495
rect 11621 29461 11655 29495
rect 11655 29461 11664 29495
rect 11612 29452 11664 29461
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 1584 29291 1636 29300
rect 1584 29257 1593 29291
rect 1593 29257 1627 29291
rect 1627 29257 1636 29291
rect 1584 29248 1636 29257
rect 2872 29248 2924 29300
rect 4804 29248 4856 29300
rect 5448 29248 5500 29300
rect 8024 29248 8076 29300
rect 8300 29248 8352 29300
rect 2320 29223 2372 29232
rect 2320 29189 2329 29223
rect 2329 29189 2363 29223
rect 2363 29189 2372 29223
rect 2320 29180 2372 29189
rect 4068 29155 4120 29164
rect 4068 29121 4077 29155
rect 4077 29121 4111 29155
rect 4111 29121 4120 29155
rect 4068 29112 4120 29121
rect 5172 29112 5224 29164
rect 7196 29180 7248 29232
rect 8208 29180 8260 29232
rect 9496 29180 9548 29232
rect 6276 29112 6328 29164
rect 11244 29155 11296 29164
rect 11244 29121 11253 29155
rect 11253 29121 11287 29155
rect 11287 29121 11296 29155
rect 11244 29112 11296 29121
rect 7012 29044 7064 29096
rect 7472 29044 7524 29096
rect 8392 29044 8444 29096
rect 7748 29019 7800 29028
rect 7748 28985 7757 29019
rect 7757 28985 7791 29019
rect 7791 28985 7800 29019
rect 7748 28976 7800 28985
rect 8576 29019 8628 29028
rect 8576 28985 8610 29019
rect 8610 28985 8628 29019
rect 8576 28976 8628 28985
rect 5908 28908 5960 28960
rect 7472 28951 7524 28960
rect 7472 28917 7481 28951
rect 7481 28917 7515 28951
rect 7515 28917 7524 28951
rect 7472 28908 7524 28917
rect 10048 28976 10100 29028
rect 10232 29019 10284 29028
rect 10232 28985 10241 29019
rect 10241 28985 10275 29019
rect 10275 28985 10284 29019
rect 10232 28976 10284 28985
rect 10416 28976 10468 29028
rect 11612 29112 11664 29164
rect 10784 28908 10836 28960
rect 10876 28908 10928 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 2780 28704 2832 28756
rect 4528 28747 4580 28756
rect 4528 28713 4537 28747
rect 4537 28713 4571 28747
rect 4571 28713 4580 28747
rect 4528 28704 4580 28713
rect 7472 28704 7524 28756
rect 8576 28704 8628 28756
rect 10876 28747 10928 28756
rect 10876 28713 10885 28747
rect 10885 28713 10919 28747
rect 10919 28713 10928 28747
rect 10876 28704 10928 28713
rect 3516 28636 3568 28688
rect 4804 28568 4856 28620
rect 4988 28543 5040 28552
rect 4988 28509 4997 28543
rect 4997 28509 5031 28543
rect 5031 28509 5040 28543
rect 4988 28500 5040 28509
rect 6184 28636 6236 28688
rect 11428 28636 11480 28688
rect 12348 28636 12400 28688
rect 5448 28568 5500 28620
rect 6368 28568 6420 28620
rect 8392 28611 8444 28620
rect 8392 28577 8401 28611
rect 8401 28577 8435 28611
rect 8435 28577 8444 28611
rect 8392 28568 8444 28577
rect 10232 28568 10284 28620
rect 11060 28568 11112 28620
rect 5264 28500 5316 28552
rect 6000 28432 6052 28484
rect 10508 28432 10560 28484
rect 5908 28407 5960 28416
rect 5908 28373 5917 28407
rect 5917 28373 5951 28407
rect 5951 28373 5960 28407
rect 5908 28364 5960 28373
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 2872 28203 2924 28212
rect 2872 28169 2881 28203
rect 2881 28169 2915 28203
rect 2915 28169 2924 28203
rect 2872 28160 2924 28169
rect 3056 28203 3108 28212
rect 3056 28169 3065 28203
rect 3065 28169 3099 28203
rect 3099 28169 3108 28203
rect 3056 28160 3108 28169
rect 4988 28203 5040 28212
rect 4988 28169 4997 28203
rect 4997 28169 5031 28203
rect 5031 28169 5040 28203
rect 4988 28160 5040 28169
rect 5264 28203 5316 28212
rect 5264 28169 5273 28203
rect 5273 28169 5307 28203
rect 5307 28169 5316 28203
rect 5264 28160 5316 28169
rect 6184 28160 6236 28212
rect 6368 28203 6420 28212
rect 6368 28169 6377 28203
rect 6377 28169 6411 28203
rect 6411 28169 6420 28203
rect 6368 28160 6420 28169
rect 8392 28160 8444 28212
rect 8852 28160 8904 28212
rect 9404 28203 9456 28212
rect 9404 28169 9413 28203
rect 9413 28169 9447 28203
rect 9447 28169 9456 28203
rect 9404 28160 9456 28169
rect 11060 28203 11112 28212
rect 11060 28169 11069 28203
rect 11069 28169 11103 28203
rect 11103 28169 11112 28203
rect 11060 28160 11112 28169
rect 11428 28203 11480 28212
rect 11428 28169 11437 28203
rect 11437 28169 11471 28203
rect 11471 28169 11480 28203
rect 11428 28160 11480 28169
rect 3516 28024 3568 28076
rect 8576 28024 8628 28076
rect 2872 27956 2924 28008
rect 7472 27956 7524 28008
rect 2412 27888 2464 27940
rect 4804 27888 4856 27940
rect 5816 27888 5868 27940
rect 7748 27931 7800 27940
rect 7748 27897 7757 27931
rect 7757 27897 7791 27931
rect 7791 27897 7800 27931
rect 7748 27888 7800 27897
rect 8024 27820 8076 27872
rect 9588 27888 9640 27940
rect 11336 27888 11388 27940
rect 8576 27820 8628 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 2412 27659 2464 27668
rect 2412 27625 2421 27659
rect 2421 27625 2455 27659
rect 2455 27625 2464 27659
rect 2412 27616 2464 27625
rect 5264 27616 5316 27668
rect 7564 27659 7616 27668
rect 7564 27625 7573 27659
rect 7573 27625 7607 27659
rect 7607 27625 7616 27659
rect 7564 27616 7616 27625
rect 8024 27659 8076 27668
rect 8024 27625 8033 27659
rect 8033 27625 8067 27659
rect 8067 27625 8076 27659
rect 8024 27616 8076 27625
rect 10876 27659 10928 27668
rect 10876 27625 10885 27659
rect 10885 27625 10919 27659
rect 10919 27625 10928 27659
rect 10876 27616 10928 27625
rect 2044 27548 2096 27600
rect 2504 27548 2556 27600
rect 2964 27548 3016 27600
rect 7932 27591 7984 27600
rect 7932 27557 7941 27591
rect 7941 27557 7975 27591
rect 7975 27557 7984 27591
rect 7932 27548 7984 27557
rect 9588 27548 9640 27600
rect 12348 27548 12400 27600
rect 2228 27480 2280 27532
rect 2780 27523 2832 27532
rect 2780 27489 2789 27523
rect 2789 27489 2823 27523
rect 2823 27489 2832 27523
rect 4344 27523 4396 27532
rect 2780 27480 2832 27489
rect 4344 27489 4378 27523
rect 4378 27489 4396 27523
rect 4344 27480 4396 27489
rect 10048 27523 10100 27532
rect 10048 27489 10057 27523
rect 10057 27489 10091 27523
rect 10091 27489 10100 27523
rect 10048 27480 10100 27489
rect 11060 27480 11112 27532
rect 11888 27523 11940 27532
rect 11888 27489 11897 27523
rect 11897 27489 11931 27523
rect 11931 27489 11940 27523
rect 11888 27480 11940 27489
rect 4068 27455 4120 27464
rect 4068 27421 4077 27455
rect 4077 27421 4111 27455
rect 4111 27421 4120 27455
rect 4068 27412 4120 27421
rect 8116 27455 8168 27464
rect 8116 27421 8125 27455
rect 8125 27421 8159 27455
rect 8159 27421 8168 27455
rect 8116 27412 8168 27421
rect 8668 27412 8720 27464
rect 8852 27412 8904 27464
rect 10876 27412 10928 27464
rect 9588 27344 9640 27396
rect 7288 27276 7340 27328
rect 13452 27276 13504 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 4344 27072 4396 27124
rect 8024 27072 8076 27124
rect 10140 27072 10192 27124
rect 2228 27004 2280 27056
rect 2504 27047 2556 27056
rect 2504 27013 2513 27047
rect 2513 27013 2547 27047
rect 2547 27013 2556 27047
rect 2504 27004 2556 27013
rect 4068 27004 4120 27056
rect 5448 27004 5500 27056
rect 6184 27004 6236 27056
rect 2688 26868 2740 26920
rect 7288 26979 7340 26988
rect 7288 26945 7297 26979
rect 7297 26945 7331 26979
rect 7331 26945 7340 26979
rect 7288 26936 7340 26945
rect 8116 27004 8168 27056
rect 11888 27004 11940 27056
rect 7656 26936 7708 26988
rect 9496 26936 9548 26988
rect 9864 26979 9916 26988
rect 9864 26945 9873 26979
rect 9873 26945 9907 26979
rect 9907 26945 9916 26979
rect 9864 26936 9916 26945
rect 10876 26936 10928 26988
rect 11244 26936 11296 26988
rect 12992 26979 13044 26988
rect 12992 26945 13001 26979
rect 13001 26945 13035 26979
rect 13035 26945 13044 26979
rect 12992 26936 13044 26945
rect 9588 26911 9640 26920
rect 9588 26877 9597 26911
rect 9597 26877 9631 26911
rect 9631 26877 9640 26911
rect 9588 26868 9640 26877
rect 10784 26868 10836 26920
rect 2964 26800 3016 26852
rect 6828 26775 6880 26784
rect 6828 26741 6837 26775
rect 6837 26741 6871 26775
rect 6871 26741 6880 26775
rect 6828 26732 6880 26741
rect 7380 26732 7432 26784
rect 8484 26732 8536 26784
rect 8852 26732 8904 26784
rect 9312 26732 9364 26784
rect 10416 26732 10468 26784
rect 11336 26800 11388 26852
rect 12256 26843 12308 26852
rect 12256 26809 12265 26843
rect 12265 26809 12299 26843
rect 12299 26809 12308 26843
rect 12256 26800 12308 26809
rect 12808 26843 12860 26852
rect 12808 26809 12817 26843
rect 12817 26809 12851 26843
rect 12851 26809 12860 26843
rect 12808 26800 12860 26809
rect 10784 26775 10836 26784
rect 10784 26741 10793 26775
rect 10793 26741 10827 26775
rect 10827 26741 10836 26775
rect 10784 26732 10836 26741
rect 10876 26732 10928 26784
rect 11520 26732 11572 26784
rect 12440 26775 12492 26784
rect 12440 26741 12449 26775
rect 12449 26741 12483 26775
rect 12483 26741 12492 26775
rect 12440 26732 12492 26741
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 2228 26528 2280 26580
rect 2688 26571 2740 26580
rect 2688 26537 2697 26571
rect 2697 26537 2731 26571
rect 2731 26537 2740 26571
rect 2688 26528 2740 26537
rect 2964 26571 3016 26580
rect 2964 26537 2973 26571
rect 2973 26537 3007 26571
rect 3007 26537 3016 26571
rect 2964 26528 3016 26537
rect 6828 26528 6880 26580
rect 7932 26571 7984 26580
rect 7932 26537 7941 26571
rect 7941 26537 7975 26571
rect 7975 26537 7984 26571
rect 7932 26528 7984 26537
rect 10876 26571 10928 26580
rect 10876 26537 10885 26571
rect 10885 26537 10919 26571
rect 10919 26537 10928 26571
rect 10876 26528 10928 26537
rect 12348 26571 12400 26580
rect 12348 26537 12357 26571
rect 12357 26537 12391 26571
rect 12391 26537 12400 26571
rect 12348 26528 12400 26537
rect 11244 26503 11296 26512
rect 11244 26469 11278 26503
rect 11278 26469 11296 26503
rect 12992 26503 13044 26512
rect 11244 26460 11296 26469
rect 12992 26469 13001 26503
rect 13001 26469 13035 26503
rect 13035 26469 13044 26503
rect 12992 26460 13044 26469
rect 6828 26392 6880 26444
rect 10876 26392 10928 26444
rect 12348 26392 12400 26444
rect 6000 26324 6052 26376
rect 7196 26324 7248 26376
rect 5908 26299 5960 26308
rect 5908 26265 5917 26299
rect 5917 26265 5951 26299
rect 5951 26265 5960 26299
rect 5908 26256 5960 26265
rect 4988 26188 5040 26240
rect 6736 26188 6788 26240
rect 8668 26231 8720 26240
rect 8668 26197 8677 26231
rect 8677 26197 8711 26231
rect 8711 26197 8720 26231
rect 8668 26188 8720 26197
rect 9864 26188 9916 26240
rect 11152 26188 11204 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 1584 26027 1636 26036
rect 1584 25993 1593 26027
rect 1593 25993 1627 26027
rect 1627 25993 1636 26027
rect 1584 25984 1636 25993
rect 6184 26027 6236 26036
rect 6184 25993 6193 26027
rect 6193 25993 6227 26027
rect 6227 25993 6236 26027
rect 6184 25984 6236 25993
rect 6828 26027 6880 26036
rect 6828 25993 6837 26027
rect 6837 25993 6871 26027
rect 6871 25993 6880 26027
rect 6828 25984 6880 25993
rect 9864 25984 9916 26036
rect 4344 25780 4396 25832
rect 8576 25959 8628 25968
rect 8576 25925 8585 25959
rect 8585 25925 8619 25959
rect 8619 25925 8628 25959
rect 8576 25916 8628 25925
rect 9404 25848 9456 25900
rect 7196 25823 7248 25832
rect 7196 25789 7205 25823
rect 7205 25789 7239 25823
rect 7239 25789 7248 25823
rect 7196 25780 7248 25789
rect 8668 25780 8720 25832
rect 10600 25891 10652 25900
rect 10600 25857 10609 25891
rect 10609 25857 10643 25891
rect 10643 25857 10652 25891
rect 10600 25848 10652 25857
rect 11060 25984 11112 26036
rect 11244 25984 11296 26036
rect 10876 25848 10928 25900
rect 9312 25712 9364 25764
rect 10784 25780 10836 25832
rect 1952 25687 2004 25696
rect 1952 25653 1961 25687
rect 1961 25653 1995 25687
rect 1995 25653 2004 25687
rect 1952 25644 2004 25653
rect 4068 25687 4120 25696
rect 4068 25653 4077 25687
rect 4077 25653 4111 25687
rect 4111 25653 4120 25687
rect 4068 25644 4120 25653
rect 4344 25687 4396 25696
rect 4344 25653 4353 25687
rect 4353 25653 4387 25687
rect 4387 25653 4396 25687
rect 4344 25644 4396 25653
rect 4528 25687 4580 25696
rect 4528 25653 4537 25687
rect 4537 25653 4571 25687
rect 4571 25653 4580 25687
rect 4528 25644 4580 25653
rect 4988 25687 5040 25696
rect 4988 25653 4997 25687
rect 4997 25653 5031 25687
rect 5031 25653 5040 25687
rect 4988 25644 5040 25653
rect 5908 25687 5960 25696
rect 5908 25653 5917 25687
rect 5917 25653 5951 25687
rect 5951 25653 5960 25687
rect 5908 25644 5960 25653
rect 7288 25687 7340 25696
rect 7288 25653 7297 25687
rect 7297 25653 7331 25687
rect 7331 25653 7340 25687
rect 7288 25644 7340 25653
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 1952 25440 2004 25492
rect 4252 25440 4304 25492
rect 4988 25440 5040 25492
rect 5908 25440 5960 25492
rect 9312 25440 9364 25492
rect 10600 25440 10652 25492
rect 2780 25372 2832 25424
rect 6184 25372 6236 25424
rect 2688 25236 2740 25288
rect 2964 25279 3016 25288
rect 2964 25245 2973 25279
rect 2973 25245 3007 25279
rect 3007 25245 3016 25279
rect 2964 25236 3016 25245
rect 4988 25236 5040 25288
rect 2596 25168 2648 25220
rect 2412 25100 2464 25152
rect 5448 25100 5500 25152
rect 7932 25143 7984 25152
rect 7932 25109 7941 25143
rect 7941 25109 7975 25143
rect 7975 25109 7984 25143
rect 7932 25100 7984 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 4068 24939 4120 24948
rect 4068 24905 4077 24939
rect 4077 24905 4111 24939
rect 4111 24905 4120 24939
rect 4068 24896 4120 24905
rect 6184 24896 6236 24948
rect 4620 24828 4672 24880
rect 5080 24803 5132 24812
rect 5080 24769 5089 24803
rect 5089 24769 5123 24803
rect 5123 24769 5132 24803
rect 5080 24760 5132 24769
rect 2228 24692 2280 24744
rect 2412 24735 2464 24744
rect 2412 24701 2446 24735
rect 2446 24701 2464 24735
rect 2412 24692 2464 24701
rect 4988 24735 5040 24744
rect 4988 24701 4997 24735
rect 4997 24701 5031 24735
rect 5031 24701 5040 24735
rect 4988 24692 5040 24701
rect 5448 24692 5500 24744
rect 2688 24624 2740 24676
rect 7932 24692 7984 24744
rect 8668 24624 8720 24676
rect 10232 24624 10284 24676
rect 10876 24624 10928 24676
rect 2596 24556 2648 24608
rect 4804 24556 4856 24608
rect 8024 24556 8076 24608
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 2596 24352 2648 24404
rect 2780 24395 2832 24404
rect 2780 24361 2789 24395
rect 2789 24361 2823 24395
rect 2823 24361 2832 24395
rect 2780 24352 2832 24361
rect 4528 24395 4580 24404
rect 4528 24361 4537 24395
rect 4537 24361 4571 24395
rect 4571 24361 4580 24395
rect 4528 24352 4580 24361
rect 5540 24284 5592 24336
rect 7748 24327 7800 24336
rect 7748 24293 7757 24327
rect 7757 24293 7791 24327
rect 7791 24293 7800 24327
rect 7748 24284 7800 24293
rect 9312 24284 9364 24336
rect 10232 24352 10284 24404
rect 4804 24216 4856 24268
rect 10140 24216 10192 24268
rect 11060 24216 11112 24268
rect 11336 24259 11388 24268
rect 11336 24225 11345 24259
rect 11345 24225 11379 24259
rect 11379 24225 11388 24259
rect 11336 24216 11388 24225
rect 12348 24216 12400 24268
rect 4160 24148 4212 24200
rect 8024 24191 8076 24200
rect 8024 24157 8033 24191
rect 8033 24157 8067 24191
rect 8067 24157 8076 24191
rect 8024 24148 8076 24157
rect 10232 24191 10284 24200
rect 10232 24157 10241 24191
rect 10241 24157 10275 24191
rect 10275 24157 10284 24191
rect 10232 24148 10284 24157
rect 6920 24055 6972 24064
rect 6920 24021 6929 24055
rect 6929 24021 6963 24055
rect 6963 24021 6972 24055
rect 6920 24012 6972 24021
rect 7196 24012 7248 24064
rect 8392 24055 8444 24064
rect 8392 24021 8401 24055
rect 8401 24021 8435 24055
rect 8435 24021 8444 24055
rect 8392 24012 8444 24021
rect 9404 24012 9456 24064
rect 12440 24012 12492 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 4160 23851 4212 23860
rect 4160 23817 4169 23851
rect 4169 23817 4203 23851
rect 4203 23817 4212 23851
rect 4160 23808 4212 23817
rect 4528 23851 4580 23860
rect 4528 23817 4537 23851
rect 4537 23817 4571 23851
rect 4571 23817 4580 23851
rect 4528 23808 4580 23817
rect 4804 23851 4856 23860
rect 4804 23817 4813 23851
rect 4813 23817 4847 23851
rect 4847 23817 4856 23851
rect 4804 23808 4856 23817
rect 7288 23808 7340 23860
rect 7748 23808 7800 23860
rect 7932 23808 7984 23860
rect 10232 23808 10284 23860
rect 11336 23808 11388 23860
rect 8024 23740 8076 23792
rect 10140 23740 10192 23792
rect 11520 23740 11572 23792
rect 6920 23672 6972 23724
rect 7196 23647 7248 23656
rect 7196 23613 7205 23647
rect 7205 23613 7239 23647
rect 7239 23613 7248 23647
rect 7196 23604 7248 23613
rect 8668 23604 8720 23656
rect 9128 23647 9180 23656
rect 9128 23613 9137 23647
rect 9137 23613 9171 23647
rect 9171 23613 9180 23647
rect 9128 23604 9180 23613
rect 9404 23647 9456 23656
rect 9404 23613 9438 23647
rect 9438 23613 9456 23647
rect 9404 23604 9456 23613
rect 8116 23536 8168 23588
rect 5816 23511 5868 23520
rect 5816 23477 5825 23511
rect 5825 23477 5859 23511
rect 5859 23477 5868 23511
rect 5816 23468 5868 23477
rect 6828 23511 6880 23520
rect 6828 23477 6837 23511
rect 6837 23477 6871 23511
rect 6871 23477 6880 23511
rect 6828 23468 6880 23477
rect 9312 23468 9364 23520
rect 12348 23468 12400 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 6828 23264 6880 23316
rect 6920 23264 6972 23316
rect 8392 23264 8444 23316
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 12532 23264 12584 23316
rect 4436 23239 4488 23248
rect 4436 23205 4445 23239
rect 4445 23205 4479 23239
rect 4479 23205 4488 23239
rect 4436 23196 4488 23205
rect 7104 23196 7156 23248
rect 8300 23196 8352 23248
rect 8668 23196 8720 23248
rect 1676 23128 1728 23180
rect 4528 23171 4580 23180
rect 4528 23137 4537 23171
rect 4537 23137 4571 23171
rect 4571 23137 4580 23171
rect 4528 23128 4580 23137
rect 5816 23128 5868 23180
rect 7380 23128 7432 23180
rect 7656 23128 7708 23180
rect 8024 23128 8076 23180
rect 4620 23103 4672 23112
rect 4620 23069 4629 23103
rect 4629 23069 4663 23103
rect 4663 23069 4672 23103
rect 4620 23060 4672 23069
rect 6276 23103 6328 23112
rect 6276 23069 6285 23103
rect 6285 23069 6319 23103
rect 6319 23069 6328 23103
rect 6276 23060 6328 23069
rect 8300 23103 8352 23112
rect 8300 23069 8309 23103
rect 8309 23069 8343 23103
rect 8343 23069 8352 23103
rect 8300 23060 8352 23069
rect 12440 23128 12492 23180
rect 12808 23128 12860 23180
rect 9128 23060 9180 23112
rect 3148 22924 3200 22976
rect 5724 22967 5776 22976
rect 5724 22933 5733 22967
rect 5733 22933 5767 22967
rect 5767 22933 5776 22967
rect 5724 22924 5776 22933
rect 12348 22992 12400 23044
rect 11336 22924 11388 22976
rect 11980 22924 12032 22976
rect 13176 22967 13228 22976
rect 13176 22933 13185 22967
rect 13185 22933 13219 22967
rect 13219 22933 13228 22967
rect 13176 22924 13228 22933
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2412 22720 2464 22772
rect 2688 22763 2740 22772
rect 1676 22695 1728 22704
rect 1676 22661 1685 22695
rect 1685 22661 1719 22695
rect 1719 22661 1728 22695
rect 1676 22652 1728 22661
rect 2688 22729 2697 22763
rect 2697 22729 2731 22763
rect 2731 22729 2740 22763
rect 2688 22720 2740 22729
rect 4436 22720 4488 22772
rect 4620 22720 4672 22772
rect 6276 22763 6328 22772
rect 6276 22729 6285 22763
rect 6285 22729 6319 22763
rect 6319 22729 6328 22763
rect 6276 22720 6328 22729
rect 7932 22720 7984 22772
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 7748 22652 7800 22704
rect 4068 22584 4120 22636
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 7656 22627 7708 22636
rect 7656 22593 7665 22627
rect 7665 22593 7699 22627
rect 7699 22593 7708 22627
rect 7656 22584 7708 22593
rect 8392 22720 8444 22772
rect 10508 22720 10560 22772
rect 8668 22652 8720 22704
rect 10784 22584 10836 22636
rect 5356 22516 5408 22568
rect 7840 22516 7892 22568
rect 8668 22516 8720 22568
rect 5908 22448 5960 22500
rect 9772 22448 9824 22500
rect 10048 22448 10100 22500
rect 11336 22720 11388 22772
rect 11520 22720 11572 22772
rect 12256 22720 12308 22772
rect 12532 22720 12584 22772
rect 12164 22448 12216 22500
rect 12900 22584 12952 22636
rect 12992 22584 13044 22636
rect 13176 22584 13228 22636
rect 12808 22516 12860 22568
rect 2412 22380 2464 22432
rect 8760 22380 8812 22432
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 10140 22380 10192 22389
rect 10876 22380 10928 22432
rect 12348 22380 12400 22432
rect 13084 22448 13136 22500
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 2412 22219 2464 22228
rect 2412 22185 2421 22219
rect 2421 22185 2455 22219
rect 2455 22185 2464 22219
rect 2412 22176 2464 22185
rect 2504 22176 2556 22228
rect 3056 22176 3108 22228
rect 3424 22176 3476 22228
rect 5908 22176 5960 22228
rect 7472 22176 7524 22228
rect 10692 22176 10744 22228
rect 2964 22108 3016 22160
rect 1676 22040 1728 22092
rect 4620 22083 4672 22092
rect 4620 22049 4629 22083
rect 4629 22049 4663 22083
rect 4663 22049 4672 22083
rect 4620 22040 4672 22049
rect 3056 22015 3108 22024
rect 3056 21981 3065 22015
rect 3065 21981 3099 22015
rect 3099 21981 3108 22015
rect 3056 21972 3108 21981
rect 5356 22108 5408 22160
rect 5080 22083 5132 22092
rect 5080 22049 5114 22083
rect 5114 22049 5132 22083
rect 5080 22040 5132 22049
rect 6092 22040 6144 22092
rect 6736 22040 6788 22092
rect 7656 22083 7708 22092
rect 7656 22049 7665 22083
rect 7665 22049 7699 22083
rect 7699 22049 7708 22083
rect 7656 22040 7708 22049
rect 7748 22083 7800 22092
rect 7748 22049 7757 22083
rect 7757 22049 7791 22083
rect 7791 22049 7800 22083
rect 7748 22040 7800 22049
rect 8024 22040 8076 22092
rect 8300 22040 8352 22092
rect 10140 22108 10192 22160
rect 10232 22108 10284 22160
rect 10784 22151 10836 22160
rect 8116 21972 8168 22024
rect 1584 21947 1636 21956
rect 1584 21913 1593 21947
rect 1593 21913 1627 21947
rect 1627 21913 1636 21947
rect 1584 21904 1636 21913
rect 7380 21904 7432 21956
rect 4252 21836 4304 21888
rect 8760 21836 8812 21888
rect 9772 21836 9824 21888
rect 10784 22117 10793 22151
rect 10793 22117 10827 22151
rect 10827 22117 10836 22151
rect 10784 22108 10836 22117
rect 10692 21972 10744 22024
rect 11060 22176 11112 22228
rect 11980 22176 12032 22228
rect 12808 22219 12860 22228
rect 12808 22185 12817 22219
rect 12817 22185 12851 22219
rect 12851 22185 12860 22219
rect 12808 22176 12860 22185
rect 12348 22040 12400 22092
rect 11336 21972 11388 22024
rect 12440 21972 12492 22024
rect 10324 21836 10376 21888
rect 11336 21836 11388 21888
rect 13084 21836 13136 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 2688 21632 2740 21684
rect 4068 21675 4120 21684
rect 4068 21641 4077 21675
rect 4077 21641 4111 21675
rect 4111 21641 4120 21675
rect 4068 21632 4120 21641
rect 4252 21632 4304 21684
rect 4528 21632 4580 21684
rect 5908 21632 5960 21684
rect 7472 21632 7524 21684
rect 8208 21632 8260 21684
rect 2504 21607 2556 21616
rect 2504 21573 2513 21607
rect 2513 21573 2547 21607
rect 2547 21573 2556 21607
rect 2504 21564 2556 21573
rect 10324 21564 10376 21616
rect 10692 21632 10744 21684
rect 11244 21632 11296 21684
rect 11520 21632 11572 21684
rect 11888 21632 11940 21684
rect 11152 21496 11204 21548
rect 11336 21539 11388 21548
rect 11336 21505 11345 21539
rect 11345 21505 11379 21539
rect 11379 21505 11388 21539
rect 11336 21496 11388 21505
rect 12992 21539 13044 21548
rect 2688 21471 2740 21480
rect 2688 21437 2697 21471
rect 2697 21437 2731 21471
rect 2731 21437 2740 21471
rect 2688 21428 2740 21437
rect 3056 21360 3108 21412
rect 5356 21428 5408 21480
rect 7564 21428 7616 21480
rect 10048 21428 10100 21480
rect 10324 21428 10376 21480
rect 10508 21471 10560 21480
rect 10508 21437 10517 21471
rect 10517 21437 10551 21471
rect 10551 21437 10560 21471
rect 10508 21428 10560 21437
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 5356 21292 5408 21344
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 5540 21292 5592 21301
rect 7288 21360 7340 21412
rect 9312 21360 9364 21412
rect 5908 21292 5960 21344
rect 7656 21292 7708 21344
rect 8116 21292 8168 21344
rect 10600 21335 10652 21344
rect 10600 21301 10609 21335
rect 10609 21301 10643 21335
rect 10643 21301 10652 21335
rect 10600 21292 10652 21301
rect 11520 21292 11572 21344
rect 13360 21292 13412 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 2688 21131 2740 21140
rect 2688 21097 2697 21131
rect 2697 21097 2731 21131
rect 2731 21097 2740 21131
rect 2688 21088 2740 21097
rect 3056 21131 3108 21140
rect 3056 21097 3065 21131
rect 3065 21097 3099 21131
rect 3099 21097 3108 21131
rect 3056 21088 3108 21097
rect 5080 21088 5132 21140
rect 6184 21088 6236 21140
rect 7564 21088 7616 21140
rect 8024 21088 8076 21140
rect 9404 21131 9456 21140
rect 9404 21097 9413 21131
rect 9413 21097 9447 21131
rect 9447 21097 9456 21131
rect 9404 21088 9456 21097
rect 10508 21131 10560 21140
rect 10508 21097 10517 21131
rect 10517 21097 10551 21131
rect 10551 21097 10560 21131
rect 10508 21088 10560 21097
rect 11060 21131 11112 21140
rect 11060 21097 11069 21131
rect 11069 21097 11103 21131
rect 11103 21097 11112 21131
rect 11060 21088 11112 21097
rect 11520 21088 11572 21140
rect 12992 21088 13044 21140
rect 5540 21020 5592 21072
rect 5632 20995 5684 21004
rect 5632 20961 5666 20995
rect 5666 20961 5684 20995
rect 7656 20995 7708 21004
rect 5632 20952 5684 20961
rect 7656 20961 7665 20995
rect 7665 20961 7699 20995
rect 7699 20961 7708 20995
rect 7656 20952 7708 20961
rect 8208 20995 8260 21004
rect 8208 20961 8217 20995
rect 8217 20961 8251 20995
rect 8251 20961 8260 20995
rect 8208 20952 8260 20961
rect 1676 20927 1728 20936
rect 1676 20893 1685 20927
rect 1685 20893 1719 20927
rect 1719 20893 1728 20927
rect 1676 20884 1728 20893
rect 5356 20927 5408 20936
rect 5356 20893 5365 20927
rect 5365 20893 5399 20927
rect 5399 20893 5408 20927
rect 5356 20884 5408 20893
rect 7748 20884 7800 20936
rect 9772 21020 9824 21072
rect 11336 21020 11388 21072
rect 9220 20952 9272 21004
rect 9404 20952 9456 21004
rect 11152 20952 11204 21004
rect 11428 20952 11480 21004
rect 13084 20952 13136 21004
rect 13268 20952 13320 21004
rect 8668 20884 8720 20936
rect 9588 20884 9640 20936
rect 11796 20927 11848 20936
rect 11796 20893 11805 20927
rect 11805 20893 11839 20927
rect 11839 20893 11848 20927
rect 11796 20884 11848 20893
rect 7840 20791 7892 20800
rect 7840 20757 7849 20791
rect 7849 20757 7883 20791
rect 7883 20757 7892 20791
rect 7840 20748 7892 20757
rect 13176 20791 13228 20800
rect 13176 20757 13185 20791
rect 13185 20757 13219 20791
rect 13219 20757 13228 20791
rect 13176 20748 13228 20757
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 5632 20544 5684 20596
rect 7840 20544 7892 20596
rect 8208 20587 8260 20596
rect 8208 20553 8217 20587
rect 8217 20553 8251 20587
rect 8251 20553 8260 20587
rect 8208 20544 8260 20553
rect 11796 20544 11848 20596
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 11336 20476 11388 20528
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 7748 20204 7800 20256
rect 8300 20204 8352 20256
rect 13176 20340 13228 20392
rect 9496 20272 9548 20324
rect 12900 20315 12952 20324
rect 12900 20281 12909 20315
rect 12909 20281 12943 20315
rect 12943 20281 12952 20315
rect 12900 20272 12952 20281
rect 11428 20204 11480 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 7564 20000 7616 20052
rect 10048 20043 10100 20052
rect 10048 20009 10057 20043
rect 10057 20009 10091 20043
rect 10091 20009 10100 20043
rect 10048 20000 10100 20009
rect 10508 20043 10560 20052
rect 10508 20009 10517 20043
rect 10517 20009 10551 20043
rect 10551 20009 10560 20043
rect 10508 20000 10560 20009
rect 12992 20043 13044 20052
rect 12992 20009 13001 20043
rect 13001 20009 13035 20043
rect 13035 20009 13044 20043
rect 12992 20000 13044 20009
rect 11980 19932 12032 19984
rect 10048 19864 10100 19916
rect 10968 19864 11020 19916
rect 11244 19864 11296 19916
rect 11152 19796 11204 19848
rect 7288 19660 7340 19712
rect 8852 19660 8904 19712
rect 9496 19660 9548 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 11244 19456 11296 19508
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 11152 19363 11204 19372
rect 8024 19252 8076 19304
rect 8208 19252 8260 19304
rect 8392 19252 8444 19304
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 9864 19252 9916 19304
rect 10692 19252 10744 19304
rect 6644 19184 6696 19236
rect 10600 19184 10652 19236
rect 10784 19184 10836 19236
rect 11520 19227 11572 19236
rect 11520 19193 11529 19227
rect 11529 19193 11563 19227
rect 11563 19193 11572 19227
rect 11520 19184 11572 19193
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 7196 19159 7248 19168
rect 6828 19116 6880 19125
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7288 19116 7340 19125
rect 8300 19116 8352 19168
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 9036 19116 9088 19168
rect 9588 19116 9640 19168
rect 9864 19116 9916 19168
rect 10048 19116 10100 19168
rect 10508 19159 10560 19168
rect 10508 19125 10517 19159
rect 10517 19125 10551 19159
rect 10551 19125 10560 19159
rect 10508 19116 10560 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 6644 18912 6696 18964
rect 7196 18912 7248 18964
rect 10324 18912 10376 18964
rect 10692 18955 10744 18964
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 11152 18955 11204 18964
rect 11152 18921 11161 18955
rect 11161 18921 11195 18955
rect 11195 18921 11204 18955
rect 11152 18912 11204 18921
rect 11980 18912 12032 18964
rect 5264 18776 5316 18828
rect 5448 18819 5500 18828
rect 5448 18785 5482 18819
rect 5482 18785 5500 18819
rect 5448 18776 5500 18785
rect 8208 18819 8260 18828
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 9864 18776 9916 18828
rect 10600 18776 10652 18828
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 7656 18640 7708 18692
rect 9496 18640 9548 18692
rect 9864 18640 9916 18692
rect 10968 18708 11020 18760
rect 10876 18640 10928 18692
rect 6184 18572 6236 18624
rect 7840 18615 7892 18624
rect 7840 18581 7849 18615
rect 7849 18581 7883 18615
rect 7883 18581 7892 18615
rect 7840 18572 7892 18581
rect 9680 18615 9732 18624
rect 9680 18581 9689 18615
rect 9689 18581 9723 18615
rect 9723 18581 9732 18615
rect 9680 18572 9732 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 8300 18368 8352 18420
rect 9496 18411 9548 18420
rect 9496 18377 9505 18411
rect 9505 18377 9539 18411
rect 9539 18377 9548 18411
rect 9496 18368 9548 18377
rect 10324 18368 10376 18420
rect 7656 18343 7708 18352
rect 7656 18309 7665 18343
rect 7665 18309 7699 18343
rect 7699 18309 7708 18343
rect 7656 18300 7708 18309
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 5356 18232 5408 18284
rect 5908 18232 5960 18284
rect 8024 18164 8076 18216
rect 3884 18139 3936 18148
rect 3884 18105 3918 18139
rect 3918 18105 3936 18139
rect 3884 18096 3936 18105
rect 3516 18071 3568 18080
rect 3516 18037 3525 18071
rect 3525 18037 3559 18071
rect 3559 18037 3568 18071
rect 3516 18028 3568 18037
rect 4068 18028 4120 18080
rect 5448 18096 5500 18148
rect 8392 18139 8444 18148
rect 8392 18105 8426 18139
rect 8426 18105 8444 18139
rect 8392 18096 8444 18105
rect 8300 18028 8352 18080
rect 9864 18028 9916 18080
rect 10968 18028 11020 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 7472 17824 7524 17876
rect 9680 17824 9732 17876
rect 11152 17824 11204 17876
rect 6184 17756 6236 17808
rect 11980 17756 12032 17808
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 4896 17731 4948 17740
rect 4896 17697 4905 17731
rect 4905 17697 4939 17731
rect 4939 17697 4948 17731
rect 4896 17688 4948 17697
rect 5724 17688 5776 17740
rect 6092 17688 6144 17740
rect 9772 17688 9824 17740
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 5908 17620 5960 17672
rect 8208 17620 8260 17672
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 11428 17620 11480 17672
rect 3884 17552 3936 17604
rect 3976 17484 4028 17536
rect 8024 17484 8076 17536
rect 8392 17552 8444 17604
rect 9680 17595 9732 17604
rect 9680 17561 9689 17595
rect 9689 17561 9723 17595
rect 9723 17561 9732 17595
rect 9680 17552 9732 17561
rect 9496 17484 9548 17536
rect 13176 17527 13228 17536
rect 13176 17493 13185 17527
rect 13185 17493 13219 17527
rect 13219 17493 13228 17527
rect 13176 17484 13228 17493
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 4804 17280 4856 17332
rect 10324 17280 10376 17332
rect 11152 17323 11204 17332
rect 11152 17289 11161 17323
rect 11161 17289 11195 17323
rect 11195 17289 11204 17323
rect 11152 17280 11204 17289
rect 11980 17280 12032 17332
rect 6184 17212 6236 17264
rect 3516 17119 3568 17128
rect 3516 17085 3525 17119
rect 3525 17085 3559 17119
rect 3559 17085 3568 17119
rect 3516 17076 3568 17085
rect 5908 17144 5960 17196
rect 6644 17144 6696 17196
rect 6828 17144 6880 17196
rect 8300 17212 8352 17264
rect 8668 17212 8720 17264
rect 5816 17076 5868 17128
rect 8392 17076 8444 17128
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 9496 17119 9548 17128
rect 9496 17085 9530 17119
rect 9530 17085 9548 17119
rect 9496 17076 9548 17085
rect 4252 17008 4304 17060
rect 4620 16940 4672 16992
rect 4988 16983 5040 16992
rect 4988 16949 4997 16983
rect 4997 16949 5031 16983
rect 5031 16949 5040 16983
rect 4988 16940 5040 16949
rect 5908 16940 5960 16992
rect 6736 17008 6788 17060
rect 7472 17008 7524 17060
rect 9772 17008 9824 17060
rect 6920 16940 6972 16992
rect 8484 16940 8536 16992
rect 9496 16940 9548 16992
rect 11428 16940 11480 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 4896 16779 4948 16788
rect 4896 16745 4905 16779
rect 4905 16745 4939 16779
rect 4939 16745 4948 16779
rect 4896 16736 4948 16745
rect 6184 16736 6236 16788
rect 7288 16736 7340 16788
rect 7656 16779 7708 16788
rect 7656 16745 7665 16779
rect 7665 16745 7699 16779
rect 7699 16745 7708 16779
rect 7656 16736 7708 16745
rect 8668 16736 8720 16788
rect 9312 16736 9364 16788
rect 5540 16668 5592 16720
rect 9588 16668 9640 16720
rect 10324 16736 10376 16788
rect 10968 16736 11020 16788
rect 4344 16600 4396 16652
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 7748 16575 7800 16584
rect 7748 16541 7757 16575
rect 7757 16541 7791 16575
rect 7791 16541 7800 16575
rect 7748 16532 7800 16541
rect 9220 16600 9272 16652
rect 11428 16668 11480 16720
rect 10784 16643 10836 16652
rect 10784 16609 10818 16643
rect 10818 16609 10836 16643
rect 10784 16600 10836 16609
rect 8392 16532 8444 16584
rect 4252 16396 4304 16448
rect 4620 16396 4672 16448
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 10784 16396 10836 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 7196 16235 7248 16244
rect 7196 16201 7205 16235
rect 7205 16201 7239 16235
rect 7239 16201 7248 16235
rect 7196 16192 7248 16201
rect 7288 16192 7340 16244
rect 7564 16192 7616 16244
rect 8392 16192 8444 16244
rect 8760 16235 8812 16244
rect 8760 16201 8769 16235
rect 8769 16201 8803 16235
rect 8803 16201 8812 16235
rect 8760 16192 8812 16201
rect 8852 16192 8904 16244
rect 1952 16099 2004 16108
rect 1952 16065 1961 16099
rect 1961 16065 1995 16099
rect 1995 16065 2004 16099
rect 1952 16056 2004 16065
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 6828 16056 6880 16108
rect 7288 16056 7340 16108
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 10232 16192 10284 16244
rect 10600 16192 10652 16244
rect 10324 16167 10376 16176
rect 10324 16133 10333 16167
rect 10333 16133 10367 16167
rect 10367 16133 10376 16167
rect 10324 16124 10376 16133
rect 3976 15988 4028 16040
rect 9404 15988 9456 16040
rect 5540 15920 5592 15972
rect 7564 15963 7616 15972
rect 7564 15929 7573 15963
rect 7573 15929 7607 15963
rect 7607 15929 7616 15963
rect 7564 15920 7616 15929
rect 8852 15920 8904 15972
rect 9312 15920 9364 15972
rect 9588 16056 9640 16108
rect 10876 16099 10928 16108
rect 10876 16065 10885 16099
rect 10885 16065 10919 16099
rect 10919 16065 10928 16099
rect 10876 16056 10928 16065
rect 10692 15963 10744 15972
rect 10692 15929 10701 15963
rect 10701 15929 10735 15963
rect 10735 15929 10744 15963
rect 10692 15920 10744 15929
rect 2780 15852 2832 15904
rect 3884 15852 3936 15904
rect 4068 15852 4120 15904
rect 4252 15852 4304 15904
rect 4712 15852 4764 15904
rect 5080 15852 5132 15904
rect 5632 15852 5684 15904
rect 7472 15852 7524 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 11428 15895 11480 15904
rect 11428 15861 11437 15895
rect 11437 15861 11471 15895
rect 11471 15861 11480 15895
rect 11428 15852 11480 15861
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 6184 15648 6236 15700
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 4252 15444 4304 15496
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 7288 15648 7340 15700
rect 7564 15648 7616 15700
rect 7656 15691 7708 15700
rect 7656 15657 7665 15691
rect 7665 15657 7699 15691
rect 7699 15657 7708 15691
rect 8852 15691 8904 15700
rect 7656 15648 7708 15657
rect 8852 15657 8861 15691
rect 8861 15657 8895 15691
rect 8895 15657 8904 15691
rect 8852 15648 8904 15657
rect 10876 15648 10928 15700
rect 12348 15580 12400 15632
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 8392 15512 8444 15564
rect 8852 15512 8904 15564
rect 7748 15487 7800 15496
rect 4620 15444 4672 15453
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 9588 15444 9640 15496
rect 12256 15444 12308 15496
rect 4068 15376 4120 15428
rect 12900 15376 12952 15428
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 12992 15351 13044 15360
rect 12992 15317 13001 15351
rect 13001 15317 13035 15351
rect 13035 15317 13044 15351
rect 12992 15308 13044 15317
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 4252 15104 4304 15156
rect 7656 15104 7708 15156
rect 7932 15104 7984 15156
rect 10692 15104 10744 15156
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 4068 15036 4120 15088
rect 11152 15036 11204 15088
rect 12716 15104 12768 15156
rect 12900 15104 12952 15156
rect 5172 14968 5224 15020
rect 7196 14968 7248 15020
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 8392 14968 8444 15020
rect 9312 14968 9364 15020
rect 10876 14968 10928 15020
rect 11980 14968 12032 15020
rect 12440 14968 12492 15020
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 4436 14832 4488 14884
rect 4620 14875 4672 14884
rect 4620 14841 4629 14875
rect 4629 14841 4663 14875
rect 4663 14841 4672 14875
rect 4620 14832 4672 14841
rect 9680 14900 9732 14952
rect 10416 14900 10468 14952
rect 11244 14900 11296 14952
rect 11888 14900 11940 14952
rect 12164 14900 12216 14952
rect 9588 14832 9640 14884
rect 2688 14764 2740 14816
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 5356 14764 5408 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7012 14764 7064 14816
rect 9312 14764 9364 14816
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 11060 14764 11112 14816
rect 13728 14832 13780 14884
rect 12716 14764 12768 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 4436 14560 4488 14612
rect 4804 14560 4856 14612
rect 6828 14560 6880 14612
rect 7564 14560 7616 14612
rect 7748 14560 7800 14612
rect 8208 14560 8260 14612
rect 9588 14560 9640 14612
rect 10784 14560 10836 14612
rect 11244 14603 11296 14612
rect 11244 14569 11253 14603
rect 11253 14569 11287 14603
rect 11287 14569 11296 14603
rect 11244 14560 11296 14569
rect 11980 14560 12032 14612
rect 6644 14535 6696 14544
rect 6644 14501 6653 14535
rect 6653 14501 6687 14535
rect 6687 14501 6696 14535
rect 6644 14492 6696 14501
rect 12164 14492 12216 14544
rect 4988 14424 5040 14476
rect 9312 14424 9364 14476
rect 10324 14424 10376 14476
rect 10968 14424 11020 14476
rect 4712 14356 4764 14408
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 7564 14356 7616 14408
rect 7932 14356 7984 14408
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 8760 14356 8812 14408
rect 10416 14356 10468 14408
rect 10876 14399 10928 14408
rect 10876 14365 10885 14399
rect 10885 14365 10919 14399
rect 10919 14365 10928 14399
rect 10876 14356 10928 14365
rect 11428 14356 11480 14408
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 7472 14288 7524 14340
rect 7656 14288 7708 14340
rect 3332 14220 3384 14272
rect 5632 14220 5684 14272
rect 12164 14220 12216 14272
rect 12440 14220 12492 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 6828 14016 6880 14068
rect 8024 14016 8076 14068
rect 8208 14016 8260 14068
rect 8760 14016 8812 14068
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 11980 14016 12032 14068
rect 5172 13948 5224 14000
rect 6644 13991 6696 14000
rect 6644 13957 6653 13991
rect 6653 13957 6687 13991
rect 6687 13957 6696 13991
rect 6644 13948 6696 13957
rect 10600 13948 10652 14000
rect 12440 14016 12492 14068
rect 2320 13812 2372 13864
rect 4988 13855 5040 13864
rect 3332 13744 3384 13796
rect 4988 13821 4997 13855
rect 4997 13821 5031 13855
rect 5031 13821 5040 13855
rect 4988 13812 5040 13821
rect 5540 13812 5592 13864
rect 6736 13812 6788 13864
rect 4896 13744 4948 13796
rect 7104 13744 7156 13796
rect 7932 13812 7984 13864
rect 8392 13812 8444 13864
rect 10600 13812 10652 13864
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 10968 13744 11020 13796
rect 12348 13744 12400 13796
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 2688 13472 2740 13524
rect 4804 13472 4856 13524
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 8484 13472 8536 13524
rect 9312 13472 9364 13524
rect 10876 13472 10928 13524
rect 12072 13515 12124 13524
rect 12072 13481 12081 13515
rect 12081 13481 12115 13515
rect 12115 13481 12124 13515
rect 12072 13472 12124 13481
rect 1768 13404 1820 13456
rect 4252 13404 4304 13456
rect 5172 13447 5224 13456
rect 5172 13413 5206 13447
rect 5206 13413 5224 13447
rect 5172 13404 5224 13413
rect 8208 13404 8260 13456
rect 1676 13336 1728 13388
rect 3056 13336 3108 13388
rect 6920 13336 6972 13388
rect 8024 13336 8076 13388
rect 10232 13336 10284 13388
rect 10784 13336 10836 13388
rect 2596 13268 2648 13320
rect 4712 13268 4764 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 8392 13200 8444 13252
rect 10324 13268 10376 13320
rect 10508 13200 10560 13252
rect 11520 13268 11572 13320
rect 11888 13268 11940 13320
rect 12440 13268 12492 13320
rect 11060 13200 11112 13252
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 1768 12971 1820 12980
rect 1768 12937 1777 12971
rect 1777 12937 1811 12971
rect 1811 12937 1820 12971
rect 1768 12928 1820 12937
rect 4344 12928 4396 12980
rect 5172 12928 5224 12980
rect 7380 12928 7432 12980
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 9864 12928 9916 12980
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 10508 12928 10560 12937
rect 11520 12928 11572 12980
rect 12072 12928 12124 12980
rect 12440 12928 12492 12980
rect 6828 12903 6880 12912
rect 6828 12869 6837 12903
rect 6837 12869 6871 12903
rect 6871 12869 6880 12903
rect 6828 12860 6880 12869
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 8392 12860 8444 12912
rect 10692 12792 10744 12844
rect 11888 12792 11940 12844
rect 2320 12724 2372 12776
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 6920 12724 6972 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 2504 12699 2556 12708
rect 2504 12665 2538 12699
rect 2538 12665 2556 12699
rect 2504 12656 2556 12665
rect 4896 12656 4948 12708
rect 2872 12588 2924 12640
rect 3332 12588 3384 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 5632 12656 5684 12708
rect 6092 12656 6144 12708
rect 7104 12588 7156 12640
rect 9312 12656 9364 12708
rect 9680 12588 9732 12640
rect 10784 12588 10836 12640
rect 12072 12588 12124 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 5816 12384 5868 12436
rect 6000 12384 6052 12436
rect 6920 12427 6972 12436
rect 6920 12393 6929 12427
rect 6929 12393 6963 12427
rect 6963 12393 6972 12427
rect 6920 12384 6972 12393
rect 7104 12384 7156 12436
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 9312 12384 9364 12436
rect 10324 12384 10376 12436
rect 5448 12316 5500 12368
rect 6184 12316 6236 12368
rect 6828 12316 6880 12368
rect 5172 12248 5224 12300
rect 5356 12248 5408 12300
rect 6000 12223 6052 12232
rect 6000 12189 6009 12223
rect 6009 12189 6043 12223
rect 6043 12189 6052 12223
rect 6000 12180 6052 12189
rect 6092 12180 6144 12232
rect 6736 12180 6788 12232
rect 7472 12316 7524 12368
rect 9680 12316 9732 12368
rect 10968 12384 11020 12436
rect 12440 12384 12492 12436
rect 9772 12248 9824 12300
rect 10140 12248 10192 12300
rect 10508 12316 10560 12368
rect 10784 12291 10836 12300
rect 10784 12257 10818 12291
rect 10818 12257 10836 12291
rect 10784 12248 10836 12257
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 2504 12112 2556 12164
rect 3516 12112 3568 12164
rect 3056 12087 3108 12096
rect 3056 12053 3065 12087
rect 3065 12053 3099 12087
rect 3099 12053 3108 12087
rect 3056 12044 3108 12053
rect 5264 12044 5316 12096
rect 10416 12044 10468 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 3516 11840 3568 11892
rect 4252 11840 4304 11892
rect 6092 11840 6144 11892
rect 10508 11883 10560 11892
rect 10508 11849 10517 11883
rect 10517 11849 10551 11883
rect 10551 11849 10560 11883
rect 10508 11840 10560 11849
rect 10784 11840 10836 11892
rect 4344 11815 4396 11824
rect 4344 11781 4353 11815
rect 4353 11781 4387 11815
rect 4387 11781 4396 11815
rect 4344 11772 4396 11781
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 2044 11568 2096 11620
rect 5080 11568 5132 11620
rect 5448 11636 5500 11688
rect 6092 11636 6144 11688
rect 7380 11636 7432 11688
rect 5448 11500 5500 11552
rect 10692 11568 10744 11620
rect 7472 11500 7524 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 3056 11296 3108 11348
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 6000 11296 6052 11348
rect 7196 11296 7248 11348
rect 4988 11228 5040 11280
rect 5448 11228 5500 11280
rect 6184 11271 6236 11280
rect 6184 11237 6193 11271
rect 6193 11237 6227 11271
rect 6227 11237 6236 11271
rect 6184 11228 6236 11237
rect 7472 11271 7524 11280
rect 7472 11237 7481 11271
rect 7481 11237 7515 11271
rect 7515 11237 7524 11271
rect 7472 11228 7524 11237
rect 5816 11160 5868 11212
rect 6460 11160 6512 11212
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 2044 10956 2096 11008
rect 3424 10999 3476 11008
rect 3424 10965 3433 10999
rect 3433 10965 3467 10999
rect 3467 10965 3476 10999
rect 3424 10956 3476 10965
rect 7380 11092 7432 11144
rect 7012 10956 7064 11008
rect 8116 10956 8168 11008
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 12532 10956 12584 10965
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 3516 10752 3568 10804
rect 5264 10752 5316 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 6092 10795 6144 10804
rect 6092 10761 6101 10795
rect 6101 10761 6135 10795
rect 6135 10761 6144 10795
rect 6092 10752 6144 10761
rect 2872 10616 2924 10668
rect 1860 10548 1912 10600
rect 3424 10616 3476 10668
rect 4988 10684 5040 10736
rect 12532 10616 12584 10668
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 3700 10523 3752 10532
rect 3700 10489 3709 10523
rect 3709 10489 3743 10523
rect 3743 10489 3752 10523
rect 3700 10480 3752 10489
rect 6460 10523 6512 10532
rect 6460 10489 6469 10523
rect 6469 10489 6503 10523
rect 6503 10489 6512 10523
rect 6460 10480 6512 10489
rect 12256 10523 12308 10532
rect 12256 10489 12265 10523
rect 12265 10489 12299 10523
rect 12299 10489 12308 10523
rect 12256 10480 12308 10489
rect 14096 10480 14148 10532
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 2412 10412 2464 10464
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 8024 10412 8076 10464
rect 12532 10412 12584 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 3700 10208 3752 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 12900 10208 12952 10260
rect 2872 10140 2924 10192
rect 4712 10115 4764 10124
rect 4712 10081 4721 10115
rect 4721 10081 4755 10115
rect 4755 10081 4764 10115
rect 4712 10072 4764 10081
rect 2412 10004 2464 10056
rect 2780 9936 2832 9988
rect 3516 10004 3568 10056
rect 4252 10004 4304 10056
rect 5632 10072 5684 10124
rect 7288 10072 7340 10124
rect 7932 10072 7984 10124
rect 8484 10072 8536 10124
rect 10508 10072 10560 10124
rect 10692 10115 10744 10124
rect 10692 10081 10726 10115
rect 10726 10081 10744 10115
rect 10692 10072 10744 10081
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13636 10072 13688 10124
rect 13452 10047 13504 10056
rect 4436 9936 4488 9988
rect 8024 9936 8076 9988
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 13544 9936 13596 9988
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 7472 9868 7524 9920
rect 9312 9868 9364 9920
rect 11980 9868 12032 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 3424 9664 3476 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 4528 9664 4580 9716
rect 10508 9664 10560 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 13268 9664 13320 9716
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 3056 9528 3108 9580
rect 12532 9596 12584 9648
rect 5540 9528 5592 9580
rect 8024 9528 8076 9580
rect 11980 9528 12032 9580
rect 13268 9528 13320 9580
rect 1768 9460 1820 9512
rect 2320 9460 2372 9512
rect 3424 9460 3476 9512
rect 4252 9460 4304 9512
rect 5816 9460 5868 9512
rect 7380 9460 7432 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 10508 9460 10560 9512
rect 12440 9460 12492 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 3332 9435 3384 9444
rect 3332 9401 3341 9435
rect 3341 9401 3375 9435
rect 3375 9401 3384 9435
rect 3332 9392 3384 9401
rect 4436 9392 4488 9444
rect 5724 9392 5776 9444
rect 3516 9324 3568 9376
rect 4712 9324 4764 9376
rect 5540 9324 5592 9376
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 8484 9392 8536 9444
rect 8300 9324 8352 9376
rect 8576 9324 8628 9376
rect 9312 9392 9364 9444
rect 10048 9392 10100 9444
rect 10692 9392 10744 9444
rect 9496 9324 9548 9376
rect 10232 9367 10284 9376
rect 10232 9333 10241 9367
rect 10241 9333 10275 9367
rect 10275 9333 10284 9367
rect 10232 9324 10284 9333
rect 12532 9324 12584 9376
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 5540 9120 5592 9172
rect 7380 9120 7432 9172
rect 10968 9120 11020 9172
rect 12624 9120 12676 9172
rect 13452 9120 13504 9172
rect 13636 9163 13688 9172
rect 13636 9129 13645 9163
rect 13645 9129 13679 9163
rect 13679 9129 13688 9163
rect 13636 9120 13688 9129
rect 2872 9052 2924 9104
rect 2688 8984 2740 9036
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 4528 9052 4580 9104
rect 6000 9052 6052 9104
rect 8116 9052 8168 9104
rect 11980 9095 12032 9104
rect 11980 9061 12014 9095
rect 12014 9061 12032 9095
rect 11980 9052 12032 9061
rect 2780 8984 2832 8993
rect 4344 9027 4396 9036
rect 4344 8993 4378 9027
rect 4378 8993 4396 9027
rect 4344 8984 4396 8993
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 8300 8916 8352 8968
rect 8208 8848 8260 8900
rect 10232 8916 10284 8968
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 10784 8916 10836 8968
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 3516 8780 3568 8832
rect 9588 8780 9640 8832
rect 13636 8848 13688 8900
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 1768 8576 1820 8628
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 2780 8576 2832 8628
rect 2872 8576 2924 8628
rect 7288 8576 7340 8628
rect 8852 8576 8904 8628
rect 10968 8619 11020 8628
rect 8300 8508 8352 8560
rect 4712 8440 4764 8492
rect 4344 8372 4396 8424
rect 6920 8372 6972 8424
rect 8760 8372 8812 8424
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 11980 8576 12032 8628
rect 10692 8551 10744 8560
rect 10692 8517 10701 8551
rect 10701 8517 10735 8551
rect 10735 8517 10744 8551
rect 10692 8508 10744 8517
rect 11888 8508 11940 8560
rect 10048 8440 10100 8492
rect 12808 8576 12860 8628
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 12440 8372 12492 8424
rect 4068 8304 4120 8356
rect 4712 8347 4764 8356
rect 4712 8313 4721 8347
rect 4721 8313 4755 8347
rect 4755 8313 4764 8347
rect 4712 8304 4764 8313
rect 6644 8347 6696 8356
rect 6644 8313 6653 8347
rect 6653 8313 6687 8347
rect 6687 8313 6696 8347
rect 6644 8304 6696 8313
rect 8024 8304 8076 8356
rect 9312 8304 9364 8356
rect 10140 8304 10192 8356
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 4528 8236 4580 8288
rect 7656 8236 7708 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 2872 8032 2924 8084
rect 6920 8032 6972 8084
rect 8392 8032 8444 8084
rect 10508 8032 10560 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 8300 7964 8352 8016
rect 10232 7964 10284 8016
rect 12992 8032 13044 8084
rect 5816 7896 5868 7948
rect 8208 7896 8260 7948
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 4068 7828 4120 7880
rect 4528 7828 4580 7880
rect 8116 7828 8168 7880
rect 8760 7828 8812 7880
rect 10048 7828 10100 7880
rect 10232 7828 10284 7880
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 6184 7760 6236 7812
rect 8300 7760 8352 7812
rect 5448 7692 5500 7744
rect 6092 7692 6144 7744
rect 9404 7692 9456 7744
rect 9680 7692 9732 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5632 7488 5684 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8392 7531 8444 7540
rect 8116 7488 8168 7497
rect 2044 7420 2096 7472
rect 6184 7420 6236 7472
rect 6736 7420 6788 7472
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 9680 7488 9732 7540
rect 10968 7488 11020 7540
rect 13820 7488 13872 7540
rect 15752 7488 15804 7540
rect 8668 7420 8720 7472
rect 10876 7420 10928 7472
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 5172 7284 5224 7336
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 5448 7216 5500 7268
rect 6828 7352 6880 7404
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 10048 7395 10100 7404
rect 10048 7361 10057 7395
rect 10057 7361 10091 7395
rect 10091 7361 10100 7395
rect 10048 7352 10100 7361
rect 7288 7284 7340 7336
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 6644 7216 6696 7268
rect 9956 7216 10008 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 6920 7148 6972 7200
rect 9680 7148 9732 7200
rect 10048 7148 10100 7200
rect 10232 7148 10284 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 5080 6944 5132 6996
rect 6644 6944 6696 6996
rect 2412 6851 2464 6860
rect 2412 6817 2421 6851
rect 2421 6817 2455 6851
rect 2455 6817 2464 6851
rect 2412 6808 2464 6817
rect 5356 6808 5408 6860
rect 6092 6876 6144 6928
rect 1492 6604 1544 6656
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 5448 6740 5500 6792
rect 5724 6808 5776 6860
rect 6184 6808 6236 6860
rect 8208 6808 8260 6860
rect 9956 6876 10008 6928
rect 11980 6808 12032 6860
rect 12624 6808 12676 6860
rect 2688 6672 2740 6724
rect 7932 6672 7984 6724
rect 2504 6604 2556 6656
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 8392 6604 8444 6656
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 13452 6647 13504 6656
rect 13452 6613 13461 6647
rect 13461 6613 13495 6647
rect 13495 6613 13504 6647
rect 13452 6604 13504 6613
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 3056 6443 3108 6452
rect 3056 6409 3065 6443
rect 3065 6409 3099 6443
rect 3099 6409 3108 6443
rect 3056 6400 3108 6409
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 6828 6400 6880 6452
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 11980 6400 12032 6452
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 9680 6332 9732 6384
rect 5172 6264 5224 6316
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 8668 6264 8720 6316
rect 9588 6264 9640 6316
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 7104 6196 7156 6248
rect 8116 6196 8168 6248
rect 9312 6196 9364 6248
rect 9772 6196 9824 6248
rect 1860 6128 1912 6180
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 8852 6128 8904 6180
rect 10048 6196 10100 6248
rect 10140 6128 10192 6180
rect 5264 6060 5316 6112
rect 5816 6103 5868 6112
rect 5816 6069 5825 6103
rect 5825 6069 5859 6103
rect 5859 6069 5868 6103
rect 5816 6060 5868 6069
rect 7656 6060 7708 6112
rect 8116 6103 8168 6112
rect 8116 6069 8125 6103
rect 8125 6069 8159 6103
rect 8159 6069 8168 6103
rect 8116 6060 8168 6069
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 1676 5856 1728 5908
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 4896 5856 4948 5908
rect 5264 5856 5316 5908
rect 6184 5856 6236 5908
rect 6736 5856 6788 5908
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 8300 5856 8352 5908
rect 8852 5856 8904 5908
rect 9588 5856 9640 5908
rect 10416 5856 10468 5908
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 2596 5788 2648 5840
rect 2688 5720 2740 5772
rect 2780 5720 2832 5772
rect 5080 5788 5132 5840
rect 5816 5788 5868 5840
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 3148 5652 3200 5704
rect 2964 5584 3016 5636
rect 4160 5652 4212 5704
rect 4804 5720 4856 5772
rect 6276 5788 6328 5840
rect 11980 5856 12032 5908
rect 13452 5788 13504 5840
rect 6644 5720 6696 5772
rect 8208 5720 8260 5772
rect 8576 5720 8628 5772
rect 10508 5720 10560 5772
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 11888 5763 11940 5772
rect 11888 5729 11922 5763
rect 11922 5729 11940 5763
rect 11888 5720 11940 5729
rect 4896 5652 4948 5704
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 4804 5584 4856 5636
rect 1308 5516 1360 5568
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 3148 5516 3200 5568
rect 6644 5516 6696 5568
rect 8300 5516 8352 5568
rect 8668 5516 8720 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 4712 5312 4764 5364
rect 5908 5312 5960 5364
rect 2688 5244 2740 5296
rect 2596 5176 2648 5228
rect 6552 5176 6604 5228
rect 7380 5176 7432 5228
rect 2320 5108 2372 5160
rect 5908 5108 5960 5160
rect 7748 5312 7800 5364
rect 7748 5176 7800 5228
rect 9312 5176 9364 5228
rect 10416 5312 10468 5364
rect 11612 5355 11664 5364
rect 11612 5321 11621 5355
rect 11621 5321 11655 5355
rect 11655 5321 11664 5355
rect 11612 5312 11664 5321
rect 10324 5176 10376 5228
rect 2964 5040 3016 5092
rect 3608 5040 3660 5092
rect 4160 5040 4212 5092
rect 6276 5040 6328 5092
rect 8208 5108 8260 5160
rect 940 4972 992 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 5448 4972 5500 5024
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 6920 4972 6972 5024
rect 7748 4972 7800 5024
rect 8576 5040 8628 5092
rect 10600 5176 10652 5228
rect 11336 5176 11388 5228
rect 11888 5176 11940 5228
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 9496 5015 9548 5024
rect 9496 4981 9505 5015
rect 9505 4981 9539 5015
rect 9539 4981 9548 5015
rect 9496 4972 9548 4981
rect 10876 4972 10928 5024
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 4436 4768 4488 4820
rect 4988 4768 5040 4820
rect 5540 4768 5592 4820
rect 6644 4811 6696 4820
rect 6644 4777 6653 4811
rect 6653 4777 6687 4811
rect 6687 4777 6696 4811
rect 6644 4768 6696 4777
rect 7840 4768 7892 4820
rect 8944 4768 8996 4820
rect 9588 4768 9640 4820
rect 10508 4768 10560 4820
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 12624 4768 12676 4820
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 3148 4700 3200 4752
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 2596 4496 2648 4548
rect 3608 4700 3660 4752
rect 3976 4700 4028 4752
rect 8300 4700 8352 4752
rect 11336 4700 11388 4752
rect 4896 4632 4948 4684
rect 6828 4632 6880 4684
rect 7380 4632 7432 4684
rect 4712 4496 4764 4548
rect 5356 4564 5408 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 9680 4632 9732 4684
rect 10048 4632 10100 4684
rect 12440 4632 12492 4684
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 6644 4496 6696 4548
rect 11244 4496 11296 4548
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 2780 4428 2832 4480
rect 6828 4428 6880 4480
rect 7380 4428 7432 4480
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 12808 4428 12860 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 2964 4224 3016 4276
rect 4988 4224 5040 4276
rect 5356 4224 5408 4276
rect 6736 4224 6788 4276
rect 6828 4267 6880 4276
rect 6828 4233 6837 4267
rect 6837 4233 6871 4267
rect 6871 4233 6880 4267
rect 6828 4224 6880 4233
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 5448 4088 5500 4140
rect 7380 4156 7432 4208
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 8024 4088 8076 4140
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 8944 4088 8996 4140
rect 9496 4088 9548 4140
rect 9772 4088 9824 4140
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 5724 4020 5776 4072
rect 6828 4020 6880 4072
rect 6920 4020 6972 4072
rect 10600 4020 10652 4072
rect 11520 4156 11572 4208
rect 10968 4088 11020 4140
rect 11336 4088 11388 4140
rect 11060 4020 11112 4072
rect 12348 4156 12400 4208
rect 12532 4156 12584 4208
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 3608 3952 3660 4004
rect 4988 3952 5040 4004
rect 1400 3884 1452 3936
rect 4896 3884 4948 3936
rect 6000 3952 6052 4004
rect 7380 3952 7432 4004
rect 8208 3952 8260 4004
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7932 3884 7984 3936
rect 8300 3884 8352 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 12532 3884 12584 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 2688 3680 2740 3732
rect 2964 3680 3016 3732
rect 3608 3680 3660 3732
rect 4712 3723 4764 3732
rect 4712 3689 4721 3723
rect 4721 3689 4755 3723
rect 4755 3689 4764 3723
rect 4712 3680 4764 3689
rect 4804 3680 4856 3732
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 5632 3680 5684 3732
rect 6000 3680 6052 3732
rect 6184 3680 6236 3732
rect 7472 3723 7524 3732
rect 7472 3689 7481 3723
rect 7481 3689 7515 3723
rect 7515 3689 7524 3723
rect 7472 3680 7524 3689
rect 7840 3680 7892 3732
rect 8484 3680 8536 3732
rect 9588 3680 9640 3732
rect 12348 3723 12400 3732
rect 12348 3689 12357 3723
rect 12357 3689 12391 3723
rect 12391 3689 12400 3723
rect 12348 3680 12400 3689
rect 12992 3723 13044 3732
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 4252 3612 4304 3664
rect 5908 3612 5960 3664
rect 11336 3612 11388 3664
rect 2320 3587 2372 3596
rect 2320 3553 2329 3587
rect 2329 3553 2363 3587
rect 2363 3553 2372 3587
rect 2320 3544 2372 3553
rect 2964 3544 3016 3596
rect 3424 3544 3476 3596
rect 4896 3544 4948 3596
rect 7932 3544 7984 3596
rect 8760 3544 8812 3596
rect 10692 3544 10744 3596
rect 10876 3544 10928 3596
rect 4160 3476 4212 3528
rect 5356 3476 5408 3528
rect 8944 3476 8996 3528
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 2596 3408 2648 3460
rect 7196 3408 7248 3460
rect 12440 3408 12492 3460
rect 3056 3383 3108 3392
rect 3056 3349 3065 3383
rect 3065 3349 3099 3383
rect 3099 3349 3108 3383
rect 3056 3340 3108 3349
rect 5448 3340 5500 3392
rect 7748 3340 7800 3392
rect 8852 3340 8904 3392
rect 9680 3340 9732 3392
rect 11336 3340 11388 3392
rect 12992 3340 13044 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 2044 3136 2096 3188
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3516 3136 3568 3188
rect 4252 3136 4304 3188
rect 5540 3136 5592 3188
rect 5908 3136 5960 3188
rect 6920 3136 6972 3188
rect 8300 3136 8352 3188
rect 8484 3136 8536 3188
rect 7288 3068 7340 3120
rect 10692 3179 10744 3188
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 11152 3136 11204 3188
rect 4160 3000 4212 3052
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 2044 2975 2096 2984
rect 2044 2941 2053 2975
rect 2053 2941 2087 2975
rect 2087 2941 2096 2975
rect 2044 2932 2096 2941
rect 3516 2932 3568 2984
rect 7472 2975 7524 2984
rect 7472 2941 7481 2975
rect 7481 2941 7515 2975
rect 7515 2941 7524 2975
rect 7472 2932 7524 2941
rect 4712 2864 4764 2916
rect 7288 2864 7340 2916
rect 204 2796 256 2848
rect 1308 2796 1360 2848
rect 2136 2796 2188 2848
rect 3516 2796 3568 2848
rect 8944 2975 8996 2984
rect 8944 2941 8978 2975
rect 8978 2941 8996 2975
rect 8944 2932 8996 2941
rect 12072 3136 12124 3188
rect 12624 3136 12676 3188
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 13268 3000 13320 3052
rect 8852 2864 8904 2916
rect 9588 2796 9640 2848
rect 11152 2796 11204 2848
rect 12072 2796 12124 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 12900 2796 12952 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 2412 2456 2464 2508
rect 4344 2592 4396 2644
rect 5264 2592 5316 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 6736 2635 6788 2644
rect 5632 2592 5684 2601
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 10876 2592 10928 2644
rect 12440 2592 12492 2644
rect 13452 2592 13504 2644
rect 7104 2524 7156 2576
rect 11060 2524 11112 2576
rect 4252 2456 4304 2508
rect 7012 2456 7064 2508
rect 9588 2499 9640 2508
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 10876 2456 10928 2508
rect 12716 2524 12768 2576
rect 5448 2388 5500 2440
rect 8484 2388 8536 2440
rect 2780 2363 2832 2372
rect 2780 2329 2789 2363
rect 2789 2329 2823 2363
rect 2823 2329 2832 2363
rect 2780 2320 2832 2329
rect 2964 2320 3016 2372
rect 8944 2388 8996 2440
rect 13268 2431 13320 2440
rect 2412 2295 2464 2304
rect 2412 2261 2421 2295
rect 2421 2261 2455 2295
rect 2455 2261 2464 2295
rect 2412 2252 2464 2261
rect 3332 2252 3384 2304
rect 5264 2295 5316 2304
rect 5264 2261 5273 2295
rect 5273 2261 5307 2295
rect 5307 2261 5316 2295
rect 5264 2252 5316 2261
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14096 2252 14148 2304
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 10600 2048 10652 2100
rect 12532 2048 12584 2100
rect 5816 552 5868 604
rect 6184 552 6236 604
rect 9772 552 9824 604
rect 9956 552 10008 604
rect 10232 552 10284 604
rect 12164 552 12216 604
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39520 10194 40000
rect 10598 39520 10654 40000
rect 10966 39520 11022 40000
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39522 13414 40000
rect 13188 39520 13414 39522
rect 13726 39520 13782 40000
rect 14186 39522 14242 40000
rect 13832 39520 14242 39522
rect 14554 39520 14610 40000
rect 14922 39522 14978 40000
rect 14922 39520 15056 39522
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34746 244 39520
rect 204 34740 256 34746
rect 204 34682 256 34688
rect 584 33969 612 39520
rect 952 35290 980 39520
rect 940 35284 992 35290
rect 940 35226 992 35232
rect 1412 34202 1440 39520
rect 1582 38720 1638 38729
rect 1582 38655 1638 38664
rect 1490 36408 1546 36417
rect 1490 36343 1546 36352
rect 1400 34196 1452 34202
rect 1400 34138 1452 34144
rect 570 33960 626 33969
rect 570 33895 626 33904
rect 1504 33658 1532 36343
rect 1596 35834 1624 38655
rect 1584 35828 1636 35834
rect 1584 35770 1636 35776
rect 1780 35193 1808 39520
rect 1860 35488 1912 35494
rect 1860 35430 1912 35436
rect 1766 35184 1822 35193
rect 1676 35148 1728 35154
rect 1766 35119 1822 35128
rect 1676 35090 1728 35096
rect 1688 34134 1716 35090
rect 1676 34128 1728 34134
rect 1582 34096 1638 34105
rect 1676 34070 1728 34076
rect 1582 34031 1638 34040
rect 1492 33652 1544 33658
rect 1492 33594 1544 33600
rect 1596 33114 1624 34031
rect 1688 33130 1716 34070
rect 1584 33108 1636 33114
rect 1688 33102 1808 33130
rect 1584 33050 1636 33056
rect 1676 32972 1728 32978
rect 1676 32914 1728 32920
rect 1688 32502 1716 32914
rect 1676 32496 1728 32502
rect 1674 32464 1676 32473
rect 1728 32464 1730 32473
rect 1674 32399 1730 32408
rect 1582 31648 1638 31657
rect 1582 31583 1638 31592
rect 1596 29850 1624 31583
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1582 29336 1638 29345
rect 1582 29271 1584 29280
rect 1636 29271 1638 29280
rect 1584 29242 1636 29248
rect 1780 29073 1808 33102
rect 1766 29064 1822 29073
rect 1766 28999 1822 29008
rect 1582 27024 1638 27033
rect 1582 26959 1638 26968
rect 1596 26042 1624 26959
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1872 25945 1900 35430
rect 2148 35290 2176 39520
rect 2608 35329 2636 39520
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2594 35320 2650 35329
rect 2136 35284 2188 35290
rect 2594 35255 2650 35264
rect 2136 35226 2188 35232
rect 2504 35148 2556 35154
rect 2504 35090 2556 35096
rect 2516 34542 2544 35090
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 2136 34536 2188 34542
rect 2136 34478 2188 34484
rect 2504 34536 2556 34542
rect 2504 34478 2556 34484
rect 1952 34060 2004 34066
rect 1952 34002 2004 34008
rect 1964 33454 1992 34002
rect 1952 33448 2004 33454
rect 1950 33416 1952 33425
rect 2004 33416 2006 33425
rect 1950 33351 2006 33360
rect 2056 27606 2084 34478
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 1858 25936 1914 25945
rect 1858 25871 1914 25880
rect 1952 25696 2004 25702
rect 1952 25638 2004 25644
rect 1964 25498 1992 25638
rect 1952 25492 2004 25498
rect 1952 25434 2004 25440
rect 1582 24576 1638 24585
rect 1582 24511 1638 24520
rect 1596 23322 1624 24511
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1688 22710 1716 23122
rect 1676 22704 1728 22710
rect 1674 22672 1676 22681
rect 1728 22672 1730 22681
rect 1674 22607 1730 22616
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 1582 21992 1638 22001
rect 1582 21927 1584 21936
rect 1636 21927 1638 21936
rect 1584 21898 1636 21904
rect 1688 20942 1716 22034
rect 1676 20936 1728 20942
rect 1674 20904 1676 20913
rect 1728 20904 1730 20913
rect 1674 20839 1730 20848
rect 1582 19952 1638 19961
rect 1582 19887 1638 19896
rect 1596 18426 1624 19887
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1950 18320 2006 18329
rect 1950 18255 1952 18264
rect 2004 18255 2006 18264
rect 1952 18226 2004 18232
rect 1582 17640 1638 17649
rect 1582 17575 1638 17584
rect 1596 16250 1624 17575
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1950 16144 2006 16153
rect 1950 16079 1952 16088
rect 2004 16079 2006 16088
rect 1952 16050 2004 16056
rect 1582 15192 1638 15201
rect 1582 15127 1638 15136
rect 1596 13530 1624 15127
rect 2148 14929 2176 34478
rect 2318 33552 2374 33561
rect 2318 33487 2320 33496
rect 2372 33487 2374 33496
rect 2320 33458 2372 33464
rect 2412 31204 2464 31210
rect 2412 31146 2464 31152
rect 2424 30938 2452 31146
rect 2792 30938 2820 35566
rect 2976 34202 3004 39520
rect 3344 35834 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4016 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3988 35834 4016 37182
rect 3332 35828 3384 35834
rect 3332 35770 3384 35776
rect 3976 35828 4028 35834
rect 3976 35770 4028 35776
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 3516 34468 3568 34474
rect 3516 34410 3568 34416
rect 2964 34196 3016 34202
rect 2964 34138 3016 34144
rect 3148 34060 3200 34066
rect 3148 34002 3200 34008
rect 3160 33318 3188 34002
rect 3528 33862 3556 34410
rect 3516 33856 3568 33862
rect 3516 33798 3568 33804
rect 3148 33312 3200 33318
rect 3148 33254 3200 33260
rect 3424 33312 3476 33318
rect 3424 33254 3476 33260
rect 3056 31680 3108 31686
rect 3056 31622 3108 31628
rect 3068 31142 3096 31622
rect 2964 31136 3016 31142
rect 2964 31078 3016 31084
rect 3056 31136 3108 31142
rect 3056 31078 3108 31084
rect 2412 30932 2464 30938
rect 2412 30874 2464 30880
rect 2780 30932 2832 30938
rect 2780 30874 2832 30880
rect 2228 30864 2280 30870
rect 2228 30806 2280 30812
rect 2240 30394 2268 30806
rect 2792 30682 2820 30874
rect 2700 30654 2820 30682
rect 2872 30728 2924 30734
rect 2872 30670 2924 30676
rect 2228 30388 2280 30394
rect 2228 30330 2280 30336
rect 2700 30274 2728 30654
rect 2884 30546 2912 30670
rect 2516 30246 2728 30274
rect 2792 30518 2912 30546
rect 2516 30054 2544 30246
rect 2504 30048 2556 30054
rect 2504 29990 2556 29996
rect 2516 29753 2544 29990
rect 2502 29744 2558 29753
rect 2320 29708 2372 29714
rect 2502 29679 2558 29688
rect 2320 29650 2372 29656
rect 2332 29238 2360 29650
rect 2792 29510 2820 30518
rect 2976 30258 3004 31078
rect 2964 30252 3016 30258
rect 2964 30194 3016 30200
rect 2872 30048 2924 30054
rect 2872 29990 2924 29996
rect 2780 29504 2832 29510
rect 2780 29446 2832 29452
rect 2320 29232 2372 29238
rect 2320 29174 2372 29180
rect 2792 28762 2820 29446
rect 2884 29306 2912 29990
rect 2976 29850 3004 30194
rect 2964 29844 3016 29850
rect 2964 29786 3016 29792
rect 2872 29300 2924 29306
rect 2872 29242 2924 29248
rect 2870 29064 2926 29073
rect 2870 28999 2926 29008
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2884 28218 2912 28999
rect 3068 28218 3096 31078
rect 3160 30705 3188 33254
rect 3146 30696 3202 30705
rect 3146 30631 3202 30640
rect 3240 30660 3292 30666
rect 2872 28212 2924 28218
rect 2872 28154 2924 28160
rect 3056 28212 3108 28218
rect 3056 28154 3108 28160
rect 2884 28014 2912 28154
rect 2962 28112 3018 28121
rect 2962 28047 3018 28056
rect 2872 28008 2924 28014
rect 2872 27950 2924 27956
rect 2412 27940 2464 27946
rect 2412 27882 2464 27888
rect 2424 27674 2452 27882
rect 2412 27668 2464 27674
rect 2412 27610 2464 27616
rect 2976 27606 3004 28047
rect 2504 27600 2556 27606
rect 2504 27542 2556 27548
rect 2964 27600 3016 27606
rect 2964 27542 3016 27548
rect 2228 27532 2280 27538
rect 2228 27474 2280 27480
rect 2240 27062 2268 27474
rect 2516 27062 2544 27542
rect 2780 27532 2832 27538
rect 2780 27474 2832 27480
rect 2792 27441 2820 27474
rect 2778 27432 2834 27441
rect 2778 27367 2834 27376
rect 2228 27056 2280 27062
rect 2228 26998 2280 27004
rect 2504 27056 2556 27062
rect 2504 26998 2556 27004
rect 2688 26920 2740 26926
rect 2688 26862 2740 26868
rect 2700 26586 2728 26862
rect 2964 26852 3016 26858
rect 2964 26794 3016 26800
rect 2976 26586 3004 26794
rect 2228 26580 2280 26586
rect 2228 26522 2280 26528
rect 2688 26580 2740 26586
rect 2688 26522 2740 26528
rect 2964 26580 3016 26586
rect 2964 26522 3016 26528
rect 2240 24750 2268 26522
rect 2780 25424 2832 25430
rect 2780 25366 2832 25372
rect 2688 25288 2740 25294
rect 2688 25230 2740 25236
rect 2596 25220 2648 25226
rect 2596 25162 2648 25168
rect 2412 25152 2464 25158
rect 2412 25094 2464 25100
rect 2424 24750 2452 25094
rect 2228 24744 2280 24750
rect 2228 24686 2280 24692
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2424 22778 2452 24686
rect 2608 24614 2636 25162
rect 2700 24682 2728 25230
rect 2688 24676 2740 24682
rect 2688 24618 2740 24624
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2608 24410 2636 24550
rect 2596 24404 2648 24410
rect 2596 24346 2648 24352
rect 2700 22778 2728 24618
rect 2792 24410 2820 25366
rect 2976 25294 3004 26522
rect 2964 25288 3016 25294
rect 2964 25230 3016 25236
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 3160 23066 3188 30631
rect 3240 30602 3292 30608
rect 3252 30190 3280 30602
rect 3436 30258 3464 33254
rect 3528 31346 3556 33798
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 4080 33454 4108 34478
rect 4172 34202 4200 39520
rect 4540 35737 4568 39520
rect 4526 35728 4582 35737
rect 4436 35692 4488 35698
rect 4526 35663 4582 35672
rect 4436 35634 4488 35640
rect 4160 34196 4212 34202
rect 4160 34138 4212 34144
rect 4160 34060 4212 34066
rect 4160 34002 4212 34008
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 4172 33318 4200 34002
rect 4250 33960 4306 33969
rect 4250 33895 4252 33904
rect 4304 33895 4306 33904
rect 4252 33866 4304 33872
rect 4252 33448 4304 33454
rect 4252 33390 4304 33396
rect 4160 33312 4212 33318
rect 4160 33254 4212 33260
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 4172 32298 4200 33254
rect 4264 33114 4292 33390
rect 4252 33108 4304 33114
rect 4252 33050 4304 33056
rect 4160 32292 4212 32298
rect 4160 32234 4212 32240
rect 4264 31958 4292 33050
rect 4252 31952 4304 31958
rect 4252 31894 4304 31900
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 4080 31482 4108 31826
rect 4448 31668 4476 35634
rect 4620 35488 4672 35494
rect 4620 35430 4672 35436
rect 4264 31640 4476 31668
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 3516 31340 3568 31346
rect 3516 31282 3568 31288
rect 4160 31204 4212 31210
rect 4080 31164 4160 31192
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3424 30252 3476 30258
rect 3424 30194 3476 30200
rect 3240 30184 3292 30190
rect 3240 30126 3292 30132
rect 3436 29714 3464 30194
rect 3424 29708 3476 29714
rect 3424 29650 3476 29656
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 4080 29170 4108 31164
rect 4160 31146 4212 31152
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 3516 28688 3568 28694
rect 3516 28630 3568 28636
rect 3528 28082 3556 28630
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 4080 27062 4108 27406
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 4264 25820 4292 31640
rect 4632 31482 4660 35430
rect 4710 35320 4766 35329
rect 5000 35290 5028 39520
rect 5368 36922 5396 39520
rect 5356 36916 5408 36922
rect 5356 36858 5408 36864
rect 5448 36236 5500 36242
rect 5448 36178 5500 36184
rect 5460 35698 5488 36178
rect 5736 35766 5764 39520
rect 5908 36576 5960 36582
rect 5908 36518 5960 36524
rect 5724 35760 5776 35766
rect 5724 35702 5776 35708
rect 5448 35692 5500 35698
rect 5448 35634 5500 35640
rect 4710 35255 4712 35264
rect 4764 35255 4766 35264
rect 4988 35284 5040 35290
rect 4712 35226 4764 35232
rect 4988 35226 5040 35232
rect 4712 35148 4764 35154
rect 4712 35090 4764 35096
rect 5632 35148 5684 35154
rect 5632 35090 5684 35096
rect 4724 33862 4752 35090
rect 5644 34678 5672 35090
rect 5632 34672 5684 34678
rect 5632 34614 5684 34620
rect 4804 34400 4856 34406
rect 4804 34342 4856 34348
rect 4712 33856 4764 33862
rect 4712 33798 4764 33804
rect 4620 31476 4672 31482
rect 4620 31418 4672 31424
rect 4620 31340 4672 31346
rect 4620 31282 4672 31288
rect 4436 31136 4488 31142
rect 4356 31084 4436 31090
rect 4356 31078 4488 31084
rect 4356 31062 4476 31078
rect 4356 30802 4384 31062
rect 4344 30796 4396 30802
rect 4344 30738 4396 30744
rect 4356 29850 4384 30738
rect 4632 30734 4660 31282
rect 4528 30728 4580 30734
rect 4528 30670 4580 30676
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4540 30054 4568 30670
rect 4632 30394 4660 30670
rect 4620 30388 4672 30394
rect 4620 30330 4672 30336
rect 4528 30048 4580 30054
rect 4528 29990 4580 29996
rect 4344 29844 4396 29850
rect 4344 29786 4396 29792
rect 4540 28762 4568 29990
rect 4528 28756 4580 28762
rect 4528 28698 4580 28704
rect 4344 27532 4396 27538
rect 4344 27474 4396 27480
rect 4356 27130 4384 27474
rect 4344 27124 4396 27130
rect 4344 27066 4396 27072
rect 4344 25832 4396 25838
rect 4264 25792 4344 25820
rect 4344 25774 4396 25780
rect 4356 25702 4384 25774
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 4344 25696 4396 25702
rect 4344 25638 4396 25644
rect 4528 25696 4580 25702
rect 4528 25638 4580 25644
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 4080 24954 4108 25638
rect 4252 25492 4304 25498
rect 4252 25434 4304 25440
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 4172 23866 4200 24142
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4172 23066 4200 23802
rect 3068 23038 3188 23066
rect 4080 23038 4200 23066
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2778 22536 2834 22545
rect 2778 22471 2834 22480
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2424 22234 2452 22374
rect 2792 22250 2820 22471
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 2700 22222 3004 22250
rect 3068 22234 3096 23038
rect 3148 22976 3200 22982
rect 3148 22918 3200 22924
rect 3160 22642 3188 22918
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 4080 22642 4108 23038
rect 4264 22964 4292 25434
rect 4172 22936 4292 22964
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 2516 21622 2544 22170
rect 2700 21690 2728 22222
rect 2976 22166 3004 22222
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2504 21616 2556 21622
rect 2504 21558 2556 21564
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 2700 21146 2728 21422
rect 3068 21418 3096 21966
rect 3056 21412 3108 21418
rect 3056 21354 3108 21360
rect 3068 21146 3096 21354
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2134 14920 2190 14929
rect 2134 14855 2190 14864
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1768 13456 1820 13462
rect 1768 13398 1820 13404
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 12481 1716 13330
rect 1780 12986 1808 13398
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 2332 12782 2360 13806
rect 2700 13530 2728 14758
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 1674 12472 1730 12481
rect 1674 12407 1676 12416
rect 1728 12407 1730 12416
rect 1676 12378 1728 12384
rect 2332 11762 2360 12718
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2516 12170 2544 12650
rect 2608 12442 2636 13262
rect 2792 12889 2820 15846
rect 3436 14362 3464 22170
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 4080 21690 4108 22578
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3528 17134 3556 18022
rect 3896 17610 3924 18090
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3884 17604 3936 17610
rect 3884 17546 3936 17552
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3988 16046 4016 17478
rect 4080 16114 4108 18022
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3884 15904 3936 15910
rect 4068 15904 4120 15910
rect 3936 15864 4016 15892
rect 3884 15846 3936 15852
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3160 14334 3464 14362
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2778 12880 2834 12889
rect 2778 12815 2834 12824
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 2056 11014 2084 11562
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 1872 10606 1900 10950
rect 1860 10600 1912 10606
rect 1582 10568 1638 10577
rect 1860 10542 1912 10548
rect 1582 10503 1638 10512
rect 1596 9654 1624 10503
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1780 9518 1808 10406
rect 2056 9586 2084 10950
rect 2884 10674 2912 12582
rect 3068 12102 3096 13330
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3068 11354 3096 12038
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10266 2452 10406
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1780 8634 1808 9454
rect 2056 8634 2084 9522
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 1584 7200 1636 7206
rect 1952 7200 2004 7206
rect 1584 7142 1636 7148
rect 1950 7168 1952 7177
rect 2004 7168 2006 7177
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1308 5568 1360 5574
rect 1308 5510 1360 5516
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 570 4312 626 4321
rect 570 4247 626 4256
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 480 244 2790
rect 584 480 612 4247
rect 952 480 980 4966
rect 1320 2854 1348 5510
rect 1400 4616 1452 4622
rect 1398 4584 1400 4593
rect 1452 4584 1454 4593
rect 1398 4519 1454 4528
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 1412 480 1440 3878
rect 1504 3505 1532 6598
rect 1596 5817 1624 7142
rect 1950 7103 2006 7112
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1688 5914 1716 6190
rect 1872 6186 1900 6598
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1582 5808 1638 5817
rect 1582 5743 1638 5752
rect 1766 4720 1822 4729
rect 1766 4655 1822 4664
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1780 480 1808 4655
rect 1872 1193 1900 6122
rect 2056 3194 2084 7414
rect 2332 5370 2360 9454
rect 2424 9178 2452 9998
rect 2780 9988 2832 9994
rect 2700 9948 2780 9976
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2700 9042 2728 9948
rect 2780 9930 2832 9936
rect 2884 9722 2912 10134
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2884 9110 2912 9658
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8634 2820 8978
rect 3068 8974 3096 9522
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2884 8634 2912 8910
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2792 8537 2820 8570
rect 2778 8528 2834 8537
rect 2778 8463 2834 8472
rect 2778 8120 2834 8129
rect 2884 8090 2912 8570
rect 2778 8055 2834 8064
rect 2872 8084 2924 8090
rect 2792 6882 2820 8055
rect 2872 8026 2924 8032
rect 3054 7304 3110 7313
rect 3054 7239 3110 7248
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2700 6854 2820 6882
rect 2870 6896 2926 6905
rect 2424 5914 2452 6802
rect 2700 6730 2728 6854
rect 2870 6831 2926 6840
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2332 5166 2360 5306
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2424 4826 2452 5850
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4185 2360 4422
rect 2318 4176 2374 4185
rect 2318 4111 2374 4120
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2332 3505 2360 3538
rect 2318 3496 2374 3505
rect 2318 3431 2374 3440
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2136 2848 2188 2854
rect 1950 2816 2006 2825
rect 2136 2790 2188 2796
rect 1950 2751 2006 2760
rect 1964 2650 1992 2751
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 1858 1184 1914 1193
rect 1858 1119 1914 1128
rect 2148 480 2176 2790
rect 2516 2553 2544 6598
rect 2884 5930 2912 6831
rect 3068 6458 3096 7239
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 2700 5902 2912 5930
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2608 5234 2636 5782
rect 2700 5778 2728 5902
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2700 5302 2728 5714
rect 2792 5370 2820 5714
rect 3160 5710 3188 14334
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3344 13802 3372 14214
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3344 12646 3372 13738
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3528 11898 3556 12106
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10674 3464 10950
rect 3528 10810 3556 11834
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3436 9722 3464 10610
rect 3528 10062 3556 10746
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 3712 10266 3740 10474
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3424 9512 3476 9518
rect 3330 9480 3386 9489
rect 3424 9454 3476 9460
rect 3330 9415 3332 9424
rect 3384 9415 3386 9424
rect 3332 9386 3384 9392
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2608 4554 2636 5170
rect 2976 5098 3004 5578
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2608 4146 2636 4490
rect 2792 4486 2820 4762
rect 2976 4622 3004 5034
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2688 3732 2740 3738
rect 2792 3720 2820 4422
rect 2976 4282 3004 4558
rect 3068 4321 3096 5510
rect 3160 4758 3188 5510
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3054 4312 3110 4321
rect 2964 4276 3016 4282
rect 3054 4247 3110 4256
rect 2964 4218 3016 4224
rect 2976 3738 3004 4218
rect 2740 3692 2820 3720
rect 2964 3732 3016 3738
rect 2688 3674 2740 3680
rect 2964 3674 3016 3680
rect 3436 3602 3464 9454
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 8838 3556 9318
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3790 8392 3846 8401
rect 3790 8327 3846 8336
rect 3804 8294 3832 8327
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3988 6066 4016 15864
rect 4068 15846 4120 15852
rect 4080 15706 4108 15846
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4080 15094 4108 15370
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 7886 4108 8298
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4080 6905 4108 7822
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 3528 6038 4016 6066
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2502 2544 2558 2553
rect 2412 2508 2464 2514
rect 2502 2479 2558 2488
rect 2412 2450 2464 2456
rect 2424 2310 2452 2450
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2424 1737 2452 2246
rect 2410 1728 2466 1737
rect 2410 1663 2466 1672
rect 2608 480 2636 3402
rect 2976 3194 3004 3538
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 3068 3097 3096 3334
rect 3528 3194 3556 6038
rect 4172 5794 4200 22936
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4264 21690 4292 21830
rect 4252 21684 4304 21690
rect 4252 21626 4304 21632
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4264 16454 4292 17002
rect 4356 16658 4384 25638
rect 4540 24410 4568 25638
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 4528 24404 4580 24410
rect 4528 24346 4580 24352
rect 4540 23866 4568 24346
rect 4528 23860 4580 23866
rect 4528 23802 4580 23808
rect 4436 23248 4488 23254
rect 4436 23190 4488 23196
rect 4448 22778 4476 23190
rect 4528 23180 4580 23186
rect 4528 23122 4580 23128
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4540 21690 4568 23122
rect 4632 23118 4660 24822
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4632 22778 4660 23054
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4632 22098 4660 22714
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4632 16454 4660 16934
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4264 15910 4292 16390
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4264 15162 4292 15438
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4448 14890 4476 15506
rect 4632 15502 4660 16390
rect 4724 16017 4752 33798
rect 4816 33386 4844 34342
rect 4988 34060 5040 34066
rect 4988 34002 5040 34008
rect 4804 33380 4856 33386
rect 4804 33322 4856 33328
rect 5000 32774 5028 34002
rect 4988 32768 5040 32774
rect 4988 32710 5040 32716
rect 5540 32768 5592 32774
rect 5540 32710 5592 32716
rect 5000 31482 5028 32710
rect 5080 31884 5132 31890
rect 5080 31826 5132 31832
rect 4896 31476 4948 31482
rect 4896 31418 4948 31424
rect 4988 31476 5040 31482
rect 4988 31418 5040 31424
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4816 29306 4844 29582
rect 4804 29300 4856 29306
rect 4804 29242 4856 29248
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 4816 27946 4844 28562
rect 4804 27940 4856 27946
rect 4804 27882 4856 27888
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4816 24274 4844 24550
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4816 23866 4844 24210
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 4908 21593 4936 31418
rect 4986 31376 5042 31385
rect 5092 31346 5120 31826
rect 5448 31680 5500 31686
rect 5448 31622 5500 31628
rect 5356 31476 5408 31482
rect 5356 31418 5408 31424
rect 4986 31311 5042 31320
rect 5080 31340 5132 31346
rect 5000 31278 5028 31311
rect 5080 31282 5132 31288
rect 4988 31272 5040 31278
rect 4988 31214 5040 31220
rect 5092 30920 5120 31282
rect 5000 30892 5120 30920
rect 5000 30666 5028 30892
rect 4988 30660 5040 30666
rect 4988 30602 5040 30608
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 5000 29714 5028 29990
rect 4988 29708 5040 29714
rect 4988 29650 5040 29656
rect 5184 29170 5212 29990
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 4988 28552 5040 28558
rect 4988 28494 5040 28500
rect 5264 28552 5316 28558
rect 5264 28494 5316 28500
rect 5000 28257 5028 28494
rect 4986 28248 5042 28257
rect 5276 28218 5304 28494
rect 4986 28183 4988 28192
rect 5040 28183 5042 28192
rect 5264 28212 5316 28218
rect 4988 28154 5040 28160
rect 5264 28154 5316 28160
rect 5276 27674 5304 28154
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 5000 25702 5028 26182
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 5000 25498 5028 25638
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 5368 25242 5396 31418
rect 5460 30734 5488 31622
rect 5552 30938 5580 32710
rect 5816 32360 5868 32366
rect 5814 32328 5816 32337
rect 5868 32328 5870 32337
rect 5814 32263 5870 32272
rect 5632 32224 5684 32230
rect 5632 32166 5684 32172
rect 5644 31929 5672 32166
rect 5630 31920 5686 31929
rect 5630 31855 5686 31864
rect 5630 31376 5686 31385
rect 5630 31311 5686 31320
rect 5540 30932 5592 30938
rect 5540 30874 5592 30880
rect 5448 30728 5500 30734
rect 5448 30670 5500 30676
rect 5552 30258 5580 30874
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 5448 29300 5500 29306
rect 5448 29242 5500 29248
rect 5460 28626 5488 29242
rect 5448 28620 5500 28626
rect 5448 28562 5500 28568
rect 5460 27062 5488 28562
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5000 24750 5028 25230
rect 5368 25214 5580 25242
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5078 24848 5134 24857
rect 5078 24783 5080 24792
rect 5132 24783 5134 24792
rect 5080 24754 5132 24760
rect 5460 24750 5488 25094
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 5460 24596 5488 24686
rect 5368 24568 5488 24596
rect 5368 22574 5396 24568
rect 5552 24342 5580 25214
rect 5540 24336 5592 24342
rect 5540 24278 5592 24284
rect 5356 22568 5408 22574
rect 5644 22556 5672 31311
rect 5816 30592 5868 30598
rect 5816 30534 5868 30540
rect 5828 30122 5856 30534
rect 5920 30190 5948 36518
rect 6196 36378 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6184 36372 6236 36378
rect 6184 36314 6236 36320
rect 6656 35834 6684 37726
rect 6644 35828 6696 35834
rect 6644 35770 6696 35776
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6276 33992 6328 33998
rect 6276 33934 6328 33940
rect 6288 33454 6316 33934
rect 6276 33448 6328 33454
rect 6276 33390 6328 33396
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6644 33108 6696 33114
rect 6644 33050 6696 33056
rect 6000 32904 6052 32910
rect 6000 32846 6052 32852
rect 6184 32904 6236 32910
rect 6184 32846 6236 32852
rect 6552 32904 6604 32910
rect 6552 32846 6604 32852
rect 6012 32502 6040 32846
rect 6000 32496 6052 32502
rect 6000 32438 6052 32444
rect 6012 32026 6040 32438
rect 6092 32292 6144 32298
rect 6092 32234 6144 32240
rect 6000 32020 6052 32026
rect 6000 31962 6052 31968
rect 6104 30666 6132 32234
rect 6196 32230 6224 32846
rect 6564 32298 6592 32846
rect 6552 32292 6604 32298
rect 6552 32234 6604 32240
rect 6184 32224 6236 32230
rect 6184 32166 6236 32172
rect 6196 31890 6224 32166
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6656 32026 6684 33050
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6196 30734 6224 30765
rect 6184 30728 6236 30734
rect 6182 30696 6184 30705
rect 6236 30696 6238 30705
rect 6092 30660 6144 30666
rect 6182 30631 6238 30640
rect 6644 30660 6696 30666
rect 6092 30602 6144 30608
rect 6196 30394 6224 30631
rect 6644 30602 6696 30608
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6000 30252 6052 30258
rect 6000 30194 6052 30200
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5816 30116 5868 30122
rect 5816 30058 5868 30064
rect 6012 29714 6040 30194
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6656 29782 6684 30602
rect 6644 29776 6696 29782
rect 6644 29718 6696 29724
rect 6000 29708 6052 29714
rect 6000 29650 6052 29656
rect 5908 28960 5960 28966
rect 5908 28902 5960 28908
rect 5920 28422 5948 28902
rect 6012 28490 6040 29650
rect 6276 29504 6328 29510
rect 6276 29446 6328 29452
rect 6288 29170 6316 29446
rect 6276 29164 6328 29170
rect 6276 29106 6328 29112
rect 6288 29050 6316 29106
rect 6196 29022 6316 29050
rect 6196 28694 6224 29022
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6184 28688 6236 28694
rect 6184 28630 6236 28636
rect 6000 28484 6052 28490
rect 6000 28426 6052 28432
rect 5908 28416 5960 28422
rect 5908 28358 5960 28364
rect 5722 28248 5778 28257
rect 5722 28183 5778 28192
rect 5736 23066 5764 28183
rect 5814 27976 5870 27985
rect 5814 27911 5816 27920
rect 5868 27911 5870 27920
rect 5816 27882 5868 27888
rect 5828 25378 5856 27882
rect 5920 26314 5948 28358
rect 6012 26382 6040 28426
rect 6196 28218 6224 28630
rect 6368 28620 6420 28626
rect 6368 28562 6420 28568
rect 6380 28393 6408 28562
rect 6366 28384 6422 28393
rect 6366 28319 6422 28328
rect 6380 28218 6408 28319
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6368 28212 6420 28218
rect 6368 28154 6420 28160
rect 6748 27985 6776 35430
rect 6932 35018 6960 39520
rect 7392 35834 7420 39520
rect 7760 36417 7788 39520
rect 7746 36408 7802 36417
rect 7746 36343 7802 36352
rect 7380 35828 7432 35834
rect 7380 35770 7432 35776
rect 8220 35714 8248 39520
rect 7944 35686 8248 35714
rect 7564 35284 7616 35290
rect 7564 35226 7616 35232
rect 7576 35193 7604 35226
rect 7562 35184 7618 35193
rect 7196 35148 7248 35154
rect 7562 35119 7618 35128
rect 7196 35090 7248 35096
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 7208 34406 7236 35090
rect 7656 34944 7708 34950
rect 7656 34886 7708 34892
rect 7380 34672 7432 34678
rect 7380 34614 7432 34620
rect 7196 34400 7248 34406
rect 7196 34342 7248 34348
rect 7012 34060 7064 34066
rect 7012 34002 7064 34008
rect 7024 33318 7052 34002
rect 7012 33312 7064 33318
rect 7012 33254 7064 33260
rect 7024 32910 7052 33254
rect 7012 32904 7064 32910
rect 7012 32846 7064 32852
rect 7012 32768 7064 32774
rect 7012 32710 7064 32716
rect 7024 32366 7052 32710
rect 7104 32564 7156 32570
rect 7104 32506 7156 32512
rect 7012 32360 7064 32366
rect 7012 32302 7064 32308
rect 6828 32292 6880 32298
rect 6828 32234 6880 32240
rect 6840 32026 6868 32234
rect 7024 32026 7052 32302
rect 6828 32020 6880 32026
rect 6828 31962 6880 31968
rect 7012 32020 7064 32026
rect 7012 31962 7064 31968
rect 6826 30968 6882 30977
rect 6826 30903 6828 30912
rect 6880 30903 6882 30912
rect 6828 30874 6880 30880
rect 6840 29866 6868 30874
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6932 30258 6960 30534
rect 6920 30252 6972 30258
rect 6920 30194 6972 30200
rect 6840 29850 6960 29866
rect 6840 29844 6972 29850
rect 6840 29838 6920 29844
rect 6734 27976 6790 27985
rect 6734 27911 6790 27920
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6184 27056 6236 27062
rect 6184 26998 6236 27004
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 5908 26308 5960 26314
rect 5908 26250 5960 26256
rect 6012 26194 6040 26318
rect 5920 26166 6040 26194
rect 5920 25702 5948 26166
rect 6196 26042 6224 26998
rect 6840 26874 6868 29838
rect 6920 29786 6972 29792
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 7024 26897 7052 29038
rect 6748 26846 6868 26874
rect 7010 26888 7066 26897
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6748 26246 6776 26846
rect 7010 26823 7066 26832
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6840 26586 6868 26726
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6828 26444 6880 26450
rect 6828 26386 6880 26392
rect 6736 26240 6788 26246
rect 6736 26182 6788 26188
rect 6840 26042 6868 26386
rect 6184 26036 6236 26042
rect 6184 25978 6236 25984
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 5908 25696 5960 25702
rect 5908 25638 5960 25644
rect 5920 25498 5948 25638
rect 5908 25492 5960 25498
rect 5908 25434 5960 25440
rect 6196 25430 6224 25978
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6184 25424 6236 25430
rect 5828 25350 6040 25378
rect 6184 25366 6236 25372
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5828 23186 5856 23462
rect 5816 23180 5868 23186
rect 5816 23122 5868 23128
rect 5736 23038 5856 23066
rect 5724 22976 5776 22982
rect 5724 22918 5776 22924
rect 5736 22681 5764 22918
rect 5722 22672 5778 22681
rect 5722 22607 5778 22616
rect 5644 22528 5764 22556
rect 5356 22510 5408 22516
rect 5368 22166 5396 22510
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 4894 21584 4950 21593
rect 4894 21519 4950 21528
rect 5092 21146 5120 22034
rect 5368 21486 5396 22102
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5538 21448 5594 21457
rect 5368 21350 5396 21422
rect 5538 21383 5594 21392
rect 5552 21350 5580 21383
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5368 20942 5396 21286
rect 5552 21078 5580 21286
rect 5540 21072 5592 21078
rect 5540 21014 5592 21020
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5368 20262 5396 20878
rect 5644 20602 5672 20946
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5264 18828 5316 18834
rect 5368 18816 5396 20198
rect 5316 18788 5396 18816
rect 5264 18770 5316 18776
rect 5368 18290 5396 18788
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5460 18154 5488 18770
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5538 17776 5594 17785
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4896 17740 4948 17746
rect 5736 17746 5764 22528
rect 5538 17711 5594 17720
rect 5724 17740 5776 17746
rect 4896 17682 4948 17688
rect 4816 17338 4844 17682
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4908 16794 4936 17682
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5000 16998 5028 17614
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5552 16726 5580 17711
rect 5724 17682 5776 17688
rect 5828 17218 5856 23038
rect 5908 22500 5960 22506
rect 5908 22442 5960 22448
rect 5920 22234 5948 22442
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5920 21690 5948 22170
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5920 21049 5948 21286
rect 5906 21040 5962 21049
rect 5906 20975 5962 20984
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5920 17678 5948 18226
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5736 17190 5856 17218
rect 5920 17202 5948 17614
rect 5908 17196 5960 17202
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 4710 16008 4766 16017
rect 5552 15978 5580 16662
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 4710 15943 4766 15952
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5644 15910 5672 16594
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4618 14920 4674 14929
rect 4436 14884 4488 14890
rect 4618 14855 4620 14864
rect 4436 14826 4488 14832
rect 4672 14855 4674 14864
rect 4620 14826 4672 14832
rect 4448 14618 4476 14826
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4264 11898 4292 13398
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4356 11830 4384 12922
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4264 9518 4292 9998
rect 4448 9994 4476 10406
rect 4436 9988 4488 9994
rect 4488 9948 4568 9976
rect 4436 9930 4488 9936
rect 4540 9722 4568 9948
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8430 4384 8978
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4448 8242 4476 9386
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4540 8294 4568 9046
rect 4356 8214 4476 8242
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4172 5766 4292 5794
rect 4160 5704 4212 5710
rect 3988 5652 4160 5658
rect 3988 5646 4212 5652
rect 3988 5630 4200 5646
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3620 4758 3648 5034
rect 3988 4758 4016 5630
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3620 3777 3648 3946
rect 3606 3768 3662 3777
rect 3606 3703 3608 3712
rect 3660 3703 3662 3712
rect 3608 3674 3660 3680
rect 4172 3534 4200 5034
rect 4264 3670 4292 5766
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3054 3088 3110 3097
rect 3054 3023 3110 3032
rect 3528 2990 3556 3130
rect 4172 3058 4200 3470
rect 4264 3194 4292 3606
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 2778 2408 2834 2417
rect 2778 2343 2780 2352
rect 2832 2343 2834 2352
rect 2964 2372 3016 2378
rect 2780 2314 2832 2320
rect 2964 2314 3016 2320
rect 2976 480 3004 2314
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 480 3372 2246
rect 3528 1442 3556 2790
rect 4264 2514 4292 3130
rect 4356 2650 4384 8214
rect 4540 7886 4568 8230
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4632 6225 4660 14826
rect 4724 14414 4752 15846
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14618 4844 14758
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4724 13326 4752 14350
rect 4816 13530 4844 14554
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5000 13870 5028 14418
rect 4988 13864 5040 13870
rect 4986 13832 4988 13841
rect 5040 13832 5042 13841
rect 4896 13796 4948 13802
rect 4986 13767 5042 13776
rect 4896 13738 4948 13744
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4908 13326 4936 13738
rect 5092 13682 5120 15846
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 15026 5212 15302
rect 5354 15056 5410 15065
rect 5172 15020 5224 15026
rect 5354 14991 5410 15000
rect 5172 14962 5224 14968
rect 5184 14006 5212 14962
rect 5368 14822 5396 14991
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5000 13654 5120 13682
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 12714 4936 13262
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 5000 12356 5028 13654
rect 5184 13462 5212 13942
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5184 12986 5212 13398
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5552 12782 5580 13806
rect 5644 12850 5672 14214
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5540 12776 5592 12782
rect 5446 12744 5502 12753
rect 5540 12718 5592 12724
rect 5446 12679 5502 12688
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12481 5212 12582
rect 5170 12472 5226 12481
rect 5170 12407 5226 12416
rect 5460 12374 5488 12679
rect 5552 12442 5580 12718
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 4816 12328 5028 12356
rect 5448 12368 5500 12374
rect 5354 12336 5410 12345
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4724 9382 4752 10066
rect 4816 9568 4844 12328
rect 5172 12300 5224 12306
rect 5448 12310 5500 12316
rect 5354 12271 5356 12280
rect 5172 12242 5224 12248
rect 5408 12271 5410 12280
rect 5356 12242 5408 12248
rect 5184 11694 5212 12242
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 5000 10742 5028 11222
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 4816 9540 4936 9568
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 8498 4752 9318
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4618 6216 4674 6225
rect 4618 6151 4674 6160
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4448 4826 4476 5714
rect 4724 5370 4752 8298
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5778 4844 6054
rect 4908 5914 4936 9540
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4816 4672 4844 5578
rect 4908 5030 4936 5646
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 5000 4826 5028 10678
rect 5092 7546 5120 11562
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7342 5212 11630
rect 5276 11354 5304 12038
rect 5446 11792 5502 11801
rect 5356 11756 5408 11762
rect 5446 11727 5502 11736
rect 5356 11698 5408 11704
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5276 10810 5304 11290
rect 5368 11150 5396 11698
rect 5460 11694 5488 11727
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11286 5488 11494
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5368 10996 5396 11086
rect 5368 10968 5580 10996
rect 5552 10810 5580 10968
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5172 7336 5224 7342
rect 5092 7284 5172 7290
rect 5092 7278 5224 7284
rect 5092 7262 5212 7278
rect 5092 7002 5120 7262
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5092 5846 5120 6938
rect 5184 6322 5212 7142
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5276 6118 5304 10746
rect 5644 10130 5672 12650
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 9382 5580 9522
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 9178 5580 9318
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5644 8945 5672 10066
rect 5736 9450 5764 17190
rect 5908 17138 5960 17144
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5828 16590 5856 17070
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12753 5856 12786
rect 5814 12744 5870 12753
rect 5814 12679 5870 12688
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5828 11218 5856 12378
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 9518 5856 11154
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5630 8936 5686 8945
rect 5630 8871 5686 8880
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7274 5488 7686
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5644 7342 5672 7482
rect 5828 7410 5856 7890
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5368 6322 5396 6802
rect 5460 6798 5488 7210
rect 5538 7168 5594 7177
rect 5538 7103 5594 7112
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4896 4684 4948 4690
rect 4816 4644 4896 4672
rect 4896 4626 4948 4632
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4724 3738 4752 4490
rect 4802 4176 4858 4185
rect 4802 4111 4858 4120
rect 4816 3738 4844 4111
rect 4908 3942 4936 4626
rect 5000 4282 5028 4762
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4526 2952 4582 2961
rect 4724 2922 4752 3674
rect 4908 3602 4936 3878
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4526 2887 4582 2896
rect 4712 2916 4764 2922
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 4158 1456 4214 1465
rect 3528 1414 3832 1442
rect 3804 480 3832 1414
rect 4158 1391 4214 1400
rect 4172 480 4200 1391
rect 4540 480 4568 2887
rect 4712 2858 4764 2864
rect 5000 480 5028 3946
rect 5276 3738 5304 5850
rect 5368 4622 5396 6258
rect 5448 5704 5500 5710
rect 5446 5672 5448 5681
rect 5500 5672 5502 5681
rect 5446 5607 5502 5616
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4282 5396 4558
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5276 3641 5304 3674
rect 5262 3632 5318 3641
rect 5262 3567 5318 3576
rect 5276 2650 5304 3567
rect 5368 3534 5396 4218
rect 5460 4146 5488 4966
rect 5552 4826 5580 7103
rect 5724 6860 5776 6866
rect 5776 6820 5856 6848
rect 5724 6802 5776 6808
rect 5828 6118 5856 6820
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5846 5856 6054
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5920 5370 5948 16934
rect 6012 12442 6040 25350
rect 6196 24954 6224 25366
rect 6184 24948 6236 24954
rect 6184 24890 6236 24896
rect 6090 24848 6146 24857
rect 6090 24783 6146 24792
rect 6104 22098 6132 24783
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23730 6960 24006
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6840 23322 6868 23462
rect 6932 23322 6960 23666
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6288 22778 6316 23054
rect 6276 22772 6328 22778
rect 6196 22732 6276 22760
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6196 21146 6224 22732
rect 6276 22714 6328 22720
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6656 18970 6684 19178
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6196 17814 6224 18566
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6104 12714 6132 17682
rect 6196 17270 6224 17750
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6196 16794 6224 17206
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6196 15706 6224 16730
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6656 14550 6684 17138
rect 6748 17066 6776 22034
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 17202 6868 19110
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6920 16992 6972 16998
rect 6840 16940 6920 16946
rect 6840 16934 6972 16940
rect 6840 16918 6960 16934
rect 6840 16454 6868 16918
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16114 6868 16390
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 7024 14906 7052 26823
rect 7116 23254 7144 32506
rect 7208 31804 7236 34342
rect 7288 33040 7340 33046
rect 7288 32982 7340 32988
rect 7300 31958 7328 32982
rect 7392 32314 7420 34614
rect 7668 34542 7696 34886
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 7748 34468 7800 34474
rect 7748 34410 7800 34416
rect 7760 33969 7788 34410
rect 7746 33960 7802 33969
rect 7746 33895 7802 33904
rect 7656 33856 7708 33862
rect 7656 33798 7708 33804
rect 7562 33416 7618 33425
rect 7562 33351 7618 33360
rect 7576 33114 7604 33351
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7472 33040 7524 33046
rect 7470 33008 7472 33017
rect 7524 33008 7526 33017
rect 7470 32943 7526 32952
rect 7576 32570 7604 33050
rect 7564 32564 7616 32570
rect 7564 32506 7616 32512
rect 7472 32496 7524 32502
rect 7470 32464 7472 32473
rect 7524 32464 7526 32473
rect 7470 32399 7526 32408
rect 7392 32286 7512 32314
rect 7288 31952 7340 31958
rect 7288 31894 7340 31900
rect 7208 31776 7328 31804
rect 7300 31736 7328 31776
rect 7300 31708 7420 31736
rect 7288 30252 7340 30258
rect 7288 30194 7340 30200
rect 7196 30048 7248 30054
rect 7196 29990 7248 29996
rect 7208 29238 7236 29990
rect 7300 29850 7328 30194
rect 7288 29844 7340 29850
rect 7288 29786 7340 29792
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7392 27577 7420 31708
rect 7484 29102 7512 32286
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7576 31142 7604 31758
rect 7668 31754 7696 33798
rect 7760 33454 7788 33895
rect 7748 33448 7800 33454
rect 7748 33390 7800 33396
rect 7748 31884 7800 31890
rect 7748 31826 7800 31832
rect 7656 31748 7708 31754
rect 7656 31690 7708 31696
rect 7564 31136 7616 31142
rect 7564 31078 7616 31084
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 7472 28960 7524 28966
rect 7472 28902 7524 28908
rect 7484 28762 7512 28902
rect 7472 28756 7524 28762
rect 7472 28698 7524 28704
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7378 27568 7434 27577
rect 7378 27503 7434 27512
rect 7484 27441 7512 27950
rect 7576 27674 7604 31078
rect 7668 30938 7696 31690
rect 7760 31482 7788 31826
rect 7748 31476 7800 31482
rect 7748 31418 7800 31424
rect 7760 30938 7788 31418
rect 7656 30932 7708 30938
rect 7656 30874 7708 30880
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7668 30258 7696 30874
rect 7840 30320 7892 30326
rect 7840 30262 7892 30268
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 7564 27668 7616 27674
rect 7564 27610 7616 27616
rect 7470 27432 7526 27441
rect 7470 27367 7526 27376
rect 7288 27328 7340 27334
rect 7288 27270 7340 27276
rect 7300 27033 7328 27270
rect 7286 27024 7342 27033
rect 7668 26994 7696 30194
rect 7748 29640 7800 29646
rect 7748 29582 7800 29588
rect 7760 29073 7788 29582
rect 7746 29064 7802 29073
rect 7746 28999 7748 29008
rect 7800 28999 7802 29008
rect 7748 28970 7800 28976
rect 7746 28112 7802 28121
rect 7746 28047 7802 28056
rect 7760 27946 7788 28047
rect 7748 27940 7800 27946
rect 7748 27882 7800 27888
rect 7286 26959 7288 26968
rect 7340 26959 7342 26968
rect 7656 26988 7708 26994
rect 7288 26930 7340 26936
rect 7656 26930 7708 26936
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7208 25838 7236 26318
rect 7196 25832 7248 25838
rect 7196 25774 7248 25780
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7300 25265 7328 25638
rect 7286 25256 7342 25265
rect 7286 25191 7342 25200
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23662 7236 24006
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7300 23508 7328 23802
rect 7208 23480 7328 23508
rect 7104 23248 7156 23254
rect 7104 23190 7156 23196
rect 7116 23089 7144 23190
rect 7102 23080 7158 23089
rect 7102 23015 7158 23024
rect 7208 19258 7236 23480
rect 7392 23338 7420 26726
rect 7748 24336 7800 24342
rect 7748 24278 7800 24284
rect 7760 23866 7788 24278
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7300 23310 7420 23338
rect 7300 21418 7328 23310
rect 7470 23216 7526 23225
rect 7380 23180 7432 23186
rect 7470 23151 7526 23160
rect 7656 23180 7708 23186
rect 7380 23122 7432 23128
rect 7392 21962 7420 23122
rect 7484 22642 7512 23151
rect 7656 23122 7708 23128
rect 7668 22642 7696 23122
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7472 22636 7524 22642
rect 7656 22636 7708 22642
rect 7472 22578 7524 22584
rect 7576 22596 7656 22624
rect 7484 22234 7512 22578
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7484 21690 7512 22170
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7576 21486 7604 22596
rect 7656 22578 7708 22584
rect 7760 22098 7788 22646
rect 7852 22574 7880 30262
rect 7944 30190 7972 35686
rect 8116 35488 8168 35494
rect 8116 35430 8168 35436
rect 8024 31816 8076 31822
rect 8024 31758 8076 31764
rect 8036 31414 8064 31758
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 8128 30938 8156 35430
rect 8588 35272 8616 39520
rect 8956 37210 8984 39520
rect 8772 37182 8984 37210
rect 8668 35488 8720 35494
rect 8668 35430 8720 35436
rect 8404 35244 8616 35272
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 8220 33674 8248 34478
rect 8220 33658 8340 33674
rect 8220 33652 8352 33658
rect 8220 33646 8300 33652
rect 8300 33594 8352 33600
rect 8208 33380 8260 33386
rect 8208 33322 8260 33328
rect 8220 33130 8248 33322
rect 8220 33102 8340 33130
rect 8312 32774 8340 33102
rect 8300 32768 8352 32774
rect 8300 32710 8352 32716
rect 8312 31686 8340 32710
rect 8404 32473 8432 35244
rect 8484 35148 8536 35154
rect 8484 35090 8536 35096
rect 8496 34542 8524 35090
rect 8484 34536 8536 34542
rect 8484 34478 8536 34484
rect 8390 32464 8446 32473
rect 8390 32399 8446 32408
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 8128 30326 8156 30874
rect 8312 30666 8340 31622
rect 8392 30728 8444 30734
rect 8392 30670 8444 30676
rect 8300 30660 8352 30666
rect 8300 30602 8352 30608
rect 8116 30320 8168 30326
rect 8116 30262 8168 30268
rect 7932 30184 7984 30190
rect 7932 30126 7984 30132
rect 8312 30054 8340 30602
rect 8300 30048 8352 30054
rect 8128 29996 8300 30002
rect 8128 29990 8352 29996
rect 8128 29974 8340 29990
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 7932 29504 7984 29510
rect 7932 29446 7984 29452
rect 7944 27606 7972 29446
rect 8036 29306 8064 29650
rect 8128 29322 8156 29974
rect 8404 29510 8432 30670
rect 8392 29504 8444 29510
rect 8392 29446 8444 29452
rect 8128 29306 8340 29322
rect 8024 29300 8076 29306
rect 8024 29242 8076 29248
rect 8128 29300 8352 29306
rect 8128 29294 8300 29300
rect 8024 27872 8076 27878
rect 8024 27814 8076 27820
rect 8036 27674 8064 27814
rect 8024 27668 8076 27674
rect 8024 27610 8076 27616
rect 7932 27600 7984 27606
rect 7932 27542 7984 27548
rect 7944 26586 7972 27542
rect 8036 27130 8064 27610
rect 8128 27470 8156 29294
rect 8300 29242 8352 29248
rect 8208 29232 8260 29238
rect 8208 29174 8260 29180
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 8128 27062 8156 27406
rect 8116 27056 8168 27062
rect 8116 26998 8168 27004
rect 7932 26580 7984 26586
rect 7932 26522 7984 26528
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7944 24750 7972 25094
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7944 23866 7972 24686
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 8036 24206 8064 24550
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 7932 23860 7984 23866
rect 7932 23802 7984 23808
rect 7944 22778 7972 23802
rect 8036 23798 8064 24142
rect 8024 23792 8076 23798
rect 8024 23734 8076 23740
rect 8036 23186 8064 23734
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8024 23180 8076 23186
rect 8024 23122 8076 23128
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 7852 22114 7880 22510
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 7748 22092 7800 22098
rect 7852 22086 7972 22114
rect 7748 22034 7800 22040
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7668 21434 7696 22034
rect 7288 21412 7340 21418
rect 7288 21354 7340 21360
rect 7576 21146 7604 21422
rect 7668 21406 7880 21434
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7746 21312 7802 21321
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7576 20058 7604 21082
rect 7668 21010 7696 21286
rect 7746 21247 7802 21256
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7760 20942 7788 21247
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 7760 20262 7788 20878
rect 7852 20806 7880 21406
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7852 20602 7880 20742
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 6932 14878 7052 14906
rect 7116 19230 7236 19258
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14618 6868 14758
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6644 14544 6696 14550
rect 6550 14512 6606 14521
rect 6644 14486 6696 14492
rect 6550 14447 6606 14456
rect 6564 13818 6592 14447
rect 6656 14006 6684 14486
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6748 13870 6776 14350
rect 6840 14074 6868 14554
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6736 13864 6788 13870
rect 6564 13790 6684 13818
rect 6736 13806 6788 13812
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6012 11354 6040 12174
rect 6104 11898 6132 12174
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6104 10810 6132 11630
rect 6196 11286 6224 12310
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6472 10577 6500 11154
rect 6458 10568 6514 10577
rect 6458 10503 6460 10512
rect 6512 10503 6514 10512
rect 6460 10474 6512 10480
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6656 10248 6684 13790
rect 6748 12238 6776 13806
rect 6932 13394 6960 14878
rect 7012 14816 7064 14822
rect 7116 14804 7144 19230
rect 7300 19174 7328 19654
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7208 18970 7236 19110
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7208 16250 7236 18906
rect 7300 16794 7328 19110
rect 7484 17882 7512 19314
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7668 18358 7696 18634
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7760 18170 7788 20198
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 18329 7880 18566
rect 7838 18320 7894 18329
rect 7838 18255 7894 18264
rect 7760 18142 7880 18170
rect 7654 17912 7710 17921
rect 7472 17876 7524 17882
rect 7392 17836 7472 17864
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7300 16114 7328 16186
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 15026 7236 15302
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7064 14776 7144 14804
rect 7012 14758 7064 14764
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 12374 6868 12854
rect 6932 12782 6960 13126
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6828 11756 6880 11762
rect 6932 11744 6960 12378
rect 7024 12322 7052 14758
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 7116 12646 7144 13738
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12442 7144 12582
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7024 12294 7144 12322
rect 6880 11716 6960 11744
rect 6828 11698 6880 11704
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 10470 7052 10950
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6196 10220 6684 10248
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5920 5166 5948 5306
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5448 4140 5500 4146
rect 5500 4100 5580 4128
rect 5448 4082 5500 4088
rect 5552 3777 5580 4100
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5538 3768 5594 3777
rect 5644 3738 5672 4014
rect 5538 3703 5594 3712
rect 5632 3732 5684 3738
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5354 2816 5410 2825
rect 5354 2751 5410 2760
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5264 2304 5316 2310
rect 5262 2272 5264 2281
rect 5316 2272 5318 2281
rect 5262 2207 5318 2216
rect 5368 480 5396 2751
rect 5460 2446 5488 3334
rect 5552 3194 5580 3703
rect 5632 3674 5684 3680
rect 5630 3496 5686 3505
rect 5630 3431 5686 3440
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5644 2650 5672 3431
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5736 480 5764 4014
rect 5828 610 5856 4966
rect 5920 3670 5948 5102
rect 6012 4010 6040 9046
rect 6196 7818 6224 10220
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6656 8362 6684 9318
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6932 8090 6960 8366
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 6934 6132 7686
rect 6196 7478 6224 7754
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6656 7002 6684 7210
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6458 6224 6802
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6196 5914 6224 6394
rect 6748 6066 6776 7414
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 6458 6868 7346
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6656 6038 6776 6066
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6288 5098 6316 5782
rect 6656 5778 6684 6038
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6656 5658 6684 5714
rect 6564 5630 6684 5658
rect 6564 5234 6592 5630
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6656 4826 6684 5510
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6748 4622 6776 5850
rect 6826 5672 6882 5681
rect 6932 5658 6960 7142
rect 7024 5828 7052 10406
rect 7116 8129 7144 12294
rect 7208 11354 7236 12718
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7300 10130 7328 15642
rect 7392 15026 7420 17836
rect 7654 17847 7710 17856
rect 7472 17818 7524 17824
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 15910 7512 17002
rect 7668 16794 7696 17847
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7668 16674 7696 16730
rect 7576 16646 7696 16674
rect 7576 16250 7604 16646
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7760 16114 7788 16526
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7654 16008 7710 16017
rect 7564 15972 7616 15978
rect 7654 15943 7710 15952
rect 7564 15914 7616 15920
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 12986 7420 14962
rect 7484 14346 7512 15846
rect 7576 15706 7604 15914
rect 7668 15706 7696 15943
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7562 15600 7618 15609
rect 7562 15535 7564 15544
rect 7616 15535 7618 15544
rect 7564 15506 7616 15512
rect 7576 14618 7604 15506
rect 7668 15162 7696 15642
rect 7760 15502 7788 16050
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7760 14618 7788 15438
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7576 14498 7604 14554
rect 7576 14470 7788 14498
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7392 11694 7420 12922
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 11150 7420 11630
rect 7484 11558 7512 12310
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11286 7512 11494
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7576 10010 7604 14350
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7208 9982 7604 10010
rect 7102 8120 7158 8129
rect 7102 8055 7158 8064
rect 7102 6760 7158 6769
rect 7102 6695 7158 6704
rect 7116 6458 7144 6695
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7116 6254 7144 6394
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7208 5896 7236 9982
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7392 9518 7420 9862
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8634 7328 9318
rect 7392 9178 7420 9454
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7300 7342 7328 8570
rect 7378 7984 7434 7993
rect 7378 7919 7434 7928
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7392 7290 7420 7919
rect 7484 7410 7512 9862
rect 7668 8537 7696 14282
rect 7654 8528 7710 8537
rect 7654 8463 7710 8472
rect 7760 8378 7788 14470
rect 7576 8350 7788 8378
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7392 7262 7512 7290
rect 7208 5868 7328 5896
rect 7024 5800 7236 5828
rect 6882 5630 6960 5658
rect 6826 5607 6882 5616
rect 6840 4690 6868 5607
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4616 6788 4622
rect 6182 4584 6238 4593
rect 6736 4558 6788 4564
rect 6182 4519 6238 4528
rect 6644 4548 6696 4554
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 6012 3738 6040 3946
rect 6196 3738 6224 4519
rect 6644 4490 6696 4496
rect 6656 4128 6684 4490
rect 6748 4282 6776 4558
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4282 6868 4422
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6932 4162 6960 4966
rect 7208 4570 7236 5800
rect 6840 4134 6960 4162
rect 7024 4542 7236 4570
rect 6656 4100 6776 4128
rect 6748 3924 6776 4100
rect 6840 4078 6868 4134
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6932 3924 6960 4014
rect 6748 3896 6960 3924
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 3194 5948 3606
rect 5908 3188 5960 3194
rect 6748 3176 6776 3896
rect 6920 3188 6972 3194
rect 6748 3148 6920 3176
rect 5908 3130 5960 3136
rect 6920 3130 6972 3136
rect 6642 3088 6698 3097
rect 6642 3023 6698 3032
rect 6918 3088 6974 3097
rect 6918 3023 6974 3032
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6656 1170 6684 3023
rect 6734 2816 6790 2825
rect 6734 2751 6790 2760
rect 6748 2650 6776 2751
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6564 1142 6684 1170
rect 5816 604 5868 610
rect 5816 546 5868 552
rect 6184 604 6236 610
rect 6184 546 6236 552
rect 6196 480 6224 546
rect 6564 480 6592 1142
rect 6932 480 6960 3023
rect 7024 2514 7052 4542
rect 7300 4468 7328 5868
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7392 4690 7420 5170
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7116 4440 7328 4468
rect 7380 4480 7432 4486
rect 7116 3505 7144 4440
rect 7380 4422 7432 4428
rect 7392 4214 7420 4422
rect 7380 4208 7432 4214
rect 7286 4176 7342 4185
rect 7380 4150 7432 4156
rect 7286 4111 7288 4120
rect 7340 4111 7342 4120
rect 7288 4082 7340 4088
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7102 3496 7158 3505
rect 7208 3466 7236 3878
rect 7286 3768 7342 3777
rect 7286 3703 7342 3712
rect 7102 3431 7158 3440
rect 7196 3460 7248 3466
rect 7116 2582 7144 3431
rect 7196 3402 7248 3408
rect 7300 3126 7328 3703
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7300 2922 7328 3062
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1465 7144 2246
rect 7102 1456 7158 1465
rect 7102 1391 7158 1400
rect 7392 480 7420 3946
rect 7484 3738 7512 7262
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7484 2990 7512 3674
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7576 2825 7604 8350
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7410 7696 8230
rect 7852 7562 7880 18142
rect 7944 15337 7972 22086
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 8036 21146 8064 22034
rect 8128 22030 8156 23530
rect 8116 22024 8168 22030
rect 8220 22001 8248 29174
rect 8392 29096 8444 29102
rect 8298 29064 8354 29073
rect 8392 29038 8444 29044
rect 8298 28999 8354 29008
rect 8312 23254 8340 28999
rect 8404 28626 8432 29038
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 8404 28393 8432 28562
rect 8390 28384 8446 28393
rect 8390 28319 8446 28328
rect 8392 28212 8444 28218
rect 8392 28154 8444 28160
rect 8404 26602 8432 28154
rect 8496 26790 8524 34478
rect 8576 34400 8628 34406
rect 8576 34342 8628 34348
rect 8588 32570 8616 34342
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 8576 31340 8628 31346
rect 8576 31282 8628 31288
rect 8588 30870 8616 31282
rect 8576 30864 8628 30870
rect 8680 30841 8708 35430
rect 8772 31346 8800 37182
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8852 33652 8904 33658
rect 8852 33594 8904 33600
rect 8864 32570 8892 33594
rect 9416 33017 9444 39520
rect 9680 36236 9732 36242
rect 9680 36178 9732 36184
rect 9692 35873 9720 36178
rect 9678 35864 9734 35873
rect 9600 35834 9678 35850
rect 9588 35828 9678 35834
rect 9640 35822 9678 35828
rect 9678 35799 9734 35808
rect 9588 35770 9640 35776
rect 9692 35739 9720 35799
rect 9496 35148 9548 35154
rect 9496 35090 9548 35096
rect 9508 34406 9536 35090
rect 9680 35080 9732 35086
rect 9680 35022 9732 35028
rect 9692 34542 9720 35022
rect 9680 34536 9732 34542
rect 9680 34478 9732 34484
rect 9496 34400 9548 34406
rect 9496 34342 9548 34348
rect 9508 34202 9536 34342
rect 9496 34196 9548 34202
rect 9496 34138 9548 34144
rect 9402 33008 9458 33017
rect 9458 32966 9720 32994
rect 9402 32943 9458 32952
rect 9416 32883 9444 32943
rect 9588 32904 9640 32910
rect 9588 32846 9640 32852
rect 9496 32836 9548 32842
rect 9496 32778 9548 32784
rect 9404 32768 9456 32774
rect 9404 32710 9456 32716
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8852 32564 8904 32570
rect 8852 32506 8904 32512
rect 8864 31822 8892 32506
rect 9416 32366 9444 32710
rect 9508 32434 9536 32778
rect 9496 32428 9548 32434
rect 9496 32370 9548 32376
rect 9404 32360 9456 32366
rect 9404 32302 9456 32308
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 9312 31680 9364 31686
rect 9312 31622 9364 31628
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9324 31346 9352 31622
rect 9416 31482 9444 32302
rect 9404 31476 9456 31482
rect 9404 31418 9456 31424
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 9312 31340 9364 31346
rect 9312 31282 9364 31288
rect 9600 31278 9628 32846
rect 9692 32570 9720 32966
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9588 31272 9640 31278
rect 9310 31240 9366 31249
rect 9588 31214 9640 31220
rect 9310 31175 9366 31184
rect 9324 31142 9352 31175
rect 9312 31136 9364 31142
rect 9312 31078 9364 31084
rect 8576 30806 8628 30812
rect 8666 30832 8722 30841
rect 8588 29866 8616 30806
rect 8666 30767 8722 30776
rect 8680 30036 8708 30767
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8760 30048 8812 30054
rect 8680 30008 8760 30036
rect 8760 29990 8812 29996
rect 8588 29838 8708 29866
rect 8680 29714 8708 29838
rect 8668 29708 8720 29714
rect 8668 29650 8720 29656
rect 8576 29640 8628 29646
rect 8576 29582 8628 29588
rect 8588 29034 8616 29582
rect 8576 29028 8628 29034
rect 8576 28970 8628 28976
rect 8588 28762 8616 28970
rect 8576 28756 8628 28762
rect 8576 28698 8628 28704
rect 8588 28082 8616 28698
rect 8576 28076 8628 28082
rect 8576 28018 8628 28024
rect 8576 27872 8628 27878
rect 8574 27840 8576 27849
rect 8628 27840 8630 27849
rect 8574 27775 8630 27784
rect 8680 27470 8708 29650
rect 8668 27464 8720 27470
rect 8668 27406 8720 27412
rect 8484 26784 8536 26790
rect 8484 26726 8536 26732
rect 8404 26574 8524 26602
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8404 23322 8432 24006
rect 8392 23316 8444 23322
rect 8392 23258 8444 23264
rect 8300 23248 8352 23254
rect 8300 23190 8352 23196
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 8312 22098 8340 23054
rect 8404 22778 8432 23258
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8116 21966 8168 21972
rect 8206 21992 8262 22001
rect 8128 21350 8156 21966
rect 8206 21927 8262 21936
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8220 21162 8248 21626
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8128 21134 8248 21162
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 8036 18222 8064 19246
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7930 15328 7986 15337
rect 7930 15263 7986 15272
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7944 14414 7972 15098
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8036 14074 8064 17478
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7944 13530 7972 13806
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 8036 12986 8064 13330
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8128 11014 8156 21134
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8220 20602 8248 20946
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8208 19304 8260 19310
rect 8312 19292 8340 20198
rect 8260 19264 8340 19292
rect 8392 19304 8444 19310
rect 8208 19246 8260 19252
rect 8392 19246 8444 19252
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8220 17678 8248 18770
rect 8312 18766 8340 19110
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8312 18426 8340 18702
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8404 18154 8432 19246
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8220 14618 8248 17614
rect 8312 17490 8340 18022
rect 8404 17610 8432 18090
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 8312 17462 8432 17490
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8220 13462 8248 14010
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10713 8156 10950
rect 8114 10704 8170 10713
rect 8114 10639 8170 10648
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7944 9489 7972 10066
rect 8036 9994 8064 10406
rect 8114 10296 8170 10305
rect 8114 10231 8116 10240
rect 8168 10231 8170 10240
rect 8116 10202 8168 10208
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8036 9586 8064 9930
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7930 9480 7986 9489
rect 7930 9415 7986 9424
rect 7944 7993 7972 9415
rect 8036 8362 8064 9522
rect 8128 9110 8156 10202
rect 8312 9382 8340 17206
rect 8404 17134 8432 17462
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8496 16998 8524 26574
rect 8668 26240 8720 26246
rect 8668 26182 8720 26188
rect 8576 25968 8628 25974
rect 8574 25936 8576 25945
rect 8628 25936 8630 25945
rect 8574 25871 8630 25880
rect 8680 25838 8708 26182
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8772 25650 8800 29990
rect 8850 29744 8906 29753
rect 8850 29679 8906 29688
rect 8864 28218 8892 29679
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8852 28212 8904 28218
rect 8852 28154 8904 28160
rect 9324 27713 9352 31078
rect 9600 30870 9628 31214
rect 9692 30938 9720 32302
rect 9680 30932 9732 30938
rect 9680 30874 9732 30880
rect 9588 30864 9640 30870
rect 9588 30806 9640 30812
rect 9784 30326 9812 39520
rect 9862 36408 9918 36417
rect 9862 36343 9864 36352
rect 9916 36343 9918 36352
rect 9864 36314 9916 36320
rect 9864 35760 9916 35766
rect 9862 35728 9864 35737
rect 9916 35728 9918 35737
rect 9862 35663 9918 35672
rect 10152 35578 10180 39520
rect 10152 35550 10364 35578
rect 9956 34400 10008 34406
rect 9956 34342 10008 34348
rect 9968 34202 9996 34342
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9968 33969 9996 34138
rect 9954 33960 10010 33969
rect 9954 33895 10010 33904
rect 10140 33448 10192 33454
rect 10138 33416 10140 33425
rect 10192 33416 10194 33425
rect 10138 33351 10194 33360
rect 10232 33380 10284 33386
rect 10232 33322 10284 33328
rect 10048 32972 10100 32978
rect 10048 32914 10100 32920
rect 10060 32026 10088 32914
rect 10140 32564 10192 32570
rect 10140 32506 10192 32512
rect 10048 32020 10100 32026
rect 10048 31962 10100 31968
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 9772 30320 9824 30326
rect 9772 30262 9824 30268
rect 9772 30184 9824 30190
rect 9772 30126 9824 30132
rect 9680 30116 9732 30122
rect 9680 30058 9732 30064
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9416 28218 9444 29446
rect 9496 29232 9548 29238
rect 9600 29209 9628 29990
rect 9496 29174 9548 29180
rect 9586 29200 9642 29209
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9310 27704 9366 27713
rect 9310 27639 9366 27648
rect 8852 27464 8904 27470
rect 8852 27406 8904 27412
rect 8864 26790 8892 27406
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9508 26994 9536 29174
rect 9586 29135 9642 29144
rect 9586 28112 9642 28121
rect 9586 28047 9642 28056
rect 9600 27946 9628 28047
rect 9588 27940 9640 27946
rect 9588 27882 9640 27888
rect 9600 27606 9628 27882
rect 9692 27849 9720 30058
rect 9784 30054 9812 30126
rect 9772 30048 9824 30054
rect 9772 29990 9824 29996
rect 9784 29510 9812 29990
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9678 27840 9734 27849
rect 9678 27775 9734 27784
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 9678 27432 9734 27441
rect 9588 27396 9640 27402
rect 9784 27418 9812 29446
rect 9734 27390 9812 27418
rect 9678 27367 9734 27376
rect 9588 27338 9640 27344
rect 9496 26988 9548 26994
rect 9496 26930 9548 26936
rect 9600 26926 9628 27338
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 9312 26784 9364 26790
rect 9692 26772 9720 27367
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9692 26744 9812 26772
rect 9312 26726 9364 26732
rect 8588 25622 8800 25650
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8390 16688 8446 16697
rect 8390 16623 8446 16632
rect 8404 16590 8432 16623
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8404 16250 8432 16526
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8404 15570 8432 16186
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8404 13870 8432 14962
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8404 13258 8432 13806
rect 8496 13530 8524 14350
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8496 12986 8524 13262
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8404 9160 8432 12854
rect 8482 12744 8538 12753
rect 8482 12679 8538 12688
rect 8496 12442 8524 12679
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8588 10146 8616 25622
rect 8668 24676 8720 24682
rect 8668 24618 8720 24624
rect 8680 23662 8708 24618
rect 8668 23656 8720 23662
rect 8668 23598 8720 23604
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8680 22710 8708 23190
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8680 22574 8708 22646
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8680 20942 8708 22510
rect 8760 22432 8812 22438
rect 8864 22420 8892 26726
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9324 25770 9352 26726
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9312 25764 9364 25770
rect 9312 25706 9364 25712
rect 9324 25498 9352 25706
rect 9312 25492 9364 25498
rect 9312 25434 9364 25440
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9416 24993 9444 25842
rect 9402 24984 9458 24993
rect 9402 24919 9458 24928
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9140 23118 9168 23598
rect 9324 23526 9352 24278
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9416 23662 9444 24006
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9312 23520 9364 23526
rect 9312 23462 9364 23468
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8812 22392 8892 22420
rect 8760 22374 8812 22380
rect 8772 21894 8800 22374
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8666 20768 8722 20777
rect 8666 20703 8722 20712
rect 8680 17270 8708 20703
rect 8772 19258 8800 21830
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 9324 21672 9352 23462
rect 9416 23361 9444 23598
rect 9402 23352 9458 23361
rect 9402 23287 9458 23296
rect 9678 23080 9734 23089
rect 9678 23015 9734 23024
rect 9692 22386 9720 23015
rect 9784 22506 9812 26744
rect 9876 26246 9904 26930
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9876 26042 9904 26182
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 9968 23746 9996 31078
rect 10046 30832 10102 30841
rect 10046 30767 10048 30776
rect 10100 30767 10102 30776
rect 10048 30738 10100 30744
rect 10048 30320 10100 30326
rect 10048 30262 10100 30268
rect 10060 29034 10088 30262
rect 10048 29028 10100 29034
rect 10048 28970 10100 28976
rect 10046 27568 10102 27577
rect 10152 27554 10180 32506
rect 10244 32026 10272 33322
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 10244 30734 10272 31282
rect 10232 30728 10284 30734
rect 10232 30670 10284 30676
rect 10244 30394 10272 30670
rect 10232 30388 10284 30394
rect 10232 30330 10284 30336
rect 10232 30116 10284 30122
rect 10232 30058 10284 30064
rect 10244 29646 10272 30058
rect 10232 29640 10284 29646
rect 10232 29582 10284 29588
rect 10244 29034 10272 29582
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 10244 28626 10272 28970
rect 10232 28620 10284 28626
rect 10232 28562 10284 28568
rect 10152 27526 10272 27554
rect 10046 27503 10048 27512
rect 10100 27503 10102 27512
rect 10048 27474 10100 27480
rect 10060 27418 10088 27474
rect 10060 27390 10180 27418
rect 10152 27130 10180 27390
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10152 24562 10180 27066
rect 10244 24682 10272 27526
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10152 24534 10272 24562
rect 10244 24410 10272 24534
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10152 23798 10180 24210
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 10244 23866 10272 24142
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 9876 23718 9996 23746
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 9772 22500 9824 22506
rect 9772 22442 9824 22448
rect 9600 22358 9720 22386
rect 9770 22400 9826 22409
rect 9600 22216 9628 22358
rect 9770 22335 9826 22344
rect 9784 22250 9812 22335
rect 9692 22222 9812 22250
rect 9692 22216 9720 22222
rect 9600 22188 9720 22216
rect 9402 22128 9458 22137
rect 9402 22063 9458 22072
rect 9586 22128 9642 22137
rect 9770 22128 9826 22137
rect 9642 22072 9770 22080
rect 9586 22063 9826 22072
rect 9416 21978 9444 22063
rect 9600 22052 9812 22063
rect 9407 21950 9444 21978
rect 9407 21842 9435 21950
rect 9772 21888 9824 21894
rect 9678 21856 9734 21865
rect 9407 21814 9444 21842
rect 9232 21644 9352 21672
rect 9232 21010 9260 21644
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 19394 8892 19654
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8864 19366 9076 19394
rect 8772 19230 8984 19258
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8668 17264 8720 17270
rect 8668 17206 8720 17212
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8496 10130 8616 10146
rect 8484 10124 8616 10130
rect 8536 10118 8616 10124
rect 8484 10066 8536 10072
rect 8496 9450 8524 10066
rect 8680 10033 8708 16730
rect 8772 16250 8800 19110
rect 8956 18714 8984 19230
rect 9048 19174 9076 19366
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8864 18686 8984 18714
rect 8864 16250 8892 18686
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9232 16658 9260 17070
rect 9324 16794 9352 21354
rect 9416 21146 9444 21814
rect 9600 21814 9678 21842
rect 9600 21457 9628 21814
rect 9876 21865 9904 23718
rect 10152 23576 10180 23734
rect 9968 23548 10180 23576
rect 9772 21830 9824 21836
rect 9862 21856 9918 21865
rect 9678 21791 9734 21800
rect 9784 21672 9812 21830
rect 9862 21791 9918 21800
rect 9692 21644 9812 21672
rect 9862 21720 9918 21729
rect 9862 21655 9918 21664
rect 9586 21448 9642 21457
rect 9586 21383 9642 21392
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8864 15978 8892 16186
rect 9416 16046 9444 20946
rect 9588 20936 9640 20942
rect 9692 20913 9720 21644
rect 9770 21584 9826 21593
rect 9770 21519 9826 21528
rect 9784 21078 9812 21519
rect 9772 21072 9824 21078
rect 9772 21014 9824 21020
rect 9588 20878 9640 20884
rect 9678 20904 9734 20913
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9508 19718 9536 20266
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 18698 9536 19654
rect 9600 19258 9628 20878
rect 9678 20839 9734 20848
rect 9876 19310 9904 21655
rect 9864 19304 9916 19310
rect 9600 19230 9812 19258
rect 9864 19246 9916 19252
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9508 18426 9536 18634
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9600 17762 9628 19110
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9692 17882 9720 18566
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9600 17734 9720 17762
rect 9784 17746 9812 19230
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9876 18834 9904 19110
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9876 18086 9904 18634
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17921 9904 18022
rect 9862 17912 9918 17921
rect 9862 17847 9918 17856
rect 9692 17610 9720 17734
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9508 17134 9536 17478
rect 9496 17128 9548 17134
rect 9494 17096 9496 17105
rect 9548 17096 9550 17105
rect 9784 17066 9812 17682
rect 9494 17031 9550 17040
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9496 16992 9548 16998
rect 9876 16946 9904 17847
rect 9496 16934 9548 16940
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 8864 15706 8892 15914
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8772 14074 8800 14350
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8666 10024 8722 10033
rect 8666 9959 8722 9968
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8404 9132 8524 9160
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8114 8528 8170 8537
rect 8114 8463 8170 8472
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7930 7984 7986 7993
rect 7930 7919 7986 7928
rect 7760 7534 7880 7562
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 2938 7696 6054
rect 7760 5370 7788 7534
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7746 5264 7802 5273
rect 7746 5199 7748 5208
rect 7800 5199 7802 5208
rect 7748 5170 7800 5176
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 3398 7788 4966
rect 7852 4826 7880 6598
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7852 3738 7880 4762
rect 7944 3942 7972 6666
rect 8036 4146 8064 8298
rect 8128 7886 8156 8463
rect 8220 7954 8248 8842
rect 8312 8566 8340 8910
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 8022 8340 8502
rect 8404 8090 8432 8978
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8390 7984 8446 7993
rect 8208 7948 8260 7954
rect 8390 7919 8392 7928
rect 8208 7890 8260 7896
rect 8444 7919 8446 7928
rect 8392 7890 8444 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7546 8156 7822
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 6118 8156 6190
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 8128 3890 8156 6054
rect 8220 5914 8248 6802
rect 8312 6361 8340 7754
rect 8404 7546 8432 7890
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8298 6352 8354 6361
rect 8298 6287 8354 6296
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5914 8340 6054
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8220 5409 8248 5714
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8206 5400 8262 5409
rect 8206 5335 8262 5344
rect 8206 5264 8262 5273
rect 8206 5199 8262 5208
rect 8220 5166 8248 5199
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8312 4842 8340 5510
rect 8220 4814 8340 4842
rect 8220 4010 8248 4814
rect 8300 4752 8352 4758
rect 8404 4729 8432 6598
rect 8300 4694 8352 4700
rect 8390 4720 8446 4729
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8312 3942 8340 4694
rect 8390 4655 8446 4664
rect 8300 3936 8352 3942
rect 8128 3862 8248 3890
rect 8300 3878 8352 3884
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3058 7788 3334
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7668 2910 7880 2938
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7852 2666 7880 2910
rect 7944 2825 7972 3538
rect 7930 2816 7986 2825
rect 7930 2751 7986 2760
rect 7760 2638 7880 2666
rect 8116 2644 8168 2650
rect 7760 480 7788 2638
rect 8116 2586 8168 2592
rect 8128 2553 8156 2586
rect 8114 2544 8170 2553
rect 8114 2479 8170 2488
rect 8220 480 8248 3862
rect 8496 3738 8524 9132
rect 8588 5778 8616 9318
rect 8772 8430 8800 9454
rect 8864 8634 8892 15506
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9324 15026 9352 15914
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14482 9352 14758
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9324 13530 9352 14418
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9324 12442 9352 12650
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 9324 9450 9352 9862
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8680 6746 8708 7414
rect 8772 7342 8800 7822
rect 8760 7336 8812 7342
rect 8758 7304 8760 7313
rect 8812 7304 8814 7313
rect 8758 7239 8814 7248
rect 8864 6905 8892 8570
rect 9310 8392 9366 8401
rect 9310 8327 9312 8336
rect 9364 8327 9366 8336
rect 9312 8298 9364 8304
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8850 6896 8906 6905
rect 8850 6831 8906 6840
rect 8680 6718 8800 6746
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8680 6322 8708 6598
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8680 5574 8708 6258
rect 8668 5568 8720 5574
rect 8588 5528 8668 5556
rect 8588 5098 8616 5528
rect 8668 5510 8720 5516
rect 8666 5128 8722 5137
rect 8576 5092 8628 5098
rect 8666 5063 8722 5072
rect 8576 5034 8628 5040
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8496 3194 8524 3674
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8312 2009 8340 3130
rect 8482 2680 8538 2689
rect 8482 2615 8484 2624
rect 8536 2615 8538 2624
rect 8484 2586 8536 2592
rect 8680 2564 8708 5063
rect 8772 3777 8800 6718
rect 8864 6186 8892 6831
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9324 6254 9352 8298
rect 9416 7750 9444 15982
rect 9508 12594 9536 16934
rect 9784 16918 9904 16946
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9600 16114 9628 16662
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9600 14890 9628 15438
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9600 14618 9628 14826
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9692 13818 9720 14894
rect 9600 13790 9720 13818
rect 9600 12753 9628 13790
rect 9586 12744 9642 12753
rect 9586 12679 9642 12688
rect 9680 12640 9732 12646
rect 9508 12566 9628 12594
rect 9680 12582 9732 12588
rect 9494 12472 9550 12481
rect 9494 12407 9550 12416
rect 9508 10305 9536 12407
rect 9494 10296 9550 10305
rect 9494 10231 9550 10240
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9508 7426 9536 9318
rect 9600 8838 9628 12566
rect 9692 12374 9720 12582
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9784 12306 9812 16918
rect 9968 13002 9996 23548
rect 10230 23352 10286 23361
rect 10230 23287 10286 23296
rect 10048 22500 10100 22506
rect 10048 22442 10100 22448
rect 10060 21486 10088 22442
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22166 10180 22374
rect 10244 22166 10272 23287
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 10336 22012 10364 35550
rect 10416 35488 10468 35494
rect 10416 35430 10468 35436
rect 10428 32230 10456 35430
rect 10506 32464 10562 32473
rect 10506 32399 10562 32408
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10520 32026 10548 32399
rect 10508 32020 10560 32026
rect 10508 31962 10560 31968
rect 10414 31920 10470 31929
rect 10414 31855 10470 31864
rect 10428 31822 10456 31855
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10428 31142 10456 31758
rect 10520 31142 10548 31962
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10520 29714 10548 30194
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10414 29064 10470 29073
rect 10414 28999 10416 29008
rect 10468 28999 10470 29008
rect 10416 28970 10468 28976
rect 10520 28490 10548 29650
rect 10508 28484 10560 28490
rect 10508 28426 10560 28432
rect 10506 27840 10562 27849
rect 10506 27775 10562 27784
rect 10416 26784 10468 26790
rect 10416 26726 10468 26732
rect 10244 21984 10364 22012
rect 10138 21856 10194 21865
rect 10138 21791 10194 21800
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10046 20360 10102 20369
rect 10046 20295 10102 20304
rect 10060 20058 10088 20295
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10060 19174 10088 19858
rect 10048 19168 10100 19174
rect 10152 19145 10180 21791
rect 10048 19110 10100 19116
rect 10138 19136 10194 19145
rect 10138 19071 10194 19080
rect 10244 19009 10272 21984
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10336 21622 10364 21830
rect 10324 21616 10376 21622
rect 10324 21558 10376 21564
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10230 19000 10286 19009
rect 10336 18970 10364 21422
rect 10230 18935 10286 18944
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10336 18426 10364 18906
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10336 17762 10364 18362
rect 10244 17734 10364 17762
rect 10244 16697 10272 17734
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10336 17338 10364 17614
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10336 16794 10364 17274
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10230 16688 10286 16697
rect 10230 16623 10286 16632
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10244 13394 10272 16186
rect 10324 16176 10376 16182
rect 10322 16144 10324 16153
rect 10376 16144 10378 16153
rect 10322 16079 10378 16088
rect 10428 14958 10456 26726
rect 10520 22778 10548 27775
rect 10612 26625 10640 39520
rect 10980 35714 11008 39520
rect 10704 35686 11008 35714
rect 10704 30977 10732 35686
rect 11152 34944 11204 34950
rect 11152 34886 11204 34892
rect 11164 34474 11192 34886
rect 11152 34468 11204 34474
rect 11152 34410 11204 34416
rect 10876 34128 10928 34134
rect 10876 34070 10928 34076
rect 10784 34060 10836 34066
rect 10784 34002 10836 34008
rect 10796 33658 10824 34002
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10782 33552 10838 33561
rect 10782 33487 10838 33496
rect 10796 33114 10824 33487
rect 10784 33108 10836 33114
rect 10784 33050 10836 33056
rect 10784 32836 10836 32842
rect 10784 32778 10836 32784
rect 10796 31822 10824 32778
rect 10888 32570 10916 34070
rect 10968 33992 11020 33998
rect 10968 33934 11020 33940
rect 10980 32774 11008 33934
rect 11060 33856 11112 33862
rect 11060 33798 11112 33804
rect 11072 33114 11100 33798
rect 11060 33108 11112 33114
rect 11060 33050 11112 33056
rect 10968 32768 11020 32774
rect 10968 32710 11020 32716
rect 10876 32564 10928 32570
rect 10876 32506 10928 32512
rect 11072 32026 11100 33050
rect 11164 32842 11192 34410
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 11256 33454 11284 34138
rect 11244 33448 11296 33454
rect 11244 33390 11296 33396
rect 11152 32836 11204 32842
rect 11152 32778 11204 32784
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 11164 31822 11192 32166
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 11152 31816 11204 31822
rect 11152 31758 11204 31764
rect 10796 31482 10824 31758
rect 10784 31476 10836 31482
rect 10784 31418 10836 31424
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10690 30968 10746 30977
rect 10690 30903 10746 30912
rect 10692 30796 10744 30802
rect 10692 30738 10744 30744
rect 10704 30433 10732 30738
rect 10690 30424 10746 30433
rect 10690 30359 10746 30368
rect 10704 30054 10732 30359
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 10598 26616 10654 26625
rect 10598 26551 10654 26560
rect 10598 26480 10654 26489
rect 10598 26415 10654 26424
rect 10612 25906 10640 26415
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10612 25498 10640 25842
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10704 25378 10732 29990
rect 10784 28960 10836 28966
rect 10784 28902 10836 28908
rect 10876 28960 10928 28966
rect 10876 28902 10928 28908
rect 10796 26926 10824 28902
rect 10888 28762 10916 28902
rect 10876 28756 10928 28762
rect 10876 28698 10928 28704
rect 10888 27674 10916 28698
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 10888 27470 10916 27610
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10888 26994 10916 27406
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10784 26920 10836 26926
rect 10784 26862 10836 26868
rect 10784 26784 10836 26790
rect 10784 26726 10836 26732
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10796 25838 10824 26726
rect 10888 26586 10916 26726
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 10888 25906 10916 26386
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10784 25832 10836 25838
rect 10784 25774 10836 25780
rect 10612 25350 10732 25378
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10506 22400 10562 22409
rect 10506 22335 10562 22344
rect 10520 21570 10548 22335
rect 10612 21729 10640 25350
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10704 22137 10732 22170
rect 10796 22166 10824 22578
rect 10888 22545 10916 24618
rect 10874 22536 10930 22545
rect 10874 22471 10930 22480
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 10784 22160 10836 22166
rect 10690 22128 10746 22137
rect 10784 22102 10836 22108
rect 10690 22063 10746 22072
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10598 21720 10654 21729
rect 10704 21690 10732 21966
rect 10598 21655 10654 21664
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10520 21542 10640 21570
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 10612 21434 10640 21542
rect 10520 21146 10548 21422
rect 10612 21406 10824 21434
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10506 21040 10562 21049
rect 10506 20975 10562 20984
rect 10520 20058 10548 20975
rect 10612 20913 10640 21286
rect 10598 20904 10654 20913
rect 10598 20839 10654 20848
rect 10508 20052 10560 20058
rect 10560 20012 10640 20040
rect 10508 19994 10560 20000
rect 10506 19952 10562 19961
rect 10506 19887 10562 19896
rect 10520 19174 10548 19887
rect 10612 19242 10640 20012
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10612 18986 10640 19178
rect 10520 18958 10640 18986
rect 10704 18970 10732 19246
rect 10796 19242 10824 21406
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10692 18964 10744 18970
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10336 14482 10364 14758
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10428 14074 10456 14350
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10520 13954 10548 18958
rect 10692 18906 10744 18912
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10612 16250 10640 18770
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10704 16130 10732 18906
rect 10888 18698 10916 22374
rect 10980 21185 11008 31078
rect 11256 30734 11284 33390
rect 11244 30728 11296 30734
rect 11244 30670 11296 30676
rect 11242 29200 11298 29209
rect 11242 29135 11244 29144
rect 11296 29135 11298 29144
rect 11244 29106 11296 29112
rect 11060 28620 11112 28626
rect 11060 28562 11112 28568
rect 11072 28218 11100 28562
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 11072 27538 11100 28154
rect 11348 27946 11376 39520
rect 11808 37754 11836 39520
rect 11808 37726 12020 37754
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 11900 33454 11928 33934
rect 11888 33448 11940 33454
rect 11888 33390 11940 33396
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11428 32904 11480 32910
rect 11428 32846 11480 32852
rect 11440 31890 11468 32846
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11428 31884 11480 31890
rect 11428 31826 11480 31832
rect 11532 30870 11560 32710
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11520 30864 11572 30870
rect 11520 30806 11572 30812
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11440 30122 11468 30670
rect 11532 30394 11560 30806
rect 11520 30388 11572 30394
rect 11520 30330 11572 30336
rect 11428 30116 11480 30122
rect 11428 30058 11480 30064
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11612 29504 11664 29510
rect 11612 29446 11664 29452
rect 11624 29170 11652 29446
rect 11612 29164 11664 29170
rect 11612 29106 11664 29112
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11428 28688 11480 28694
rect 11428 28630 11480 28636
rect 11440 28218 11468 28630
rect 11428 28212 11480 28218
rect 11428 28154 11480 28160
rect 11336 27940 11388 27946
rect 11336 27882 11388 27888
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 11888 27532 11940 27538
rect 11888 27474 11940 27480
rect 11072 26194 11100 27474
rect 11334 27160 11390 27169
rect 11334 27095 11390 27104
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 11256 26518 11284 26930
rect 11348 26858 11376 27095
rect 11900 27062 11928 27474
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11992 26908 12020 37726
rect 12070 35864 12126 35873
rect 12070 35799 12126 35808
rect 12084 34746 12112 35799
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 12084 34542 12112 34682
rect 12072 34536 12124 34542
rect 12072 34478 12124 34484
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 12084 34134 12112 34342
rect 12072 34128 12124 34134
rect 12072 34070 12124 34076
rect 12084 33522 12112 34070
rect 12072 33516 12124 33522
rect 12072 33458 12124 33464
rect 12084 33046 12112 33458
rect 12072 33040 12124 33046
rect 12072 32982 12124 32988
rect 12084 32774 12112 32982
rect 12072 32768 12124 32774
rect 12072 32710 12124 32716
rect 12084 32434 12112 32710
rect 12072 32428 12124 32434
rect 12072 32370 12124 32376
rect 12084 32230 12112 32370
rect 12072 32224 12124 32230
rect 12072 32166 12124 32172
rect 12084 32026 12112 32166
rect 12072 32020 12124 32026
rect 12072 31962 12124 31968
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 11440 26880 12020 26908
rect 11336 26852 11388 26858
rect 11336 26794 11388 26800
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 11152 26240 11204 26246
rect 11072 26188 11152 26194
rect 11072 26182 11204 26188
rect 11072 26166 11192 26182
rect 11072 26042 11100 26166
rect 11256 26042 11284 26454
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 11072 24274 11100 25978
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11348 23866 11376 24210
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11058 23352 11114 23361
rect 11058 23287 11060 23296
rect 11112 23287 11114 23296
rect 11060 23258 11112 23264
rect 11348 22982 11376 23802
rect 11336 22976 11388 22982
rect 11336 22918 11388 22924
rect 11348 22778 11376 22918
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 10966 21176 11022 21185
rect 11072 21146 11100 22170
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11348 21894 11376 21966
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 10966 21111 11022 21120
rect 11060 21140 11112 21146
rect 10980 19922 11008 21111
rect 11060 21082 11112 21088
rect 11164 21010 11192 21490
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11256 19922 11284 21626
rect 11348 21554 11376 21830
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11336 21072 11388 21078
rect 11336 21014 11388 21020
rect 11348 20534 11376 21014
rect 11440 21010 11468 26880
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11532 23798 11560 26726
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11520 23792 11572 23798
rect 11520 23734 11572 23740
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11980 22976 12032 22982
rect 11980 22918 12032 22924
rect 11520 22772 11572 22778
rect 11520 22714 11572 22720
rect 11532 21690 11560 22714
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11992 22234 12020 22918
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 11886 21992 11942 22001
rect 11886 21927 11942 21936
rect 11900 21690 11928 21927
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 21146 11560 21286
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11164 19378 11192 19790
rect 11256 19514 11284 19858
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11164 18970 11192 19314
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10980 18086 11008 18702
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 17105 11008 18022
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11164 17338 11192 17818
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10966 17096 11022 17105
rect 10966 17031 11022 17040
rect 10980 16794 11008 17031
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10782 16688 10838 16697
rect 10782 16623 10784 16632
rect 10836 16623 10838 16632
rect 10784 16594 10836 16600
rect 10796 16538 10824 16594
rect 10796 16510 10916 16538
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10612 16102 10732 16130
rect 10612 14006 10640 16102
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10704 15162 10732 15914
rect 10796 15910 10824 16390
rect 10888 16114 10916 16510
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10796 14618 10824 15846
rect 10888 15706 10916 16050
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10888 14414 10916 14962
rect 10980 14804 11008 15302
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11060 14816 11112 14822
rect 10980 14776 11060 14804
rect 11060 14758 11112 14764
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10980 14362 11008 14418
rect 10980 14334 11100 14362
rect 10336 13926 10548 13954
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10336 13326 10364 13926
rect 10612 13870 10640 13942
rect 10600 13864 10652 13870
rect 10428 13812 10600 13818
rect 10428 13806 10652 13812
rect 10428 13790 10640 13806
rect 10968 13796 11020 13802
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 9876 12986 9996 13002
rect 9864 12980 9996 12986
rect 9916 12974 9996 12980
rect 9864 12922 9916 12928
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8537 9628 8774
rect 9586 8528 9642 8537
rect 9586 8463 9642 8472
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9692 7546 9720 7686
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9416 7398 9536 7426
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8864 4146 8892 5850
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 8942 5264 8998 5273
rect 8942 5199 8998 5208
rect 9312 5228 9364 5234
rect 8956 4826 8984 5199
rect 9312 5170 9364 5176
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8758 3768 8814 3777
rect 8758 3703 8814 3712
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8588 2536 8708 2564
rect 8484 2440 8536 2446
rect 8482 2408 8484 2417
rect 8536 2408 8538 2417
rect 8482 2343 8538 2352
rect 8298 2000 8354 2009
rect 8298 1935 8354 1944
rect 8588 480 8616 2536
rect 8772 2281 8800 3538
rect 8956 3534 8984 4082
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 3074 8892 3334
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8864 3046 8984 3074
rect 8956 2990 8984 3046
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8758 2272 8814 2281
rect 8758 2207 8814 2216
rect 8864 1034 8892 2858
rect 8956 2446 8984 2926
rect 9324 2632 9352 5170
rect 9416 3641 9444 7398
rect 9692 7206 9720 7482
rect 9968 7274 9996 12974
rect 10336 12442 10364 13262
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10060 8498 10088 9386
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10060 7886 10088 8434
rect 10152 8362 10180 12242
rect 10336 11801 10364 12378
rect 10428 12102 10456 13790
rect 10968 13738 11020 13744
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13530 10916 13670
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12986 10548 13194
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10520 12374 10548 12922
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10322 11792 10378 11801
rect 10322 11727 10378 11736
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 8974 10272 9318
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10138 8120 10194 8129
rect 10138 8055 10194 8064
rect 10048 7880 10100 7886
rect 10152 7868 10180 8055
rect 10244 8022 10272 8910
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10232 7880 10284 7886
rect 10152 7840 10232 7868
rect 10048 7822 10100 7828
rect 10232 7822 10284 7828
rect 10060 7410 10088 7822
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9968 6934 9996 7210
rect 10244 7206 10272 7822
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 10060 6746 10088 7142
rect 9968 6718 10088 6746
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9600 6118 9628 6258
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5914 9628 6054
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4146 9536 4966
rect 9588 4820 9640 4826
rect 9692 4808 9720 6326
rect 9772 6248 9824 6254
rect 9770 6216 9772 6225
rect 9824 6216 9826 6225
rect 9770 6151 9826 6160
rect 9640 4780 9812 4808
rect 9588 4762 9640 4768
rect 9680 4684 9732 4690
rect 9600 4644 9680 4672
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9600 3738 9628 4644
rect 9680 4626 9732 4632
rect 9784 4146 9812 4780
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9402 3632 9458 3641
rect 9402 3567 9458 3576
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 3097 9720 3334
rect 9678 3088 9734 3097
rect 9678 3023 9734 3032
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9324 2604 9444 2632
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8864 1006 8984 1034
rect 8956 480 8984 1006
rect 9416 480 9444 2604
rect 9600 2514 9628 2790
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9968 610 9996 6718
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6361 10088 6598
rect 10046 6352 10102 6361
rect 10046 6287 10102 6296
rect 10060 6254 10088 6287
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 4690 10088 5510
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9772 604 9824 610
rect 9772 546 9824 552
rect 9956 604 10008 610
rect 9956 546 10008 552
rect 9784 480 9812 546
rect 10152 480 10180 6122
rect 10244 610 10272 7142
rect 10336 5234 10364 11727
rect 10428 5914 10456 12038
rect 10520 11898 10548 12174
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10520 10130 10548 11834
rect 10704 11626 10732 12786
rect 10796 12646 10824 13330
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10980 12442 11008 13738
rect 11072 13258 11100 14334
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11058 12336 11114 12345
rect 10784 12300 10836 12306
rect 11058 12271 11114 12280
rect 10784 12242 10836 12248
rect 10796 11898 10824 12242
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10704 10248 10732 11562
rect 10612 10220 10732 10248
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10520 9722 10548 10066
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10520 9518 10548 9658
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8090 10548 8978
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10612 6440 10640 10220
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10704 9450 10732 10066
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10796 8974 10824 9658
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10704 8566 10732 8910
rect 10980 8634 11008 9114
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10888 7478 10916 7822
rect 10980 7546 11008 7822
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10520 6412 10640 6440
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10428 5370 10456 5850
rect 10520 5778 10548 6412
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10336 5137 10364 5170
rect 10322 5128 10378 5137
rect 10322 5063 10378 5072
rect 10520 4826 10548 5714
rect 10612 5710 10640 6258
rect 11072 5914 11100 12271
rect 11060 5908 11112 5914
rect 10980 5868 11060 5896
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10612 5234 10640 5646
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10980 5166 11008 5868
rect 11060 5850 11112 5856
rect 11058 5264 11114 5273
rect 11058 5199 11114 5208
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 4826 10916 4966
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11072 4706 11100 5199
rect 10888 4678 11100 4706
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4185 10456 4422
rect 10414 4176 10470 4185
rect 10414 4111 10470 4120
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10612 3942 10640 4014
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10506 3496 10562 3505
rect 10506 3431 10562 3440
rect 10520 626 10548 3431
rect 10612 2106 10640 3878
rect 10782 3768 10838 3777
rect 10782 3703 10838 3712
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10704 3233 10732 3538
rect 10796 3505 10824 3703
rect 10888 3602 10916 4678
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10980 4146 11008 4558
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10782 3496 10838 3505
rect 10782 3431 10838 3440
rect 10690 3224 10746 3233
rect 10690 3159 10692 3168
rect 10744 3159 10746 3168
rect 10692 3130 10744 3136
rect 10888 2650 10916 3538
rect 10966 2816 11022 2825
rect 10966 2751 11022 2760
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10888 2514 10916 2586
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10600 2100 10652 2106
rect 10600 2042 10652 2048
rect 10232 604 10284 610
rect 10520 598 10640 626
rect 10232 546 10284 552
rect 10612 480 10640 598
rect 10980 480 11008 2751
rect 11072 2582 11100 4014
rect 11164 3194 11192 15030
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11256 14618 11284 14894
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11348 14260 11376 20470
rect 11440 20262 11468 20946
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11808 20602 11836 20878
rect 11796 20596 11848 20602
rect 11848 20556 11928 20584
rect 11796 20538 11848 20544
rect 11900 20346 11928 20556
rect 11900 20318 12020 20346
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11440 17785 11468 20198
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11992 19990 12020 20318
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 11520 19236 11572 19242
rect 11520 19178 11572 19184
rect 11426 17776 11482 17785
rect 11426 17711 11482 17720
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11440 16998 11468 17614
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11440 16726 11468 16934
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11440 15910 11468 16662
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 14414 11468 15846
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11256 14232 11376 14260
rect 11256 13841 11284 14232
rect 11242 13832 11298 13841
rect 11242 13767 11298 13776
rect 11256 5352 11284 13767
rect 11532 13326 11560 19178
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11992 18970 12020 19926
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11980 17808 12032 17814
rect 11980 17750 12032 17756
rect 11992 17338 12020 17750
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11900 14958 11928 15302
rect 11992 15026 12020 17274
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11992 14618 12020 14962
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 13870 11836 14350
rect 11992 14074 12020 14554
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 12084 13530 12112 31758
rect 12176 23225 12204 39520
rect 12544 35290 12572 39520
rect 12532 35284 12584 35290
rect 12532 35226 12584 35232
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12268 34406 12296 34546
rect 12544 34542 12572 35226
rect 12532 34536 12584 34542
rect 12532 34478 12584 34484
rect 12256 34400 12308 34406
rect 12256 34342 12308 34348
rect 12440 34400 12492 34406
rect 12440 34342 12492 34348
rect 12452 33522 12480 34342
rect 12440 33516 12492 33522
rect 12440 33458 12492 33464
rect 12348 33380 12400 33386
rect 12348 33322 12400 33328
rect 12360 33114 12388 33322
rect 12440 33312 12492 33318
rect 12440 33254 12492 33260
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 12452 32994 12480 33254
rect 12360 32978 12480 32994
rect 12348 32972 12480 32978
rect 12400 32966 12480 32972
rect 12348 32914 12400 32920
rect 12544 32722 12572 34478
rect 12808 34400 12860 34406
rect 12808 34342 12860 34348
rect 12716 32972 12768 32978
rect 12716 32914 12768 32920
rect 12544 32694 12664 32722
rect 12636 32314 12664 32694
rect 12728 32434 12756 32914
rect 12716 32428 12768 32434
rect 12716 32370 12768 32376
rect 12636 32286 12756 32314
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 12360 30954 12388 31826
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12360 30938 12480 30954
rect 12360 30932 12492 30938
rect 12360 30926 12440 30932
rect 12360 28694 12388 30926
rect 12440 30874 12492 30880
rect 12636 28948 12664 31282
rect 12544 28920 12664 28948
rect 12348 28688 12400 28694
rect 12348 28630 12400 28636
rect 12348 27600 12400 27606
rect 12348 27542 12400 27548
rect 12254 26888 12310 26897
rect 12254 26823 12256 26832
rect 12308 26823 12310 26832
rect 12256 26794 12308 26800
rect 12360 26586 12388 27542
rect 12440 26784 12492 26790
rect 12440 26726 12492 26732
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12360 26450 12388 26522
rect 12452 26489 12480 26726
rect 12438 26480 12494 26489
rect 12348 26444 12400 26450
rect 12438 26415 12494 26424
rect 12348 26386 12400 26392
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12360 23526 12388 24210
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12162 23216 12218 23225
rect 12162 23151 12218 23160
rect 12360 23050 12388 23462
rect 12452 23186 12480 24006
rect 12544 23322 12572 28920
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12348 23044 12400 23050
rect 12348 22986 12400 22992
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 12176 15162 12204 22442
rect 12268 15502 12296 22714
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12360 22098 12388 22374
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 12452 22030 12480 23122
rect 12544 22778 12572 23258
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12438 20904 12494 20913
rect 12438 20839 12494 20848
rect 12452 20602 12480 20839
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12256 15496 12308 15502
rect 12254 15464 12256 15473
rect 12308 15464 12310 15473
rect 12254 15399 12310 15408
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12176 14958 12204 15098
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12176 14278 12204 14486
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12360 13802 12388 15574
rect 12728 15162 12756 32286
rect 12820 26976 12848 34342
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 12912 32570 12940 33050
rect 12900 32564 12952 32570
rect 12900 32506 12952 32512
rect 12912 31346 12940 32506
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 13004 27169 13032 39520
rect 13188 39494 13400 39520
rect 13084 33856 13136 33862
rect 13084 33798 13136 33804
rect 13096 33522 13124 33798
rect 13084 33516 13136 33522
rect 13084 33458 13136 33464
rect 12990 27160 13046 27169
rect 12990 27095 13046 27104
rect 13188 27033 13216 39494
rect 13740 35714 13768 39520
rect 13648 35686 13768 35714
rect 13832 39494 14228 39520
rect 13544 31272 13596 31278
rect 13544 31214 13596 31220
rect 13452 27328 13504 27334
rect 13452 27270 13504 27276
rect 13174 27024 13230 27033
rect 12992 26988 13044 26994
rect 12820 26948 12940 26976
rect 12806 26888 12862 26897
rect 12806 26823 12808 26832
rect 12860 26823 12862 26832
rect 12808 26794 12860 26800
rect 12808 23180 12860 23186
rect 12808 23122 12860 23128
rect 12820 22574 12848 23122
rect 12912 22642 12940 26948
rect 12992 26930 13044 26936
rect 13096 26982 13174 27010
rect 13004 26518 13032 26930
rect 12992 26512 13044 26518
rect 12992 26454 13044 26460
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12820 22234 12848 22510
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 13004 21554 13032 22578
rect 13096 22506 13124 26982
rect 13174 26959 13230 26968
rect 13266 25256 13322 25265
rect 13266 25191 13322 25200
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13188 22642 13216 22918
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13084 22500 13136 22506
rect 13084 22442 13136 22448
rect 13096 21894 13124 22442
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13004 21146 13032 21490
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13004 20466 13032 21082
rect 13096 21010 13124 21830
rect 13280 21128 13308 25191
rect 13464 24993 13492 27270
rect 13450 24984 13506 24993
rect 13450 24919 13506 24928
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13188 21100 13308 21128
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 13188 20890 13216 21100
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13096 20862 13216 20890
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12898 20360 12954 20369
rect 12898 20295 12900 20304
rect 12952 20295 12954 20304
rect 12900 20266 12952 20272
rect 13004 20058 13032 20402
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 12912 15162 12940 15370
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 14278 12480 14962
rect 12728 14822 12756 15098
rect 13004 15026 13032 15302
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 13096 14362 13124 20862
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 13188 20398 13216 20742
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13188 19961 13216 20334
rect 13174 19952 13230 19961
rect 13174 19887 13230 19896
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 16697 13216 17478
rect 13174 16688 13230 16697
rect 13174 16623 13230 16632
rect 12544 14334 13124 14362
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 14074 12480 14214
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11256 5324 11468 5352
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11348 4758 11376 5170
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11150 2952 11206 2961
rect 11150 2887 11206 2896
rect 11164 2854 11192 2887
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11256 2689 11284 4490
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11348 3942 11376 4082
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3670 11376 3878
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11348 3398 11376 3606
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11334 3088 11390 3097
rect 11334 3023 11390 3032
rect 11242 2680 11298 2689
rect 11242 2615 11298 2624
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11256 2281 11284 2615
rect 11242 2272 11298 2281
rect 11242 2207 11298 2216
rect 11348 480 11376 3023
rect 11440 2666 11468 5324
rect 11532 4214 11560 12922
rect 11900 12850 11928 13262
rect 12084 12986 12112 13466
rect 12452 13326 12480 14010
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12452 12986 12480 13262
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 12084 12345 12112 12582
rect 12452 12442 12480 12922
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12070 12336 12126 12345
rect 12070 12271 12126 12280
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 12544 11098 12572 14334
rect 13280 14226 13308 20946
rect 13096 14198 13308 14226
rect 12544 11070 12756 11098
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12346 10704 12402 10713
rect 12544 10674 12572 10950
rect 12346 10639 12402 10648
rect 12532 10668 12584 10674
rect 12254 10568 12310 10577
rect 12254 10503 12256 10512
rect 12308 10503 12310 10512
rect 12256 10474 12308 10480
rect 12254 10432 12310 10441
rect 11622 10364 11918 10384
rect 12254 10367 12310 10376
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 12070 10024 12126 10033
rect 12070 9959 12126 9968
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9586 12020 9862
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11992 9110 12020 9522
rect 11980 9104 12032 9110
rect 11900 9052 11980 9058
rect 11900 9046 12032 9052
rect 11900 9030 12020 9046
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 8634 11744 8910
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11716 8378 11744 8570
rect 11900 8566 11928 9030
rect 11978 8936 12034 8945
rect 11978 8871 12034 8880
rect 11992 8634 12020 8871
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11716 8350 12020 8378
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11992 6905 12020 8350
rect 11978 6896 12034 6905
rect 11978 6831 11980 6840
rect 12032 6831 12034 6840
rect 11980 6802 12032 6808
rect 11992 6458 12020 6802
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11992 5914 12020 6394
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11624 5370 11652 5714
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11624 5273 11652 5306
rect 11610 5264 11666 5273
rect 11900 5234 11928 5714
rect 11610 5199 11666 5208
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 12084 3194 12112 9959
rect 12268 6769 12296 10367
rect 12360 10033 12388 10639
rect 12532 10610 12584 10616
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12346 10024 12402 10033
rect 12346 9959 12402 9968
rect 12544 9654 12572 10406
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12452 8430 12480 9454
rect 12544 9382 12572 9590
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12452 8090 12480 8366
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12636 6866 12664 9114
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12254 6760 12310 6769
rect 12254 6695 12310 6704
rect 12636 6458 12664 6802
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 4826 12664 4966
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12360 3738 12388 4150
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12452 3466 12480 4626
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12544 4214 12572 4558
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12084 2854 12112 3130
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11440 2638 11560 2666
rect 12452 2650 12480 3402
rect 11532 2632 11560 2638
rect 12440 2644 12492 2650
rect 11532 2604 11836 2632
rect 11808 480 11836 2604
rect 12440 2586 12492 2592
rect 12544 2553 12572 3878
rect 12636 3194 12664 4762
rect 12728 3210 12756 11070
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 10266 12940 10406
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12912 10033 12940 10202
rect 12898 10024 12954 10033
rect 12898 9959 12954 9968
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12820 8634 12848 9454
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13004 8498 13032 10610
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8090 13032 8434
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4078 12848 4422
rect 12898 4176 12954 4185
rect 12898 4111 12900 4120
rect 12952 4111 12954 4120
rect 12900 4082 12952 4088
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13004 3738 13032 5510
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13004 3398 13032 3674
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12806 3224 12862 3233
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12728 3182 12806 3210
rect 12728 2582 12756 3182
rect 12806 3159 12862 3168
rect 13004 3058 13032 3334
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12808 2848 12860 2854
rect 12806 2816 12808 2825
rect 12900 2848 12952 2854
rect 12860 2816 12862 2825
rect 12900 2790 12952 2796
rect 12806 2751 12862 2760
rect 12716 2576 12768 2582
rect 12530 2544 12586 2553
rect 12716 2518 12768 2524
rect 12530 2479 12586 2488
rect 12912 2417 12940 2790
rect 12898 2408 12954 2417
rect 12898 2343 12954 2352
rect 12532 2100 12584 2106
rect 12532 2042 12584 2048
rect 12164 604 12216 610
rect 12164 546 12216 552
rect 12176 480 12204 546
rect 12544 480 12572 2042
rect 12990 2000 13046 2009
rect 12990 1935 13046 1944
rect 13004 480 13032 1935
rect 13096 1737 13124 14198
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9722 13308 10066
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13280 9586 13308 9658
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13280 2446 13308 2994
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13082 1728 13138 1737
rect 13082 1663 13138 1672
rect 13372 480 13400 21286
rect 13464 20097 13492 24919
rect 13450 20088 13506 20097
rect 13450 20023 13506 20032
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13464 9382 13492 9998
rect 13556 9994 13584 31214
rect 13648 30433 13676 35686
rect 13726 33416 13782 33425
rect 13726 33351 13782 33360
rect 13740 31482 13768 33351
rect 13728 31476 13780 31482
rect 13728 31418 13780 31424
rect 13634 30424 13690 30433
rect 13634 30359 13690 30368
rect 13832 24857 13860 39494
rect 14568 37210 14596 39520
rect 14936 39494 15056 39520
rect 14568 37182 14688 37210
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14660 31385 14688 37182
rect 14646 31376 14702 31385
rect 14646 31311 14702 31320
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 15028 25265 15056 39494
rect 15396 31249 15424 39520
rect 15764 33114 15792 39520
rect 15752 33108 15804 33114
rect 15752 33050 15804 33056
rect 15382 31240 15438 31249
rect 15382 31175 15438 31184
rect 15014 25256 15070 25265
rect 15014 25191 15070 25200
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 13818 24848 13874 24857
rect 13818 24783 13874 24792
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14770 13768 14826
rect 13740 14742 13860 14770
rect 13726 10160 13782 10169
rect 13636 10124 13688 10130
rect 13726 10095 13782 10104
rect 13636 10066 13688 10072
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 9178 13492 9318
rect 13648 9178 13676 10066
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13648 8906 13676 9114
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 5846 13492 6598
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13464 2650 13492 3470
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13740 480 13768 10095
rect 13832 7546 13860 14742
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14002 3496 14058 3505
rect 14002 3431 14058 3440
rect 14016 1850 14044 3431
rect 14108 2394 14136 10474
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 15382 3632 15438 3641
rect 15382 3567 15438 3576
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14922 2816 14978 2825
rect 14922 2751 14978 2760
rect 14108 2366 14228 2394
rect 14096 2304 14148 2310
rect 14094 2272 14096 2281
rect 14148 2272 14150 2281
rect 14094 2207 14150 2216
rect 14200 1986 14228 2366
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14200 1958 14596 1986
rect 14016 1822 14228 1850
rect 14200 480 14228 1822
rect 14568 480 14596 1958
rect 14936 480 14964 2751
rect 15396 480 15424 3567
rect 15764 480 15792 7482
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 1582 38664 1638 38720
rect 1490 36352 1546 36408
rect 570 33904 626 33960
rect 1766 35128 1822 35184
rect 1582 34040 1638 34096
rect 1674 32444 1676 32464
rect 1676 32444 1728 32464
rect 1728 32444 1730 32464
rect 1674 32408 1730 32444
rect 1582 31592 1638 31648
rect 1582 29300 1638 29336
rect 1582 29280 1584 29300
rect 1584 29280 1636 29300
rect 1636 29280 1638 29300
rect 1766 29008 1822 29064
rect 1582 26968 1638 27024
rect 2594 35264 2650 35320
rect 1950 33396 1952 33416
rect 1952 33396 2004 33416
rect 2004 33396 2006 33416
rect 1950 33360 2006 33396
rect 1858 25880 1914 25936
rect 1582 24520 1638 24576
rect 1674 22652 1676 22672
rect 1676 22652 1728 22672
rect 1728 22652 1730 22672
rect 1674 22616 1730 22652
rect 1582 21956 1638 21992
rect 1582 21936 1584 21956
rect 1584 21936 1636 21956
rect 1636 21936 1638 21956
rect 1674 20884 1676 20904
rect 1676 20884 1728 20904
rect 1728 20884 1730 20904
rect 1674 20848 1730 20884
rect 1582 19896 1638 19952
rect 1950 18284 2006 18320
rect 1950 18264 1952 18284
rect 1952 18264 2004 18284
rect 2004 18264 2006 18284
rect 1582 17584 1638 17640
rect 1950 16108 2006 16144
rect 1950 16088 1952 16108
rect 1952 16088 2004 16108
rect 2004 16088 2006 16108
rect 1582 15136 1638 15192
rect 2318 33516 2374 33552
rect 2318 33496 2320 33516
rect 2320 33496 2372 33516
rect 2372 33496 2374 33516
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 2502 29688 2558 29744
rect 2870 29008 2926 29064
rect 3146 30640 3202 30696
rect 2962 28056 3018 28112
rect 2778 27376 2834 27432
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 4526 35672 4582 35728
rect 4250 33924 4306 33960
rect 4250 33904 4252 33924
rect 4252 33904 4304 33924
rect 4304 33904 4306 33924
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 4710 35284 4766 35320
rect 4710 35264 4712 35284
rect 4712 35264 4764 35284
rect 4764 35264 4766 35284
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 2778 22480 2834 22536
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 2134 14864 2190 14920
rect 1674 12436 1730 12472
rect 1674 12416 1676 12436
rect 1676 12416 1728 12436
rect 1728 12416 1730 12436
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 2778 12824 2834 12880
rect 1582 10512 1638 10568
rect 1950 7148 1952 7168
rect 1952 7148 2004 7168
rect 2004 7148 2006 7168
rect 570 4256 626 4312
rect 1398 4564 1400 4584
rect 1400 4564 1452 4584
rect 1452 4564 1454 4584
rect 1398 4528 1454 4564
rect 1950 7112 2006 7148
rect 1582 5752 1638 5808
rect 1766 4664 1822 4720
rect 1490 3440 1546 3496
rect 2778 8472 2834 8528
rect 2778 8064 2834 8120
rect 3054 7248 3110 7304
rect 2870 6840 2926 6896
rect 2318 4120 2374 4176
rect 2318 3440 2374 3496
rect 1950 2760 2006 2816
rect 1858 1128 1914 1184
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3330 9444 3386 9480
rect 3330 9424 3332 9444
rect 3332 9424 3384 9444
rect 3384 9424 3386 9444
rect 3054 4256 3110 4312
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3790 8336 3846 8392
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 4066 6840 4122 6896
rect 2502 2488 2558 2544
rect 2410 1672 2466 1728
rect 4986 31320 5042 31376
rect 4986 28212 5042 28248
rect 4986 28192 4988 28212
rect 4988 28192 5040 28212
rect 5040 28192 5042 28212
rect 5814 32308 5816 32328
rect 5816 32308 5868 32328
rect 5868 32308 5870 32328
rect 5814 32272 5870 32308
rect 5630 31864 5686 31920
rect 5630 31320 5686 31376
rect 5078 24812 5134 24848
rect 5078 24792 5080 24812
rect 5080 24792 5132 24812
rect 5132 24792 5134 24812
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6182 30676 6184 30696
rect 6184 30676 6236 30696
rect 6236 30676 6238 30696
rect 6182 30640 6238 30676
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 5722 28192 5778 28248
rect 5814 27940 5870 27976
rect 5814 27920 5816 27940
rect 5816 27920 5868 27940
rect 5868 27920 5870 27940
rect 6366 28328 6422 28384
rect 7746 36352 7802 36408
rect 7562 35128 7618 35184
rect 6826 30932 6882 30968
rect 6826 30912 6828 30932
rect 6828 30912 6880 30932
rect 6880 30912 6882 30932
rect 6734 27920 6790 27976
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 7010 26832 7066 26888
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 5722 22616 5778 22672
rect 4894 21528 4950 21584
rect 5538 21392 5594 21448
rect 5538 17720 5594 17776
rect 5906 20984 5962 21040
rect 4710 15952 4766 16008
rect 4618 14884 4674 14920
rect 4618 14864 4620 14884
rect 4620 14864 4672 14884
rect 4672 14864 4674 14884
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3606 3732 3662 3768
rect 3606 3712 3608 3732
rect 3608 3712 3660 3732
rect 3660 3712 3662 3732
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3054 3032 3110 3088
rect 2778 2372 2834 2408
rect 2778 2352 2780 2372
rect 2780 2352 2832 2372
rect 2832 2352 2834 2372
rect 4986 13812 4988 13832
rect 4988 13812 5040 13832
rect 5040 13812 5042 13832
rect 4986 13776 5042 13812
rect 5354 15000 5410 15056
rect 5446 12688 5502 12744
rect 5170 12416 5226 12472
rect 5354 12300 5410 12336
rect 5354 12280 5356 12300
rect 5356 12280 5408 12300
rect 5408 12280 5410 12300
rect 4618 6160 4674 6216
rect 5446 11736 5502 11792
rect 5814 12688 5870 12744
rect 5630 8880 5686 8936
rect 5538 7112 5594 7168
rect 4802 4120 4858 4176
rect 4526 2896 4582 2952
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 4158 1400 4214 1456
rect 5446 5652 5448 5672
rect 5448 5652 5500 5672
rect 5500 5652 5502 5672
rect 5446 5616 5502 5652
rect 5262 3576 5318 3632
rect 6090 24792 6146 24848
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 7746 33904 7802 33960
rect 7562 33360 7618 33416
rect 7470 32988 7472 33008
rect 7472 32988 7524 33008
rect 7524 32988 7526 33008
rect 7470 32952 7526 32988
rect 7470 32444 7472 32464
rect 7472 32444 7524 32464
rect 7524 32444 7526 32464
rect 7470 32408 7526 32444
rect 7378 27512 7434 27568
rect 7470 27376 7526 27432
rect 7286 26988 7342 27024
rect 7746 29028 7802 29064
rect 7746 29008 7748 29028
rect 7748 29008 7800 29028
rect 7800 29008 7802 29028
rect 7746 28056 7802 28112
rect 7286 26968 7288 26988
rect 7288 26968 7340 26988
rect 7340 26968 7342 26988
rect 7286 25200 7342 25256
rect 7102 23024 7158 23080
rect 7470 23160 7526 23216
rect 8390 32408 8446 32464
rect 7746 21256 7802 21312
rect 6550 14456 6606 14512
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6458 10532 6514 10568
rect 6458 10512 6460 10532
rect 6460 10512 6512 10532
rect 6512 10512 6514 10532
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 7838 18264 7894 18320
rect 5538 3712 5594 3768
rect 5354 2760 5410 2816
rect 5262 2252 5264 2272
rect 5264 2252 5316 2272
rect 5316 2252 5318 2272
rect 5262 2216 5318 2252
rect 5630 3440 5686 3496
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6826 5616 6882 5672
rect 7654 17856 7710 17912
rect 7654 15952 7710 16008
rect 7562 15564 7618 15600
rect 7562 15544 7564 15564
rect 7564 15544 7616 15564
rect 7616 15544 7618 15564
rect 7102 8064 7158 8120
rect 7102 6704 7158 6760
rect 7378 7928 7434 7984
rect 7654 8472 7710 8528
rect 6182 4528 6238 4584
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6642 3032 6698 3088
rect 6918 3032 6974 3088
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 6734 2760 6790 2816
rect 7286 4140 7342 4176
rect 7286 4120 7288 4140
rect 7288 4120 7340 4140
rect 7340 4120 7342 4140
rect 7102 3440 7158 3496
rect 7286 3712 7342 3768
rect 7102 1400 7158 1456
rect 8298 29008 8354 29064
rect 8390 28328 8446 28384
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 9678 35808 9734 35864
rect 9402 32952 9458 33008
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 9310 31184 9366 31240
rect 8666 30776 8722 30832
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8574 27820 8576 27840
rect 8576 27820 8628 27840
rect 8628 27820 8630 27840
rect 8574 27784 8630 27820
rect 8206 21936 8262 21992
rect 7930 15272 7986 15328
rect 8114 10648 8170 10704
rect 8114 10260 8170 10296
rect 8114 10240 8116 10260
rect 8116 10240 8168 10260
rect 8168 10240 8170 10260
rect 7930 9424 7986 9480
rect 8574 25916 8576 25936
rect 8576 25916 8628 25936
rect 8628 25916 8630 25936
rect 8574 25880 8630 25916
rect 8850 29688 8906 29744
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 9862 36372 9918 36408
rect 9862 36352 9864 36372
rect 9864 36352 9916 36372
rect 9916 36352 9918 36372
rect 9862 35708 9864 35728
rect 9864 35708 9916 35728
rect 9916 35708 9918 35728
rect 9862 35672 9918 35708
rect 9954 33904 10010 33960
rect 10138 33396 10140 33416
rect 10140 33396 10192 33416
rect 10192 33396 10194 33416
rect 10138 33360 10194 33396
rect 9310 27648 9366 27704
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 9586 29144 9642 29200
rect 9586 28056 9642 28112
rect 9678 27784 9734 27840
rect 9678 27376 9734 27432
rect 8390 16632 8446 16688
rect 8482 12688 8538 12744
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 9402 24928 9458 24984
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8666 20712 8722 20768
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 9402 23296 9458 23352
rect 9678 23024 9734 23080
rect 10046 30796 10102 30832
rect 10046 30776 10048 30796
rect 10048 30776 10100 30796
rect 10100 30776 10102 30796
rect 10046 27532 10102 27568
rect 10046 27512 10048 27532
rect 10048 27512 10100 27532
rect 10100 27512 10102 27532
rect 9770 22344 9826 22400
rect 9402 22072 9458 22128
rect 9586 22072 9642 22128
rect 9770 22072 9826 22128
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 9678 21800 9734 21856
rect 9862 21800 9918 21856
rect 9862 21664 9918 21720
rect 9586 21392 9642 21448
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 9770 21528 9826 21584
rect 9678 20848 9734 20904
rect 9862 17856 9918 17912
rect 9494 17076 9496 17096
rect 9496 17076 9548 17096
rect 9548 17076 9550 17096
rect 9494 17040 9550 17076
rect 8666 9968 8722 10024
rect 8114 8472 8170 8528
rect 7930 7928 7986 7984
rect 7746 5228 7802 5264
rect 7746 5208 7748 5228
rect 7748 5208 7800 5228
rect 7800 5208 7802 5228
rect 8390 7948 8446 7984
rect 8390 7928 8392 7948
rect 8392 7928 8444 7948
rect 8444 7928 8446 7948
rect 8298 6296 8354 6352
rect 8206 5344 8262 5400
rect 8206 5208 8262 5264
rect 8390 4664 8446 4720
rect 7562 2760 7618 2816
rect 7930 2760 7986 2816
rect 8114 2488 8170 2544
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8758 7284 8760 7304
rect 8760 7284 8812 7304
rect 8812 7284 8814 7304
rect 8758 7248 8814 7284
rect 9310 8356 9366 8392
rect 9310 8336 9312 8356
rect 9312 8336 9364 8356
rect 9364 8336 9366 8356
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8850 6840 8906 6896
rect 8666 5072 8722 5128
rect 8482 2644 8538 2680
rect 8482 2624 8484 2644
rect 8484 2624 8536 2644
rect 8536 2624 8538 2644
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 9586 12688 9642 12744
rect 9494 12416 9550 12472
rect 9494 10240 9550 10296
rect 10230 23296 10286 23352
rect 10506 32408 10562 32464
rect 10414 31864 10470 31920
rect 10414 29028 10470 29064
rect 10414 29008 10416 29028
rect 10416 29008 10468 29028
rect 10468 29008 10470 29028
rect 10506 27784 10562 27840
rect 10138 21800 10194 21856
rect 10046 20304 10102 20360
rect 10138 19080 10194 19136
rect 10230 18944 10286 19000
rect 10230 16632 10286 16688
rect 10322 16124 10324 16144
rect 10324 16124 10376 16144
rect 10376 16124 10378 16144
rect 10322 16088 10378 16124
rect 10782 33496 10838 33552
rect 10690 30912 10746 30968
rect 10690 30368 10746 30424
rect 10598 26560 10654 26616
rect 10598 26424 10654 26480
rect 10506 22344 10562 22400
rect 10874 22480 10930 22536
rect 10690 22072 10746 22128
rect 10598 21664 10654 21720
rect 10506 20984 10562 21040
rect 10598 20848 10654 20904
rect 10506 19896 10562 19952
rect 11242 29164 11298 29200
rect 11242 29144 11244 29164
rect 11244 29144 11296 29164
rect 11296 29144 11298 29164
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11334 27104 11390 27160
rect 12070 35808 12126 35864
rect 11058 23316 11114 23352
rect 11058 23296 11060 23316
rect 11060 23296 11112 23316
rect 11112 23296 11114 23316
rect 10966 21120 11022 21176
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11886 21936 11942 21992
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 10966 17040 11022 17096
rect 10782 16652 10838 16688
rect 10782 16632 10784 16652
rect 10784 16632 10836 16652
rect 10836 16632 10838 16652
rect 9586 8472 9642 8528
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8942 5208 8998 5264
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8758 3712 8814 3768
rect 8482 2388 8484 2408
rect 8484 2388 8536 2408
rect 8536 2388 8538 2408
rect 8482 2352 8538 2388
rect 8298 1944 8354 2000
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8758 2216 8814 2272
rect 10322 11736 10378 11792
rect 10138 8064 10194 8120
rect 9770 6196 9772 6216
rect 9772 6196 9824 6216
rect 9824 6196 9826 6216
rect 9770 6160 9826 6196
rect 9402 3576 9458 3632
rect 9678 3032 9734 3088
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 10046 6296 10102 6352
rect 11058 12280 11114 12336
rect 10322 5072 10378 5128
rect 11058 5208 11114 5264
rect 10414 4120 10470 4176
rect 10506 3440 10562 3496
rect 10782 3712 10838 3768
rect 10782 3440 10838 3496
rect 10690 3188 10746 3224
rect 10690 3168 10692 3188
rect 10692 3168 10744 3188
rect 10744 3168 10746 3188
rect 10966 2760 11022 2816
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11426 17720 11482 17776
rect 11242 13776 11298 13832
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 12254 26852 12310 26888
rect 12254 26832 12256 26852
rect 12256 26832 12308 26852
rect 12308 26832 12310 26852
rect 12438 26424 12494 26480
rect 12162 23160 12218 23216
rect 12438 20848 12494 20904
rect 12254 15444 12256 15464
rect 12256 15444 12308 15464
rect 12308 15444 12310 15464
rect 12254 15408 12310 15444
rect 12990 27104 13046 27160
rect 12806 26852 12862 26888
rect 12806 26832 12808 26852
rect 12808 26832 12860 26852
rect 12860 26832 12862 26852
rect 13174 26968 13230 27024
rect 13266 25200 13322 25256
rect 13450 24928 13506 24984
rect 12898 20324 12954 20360
rect 12898 20304 12900 20324
rect 12900 20304 12952 20324
rect 12952 20304 12954 20324
rect 13174 19896 13230 19952
rect 13174 16632 13230 16688
rect 11150 2896 11206 2952
rect 11334 3032 11390 3088
rect 11242 2624 11298 2680
rect 11242 2216 11298 2272
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 12070 12280 12126 12336
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 12346 10648 12402 10704
rect 12254 10532 12310 10568
rect 12254 10512 12256 10532
rect 12256 10512 12308 10532
rect 12308 10512 12310 10532
rect 12254 10376 12310 10432
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 12070 9968 12126 10024
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11978 8880 12034 8936
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11978 6860 12034 6896
rect 11978 6840 11980 6860
rect 11980 6840 12032 6860
rect 12032 6840 12034 6860
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11610 5208 11666 5264
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 12346 9968 12402 10024
rect 12254 6704 12310 6760
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12898 9968 12954 10024
rect 12898 4140 12954 4176
rect 12898 4120 12900 4140
rect 12900 4120 12952 4140
rect 12952 4120 12954 4140
rect 12806 3168 12862 3224
rect 12806 2796 12808 2816
rect 12808 2796 12860 2816
rect 12860 2796 12862 2816
rect 12806 2760 12862 2796
rect 12530 2488 12586 2544
rect 12898 2352 12954 2408
rect 12990 1944 13046 2000
rect 13082 1672 13138 1728
rect 13450 20032 13506 20088
rect 13726 33360 13782 33416
rect 13634 30368 13690 30424
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14646 31320 14702 31376
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 15382 31184 15438 31240
rect 15014 25200 15070 25256
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 13818 24792 13874 24848
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 13726 10104 13782 10160
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14002 3440 14058 3496
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 15382 3576 15438 3632
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14922 2760 14978 2816
rect 14094 2252 14096 2272
rect 14096 2252 14148 2272
rect 14148 2252 14150 2272
rect 14094 2216 14150 2252
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 0 38722 480 38752
rect 1577 38722 1643 38725
rect 0 38720 1643 38722
rect 0 38664 1582 38720
rect 1638 38664 1643 38720
rect 0 38662 1643 38664
rect 0 38632 480 38662
rect 1577 38659 1643 38662
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 0 36410 480 36440
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 1485 36410 1551 36413
rect 0 36408 1551 36410
rect 0 36352 1490 36408
rect 1546 36352 1551 36408
rect 0 36350 1551 36352
rect 0 36320 480 36350
rect 1485 36347 1551 36350
rect 7741 36410 7807 36413
rect 9857 36410 9923 36413
rect 7741 36408 9923 36410
rect 7741 36352 7746 36408
rect 7802 36352 9862 36408
rect 9918 36352 9923 36408
rect 7741 36350 9923 36352
rect 7741 36347 7807 36350
rect 9857 36347 9923 36350
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 9673 35866 9739 35869
rect 12065 35866 12131 35869
rect 9673 35864 12131 35866
rect 9673 35808 9678 35864
rect 9734 35808 12070 35864
rect 12126 35808 12131 35864
rect 9673 35806 12131 35808
rect 9673 35803 9739 35806
rect 12065 35803 12131 35806
rect 4521 35730 4587 35733
rect 9857 35730 9923 35733
rect 4521 35728 9923 35730
rect 4521 35672 4526 35728
rect 4582 35672 9862 35728
rect 9918 35672 9923 35728
rect 4521 35670 9923 35672
rect 4521 35667 4587 35670
rect 9857 35667 9923 35670
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 2589 35322 2655 35325
rect 4705 35322 4771 35325
rect 2589 35320 4771 35322
rect 2589 35264 2594 35320
rect 2650 35264 4710 35320
rect 4766 35264 4771 35320
rect 2589 35262 4771 35264
rect 2589 35259 2655 35262
rect 4705 35259 4771 35262
rect 1761 35186 1827 35189
rect 7557 35186 7623 35189
rect 1761 35184 7623 35186
rect 1761 35128 1766 35184
rect 1822 35128 7562 35184
rect 7618 35128 7623 35184
rect 1761 35126 7623 35128
rect 1761 35123 1827 35126
rect 7557 35123 7623 35126
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 0 34098 480 34128
rect 1577 34098 1643 34101
rect 0 34096 1643 34098
rect 0 34040 1582 34096
rect 1638 34040 1643 34096
rect 0 34038 1643 34040
rect 0 34008 480 34038
rect 1577 34035 1643 34038
rect 565 33962 631 33965
rect 4245 33962 4311 33965
rect 565 33960 4311 33962
rect 565 33904 570 33960
rect 626 33904 4250 33960
rect 4306 33904 4311 33960
rect 565 33902 4311 33904
rect 565 33899 631 33902
rect 4245 33899 4311 33902
rect 7741 33962 7807 33965
rect 9949 33962 10015 33965
rect 7741 33960 10015 33962
rect 7741 33904 7746 33960
rect 7802 33904 9954 33960
rect 10010 33904 10015 33960
rect 7741 33902 10015 33904
rect 7741 33899 7807 33902
rect 9949 33899 10015 33902
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 2313 33554 2379 33557
rect 10777 33554 10843 33557
rect 2313 33552 10843 33554
rect 2313 33496 2318 33552
rect 2374 33496 10782 33552
rect 10838 33496 10843 33552
rect 2313 33494 10843 33496
rect 2313 33491 2379 33494
rect 10777 33491 10843 33494
rect 1945 33418 2011 33421
rect 7557 33418 7623 33421
rect 10133 33418 10199 33421
rect 1945 33416 10199 33418
rect 1945 33360 1950 33416
rect 2006 33360 7562 33416
rect 7618 33360 10138 33416
rect 10194 33360 10199 33416
rect 1945 33358 10199 33360
rect 1945 33355 2011 33358
rect 7557 33355 7623 33358
rect 10133 33355 10199 33358
rect 13721 33418 13787 33421
rect 15520 33418 16000 33448
rect 13721 33416 16000 33418
rect 13721 33360 13726 33416
rect 13782 33360 16000 33416
rect 13721 33358 16000 33360
rect 13721 33355 13787 33358
rect 15520 33328 16000 33358
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 7465 33010 7531 33013
rect 9397 33010 9463 33013
rect 7465 33008 9463 33010
rect 7465 32952 7470 33008
rect 7526 32952 9402 33008
rect 9458 32952 9463 33008
rect 7465 32950 9463 32952
rect 7465 32947 7531 32950
rect 9397 32947 9463 32950
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 1669 32466 1735 32469
rect 7465 32466 7531 32469
rect 8385 32466 8451 32469
rect 10501 32466 10567 32469
rect 1669 32464 7531 32466
rect 1669 32408 1674 32464
rect 1730 32408 7470 32464
rect 7526 32408 7531 32464
rect 1669 32406 7531 32408
rect 1669 32403 1735 32406
rect 7465 32403 7531 32406
rect 7974 32464 10567 32466
rect 7974 32408 8390 32464
rect 8446 32408 10506 32464
rect 10562 32408 10567 32464
rect 7974 32406 10567 32408
rect 5809 32330 5875 32333
rect 7974 32330 8034 32406
rect 8385 32403 8451 32406
rect 10501 32403 10567 32406
rect 5809 32328 8034 32330
rect 5809 32272 5814 32328
rect 5870 32272 8034 32328
rect 5809 32270 8034 32272
rect 5809 32267 5875 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 5625 31922 5691 31925
rect 10409 31922 10475 31925
rect 5625 31920 10475 31922
rect 5625 31864 5630 31920
rect 5686 31864 10414 31920
rect 10470 31864 10475 31920
rect 5625 31862 10475 31864
rect 5625 31859 5691 31862
rect 10409 31859 10475 31862
rect 0 31650 480 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 480 31590
rect 1577 31587 1643 31590
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 4981 31378 5047 31381
rect 5625 31378 5691 31381
rect 14641 31378 14707 31381
rect 4981 31376 14707 31378
rect 4981 31320 4986 31376
rect 5042 31320 5630 31376
rect 5686 31320 14646 31376
rect 14702 31320 14707 31376
rect 4981 31318 14707 31320
rect 4981 31315 5047 31318
rect 5625 31315 5691 31318
rect 14641 31315 14707 31318
rect 9305 31242 9371 31245
rect 15377 31242 15443 31245
rect 9305 31240 15443 31242
rect 9305 31184 9310 31240
rect 9366 31184 15382 31240
rect 15438 31184 15443 31240
rect 9305 31182 15443 31184
rect 9305 31179 9371 31182
rect 15377 31179 15443 31182
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 6821 30970 6887 30973
rect 10685 30970 10751 30973
rect 6821 30968 10751 30970
rect 6821 30912 6826 30968
rect 6882 30912 10690 30968
rect 10746 30912 10751 30968
rect 6821 30910 10751 30912
rect 6821 30907 6887 30910
rect 10685 30907 10751 30910
rect 8661 30834 8727 30837
rect 10041 30834 10107 30837
rect 8661 30832 10107 30834
rect 8661 30776 8666 30832
rect 8722 30776 10046 30832
rect 10102 30776 10107 30832
rect 8661 30774 10107 30776
rect 8661 30771 8727 30774
rect 10041 30771 10107 30774
rect 3141 30698 3207 30701
rect 6177 30698 6243 30701
rect 3141 30696 6243 30698
rect 3141 30640 3146 30696
rect 3202 30640 6182 30696
rect 6238 30640 6243 30696
rect 3141 30638 6243 30640
rect 3141 30635 3207 30638
rect 6177 30635 6243 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 10685 30426 10751 30429
rect 13629 30426 13695 30429
rect 10685 30424 13695 30426
rect 10685 30368 10690 30424
rect 10746 30368 13634 30424
rect 13690 30368 13695 30424
rect 10685 30366 13695 30368
rect 10685 30363 10751 30366
rect 13629 30363 13695 30366
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 2497 29746 2563 29749
rect 8845 29746 8911 29749
rect 2497 29744 8911 29746
rect 2497 29688 2502 29744
rect 2558 29688 8850 29744
rect 8906 29688 8911 29744
rect 2497 29686 8911 29688
rect 2497 29683 2563 29686
rect 8845 29683 8911 29686
rect 3610 29408 3930 29409
rect 0 29338 480 29368
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 1577 29338 1643 29341
rect 0 29336 1643 29338
rect 0 29280 1582 29336
rect 1638 29280 1643 29336
rect 0 29278 1643 29280
rect 0 29248 480 29278
rect 1577 29275 1643 29278
rect 9581 29202 9647 29205
rect 11237 29202 11303 29205
rect 9581 29200 11303 29202
rect 9581 29144 9586 29200
rect 9642 29144 11242 29200
rect 11298 29144 11303 29200
rect 9581 29142 11303 29144
rect 9581 29139 9647 29142
rect 11237 29139 11303 29142
rect 1761 29066 1827 29069
rect 2865 29066 2931 29069
rect 7741 29066 7807 29069
rect 8293 29066 8359 29069
rect 10409 29066 10475 29069
rect 1761 29064 10475 29066
rect 1761 29008 1766 29064
rect 1822 29008 2870 29064
rect 2926 29008 7746 29064
rect 7802 29008 8298 29064
rect 8354 29008 10414 29064
rect 10470 29008 10475 29064
rect 1761 29006 10475 29008
rect 1761 29003 1827 29006
rect 2865 29003 2931 29006
rect 7741 29003 7807 29006
rect 8293 29003 8359 29006
rect 10409 29003 10475 29006
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 6361 28386 6427 28389
rect 8385 28386 8451 28389
rect 6361 28384 8451 28386
rect 6361 28328 6366 28384
rect 6422 28328 8390 28384
rect 8446 28328 8451 28384
rect 6361 28326 8451 28328
rect 6361 28323 6427 28326
rect 8385 28323 8451 28326
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 4981 28250 5047 28253
rect 5717 28250 5783 28253
rect 4981 28248 8034 28250
rect 4981 28192 4986 28248
rect 5042 28192 5722 28248
rect 5778 28192 8034 28248
rect 4981 28190 8034 28192
rect 4981 28187 5047 28190
rect 5717 28187 5783 28190
rect 2957 28114 3023 28117
rect 7741 28114 7807 28117
rect 2957 28112 7807 28114
rect 2957 28056 2962 28112
rect 3018 28056 7746 28112
rect 7802 28056 7807 28112
rect 2957 28054 7807 28056
rect 7974 28114 8034 28190
rect 9581 28114 9647 28117
rect 7974 28112 9647 28114
rect 7974 28056 9586 28112
rect 9642 28056 9647 28112
rect 7974 28054 9647 28056
rect 2957 28051 3023 28054
rect 7741 28051 7807 28054
rect 9581 28051 9647 28054
rect 5809 27978 5875 27981
rect 6729 27978 6795 27981
rect 5809 27976 6795 27978
rect 5809 27920 5814 27976
rect 5870 27920 6734 27976
rect 6790 27920 6795 27976
rect 5809 27918 6795 27920
rect 5809 27915 5875 27918
rect 6729 27915 6795 27918
rect 8569 27842 8635 27845
rect 9673 27842 9739 27845
rect 10501 27842 10567 27845
rect 8569 27840 10567 27842
rect 8569 27784 8574 27840
rect 8630 27784 9678 27840
rect 9734 27784 10506 27840
rect 10562 27784 10567 27840
rect 8569 27782 10567 27784
rect 8569 27779 8635 27782
rect 9673 27779 9739 27782
rect 10501 27779 10567 27782
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 8702 27644 8708 27708
rect 8772 27706 8778 27708
rect 9305 27706 9371 27709
rect 8772 27704 9371 27706
rect 8772 27648 9310 27704
rect 9366 27648 9371 27704
rect 8772 27646 9371 27648
rect 8772 27644 8778 27646
rect 9305 27643 9371 27646
rect 7373 27570 7439 27573
rect 10041 27570 10107 27573
rect 7373 27568 10107 27570
rect 7373 27512 7378 27568
rect 7434 27512 10046 27568
rect 10102 27512 10107 27568
rect 7373 27510 10107 27512
rect 7373 27507 7439 27510
rect 10041 27507 10107 27510
rect 2773 27434 2839 27437
rect 7465 27434 7531 27437
rect 9673 27434 9739 27437
rect 2773 27432 9739 27434
rect 2773 27376 2778 27432
rect 2834 27376 7470 27432
rect 7526 27376 9678 27432
rect 9734 27376 9739 27432
rect 2773 27374 9739 27376
rect 2773 27371 2839 27374
rect 7465 27371 7531 27374
rect 9673 27371 9739 27374
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 11329 27162 11395 27165
rect 12985 27162 13051 27165
rect 11329 27160 13051 27162
rect 11329 27104 11334 27160
rect 11390 27104 12990 27160
rect 13046 27104 13051 27160
rect 11329 27102 13051 27104
rect 11329 27099 11395 27102
rect 12985 27099 13051 27102
rect 0 27026 480 27056
rect 1577 27026 1643 27029
rect 0 27024 1643 27026
rect 0 26968 1582 27024
rect 1638 26968 1643 27024
rect 0 26966 1643 26968
rect 0 26936 480 26966
rect 1577 26963 1643 26966
rect 7281 27026 7347 27029
rect 13169 27026 13235 27029
rect 7281 27024 13235 27026
rect 7281 26968 7286 27024
rect 7342 26968 13174 27024
rect 13230 26968 13235 27024
rect 7281 26966 13235 26968
rect 7281 26963 7347 26966
rect 13169 26963 13235 26966
rect 7005 26890 7071 26893
rect 12249 26890 12315 26893
rect 12801 26890 12867 26893
rect 7005 26888 12867 26890
rect 7005 26832 7010 26888
rect 7066 26832 12254 26888
rect 12310 26832 12806 26888
rect 12862 26832 12867 26888
rect 7005 26830 12867 26832
rect 7005 26827 7071 26830
rect 12249 26827 12315 26830
rect 12801 26827 12867 26830
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 10174 26556 10180 26620
rect 10244 26618 10250 26620
rect 10593 26618 10659 26621
rect 10244 26616 10659 26618
rect 10244 26560 10598 26616
rect 10654 26560 10659 26616
rect 10244 26558 10659 26560
rect 10244 26556 10250 26558
rect 10593 26555 10659 26558
rect 10593 26482 10659 26485
rect 12433 26482 12499 26485
rect 10593 26480 12499 26482
rect 10593 26424 10598 26480
rect 10654 26424 12438 26480
rect 12494 26424 12499 26480
rect 10593 26422 12499 26424
rect 10593 26419 10659 26422
rect 12433 26419 12499 26422
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 1853 25938 1919 25941
rect 8569 25938 8635 25941
rect 1853 25936 8635 25938
rect 1853 25880 1858 25936
rect 1914 25880 8574 25936
rect 8630 25880 8635 25936
rect 1853 25878 8635 25880
rect 1853 25875 1919 25878
rect 8569 25875 8635 25878
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 7281 25258 7347 25261
rect 13261 25258 13327 25261
rect 15009 25258 15075 25261
rect 7281 25256 15075 25258
rect 7281 25200 7286 25256
rect 7342 25200 13266 25256
rect 13322 25200 15014 25256
rect 15070 25200 15075 25256
rect 7281 25198 15075 25200
rect 7281 25195 7347 25198
rect 13261 25195 13327 25198
rect 15009 25195 15075 25198
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 9397 24986 9463 24989
rect 13445 24986 13511 24989
rect 9397 24984 13511 24986
rect 9397 24928 9402 24984
rect 9458 24928 13450 24984
rect 13506 24928 13511 24984
rect 9397 24926 13511 24928
rect 9397 24923 9463 24926
rect 13445 24923 13511 24926
rect 5073 24850 5139 24853
rect 6085 24850 6151 24853
rect 13813 24850 13879 24853
rect 5073 24848 13879 24850
rect 5073 24792 5078 24848
rect 5134 24792 6090 24848
rect 6146 24792 13818 24848
rect 13874 24792 13879 24848
rect 5073 24790 13879 24792
rect 5073 24787 5139 24790
rect 6085 24787 6151 24790
rect 13813 24787 13879 24790
rect 0 24578 480 24608
rect 1577 24578 1643 24581
rect 0 24576 1643 24578
rect 0 24520 1582 24576
rect 1638 24520 1643 24576
rect 0 24518 1643 24520
rect 0 24488 480 24518
rect 1577 24515 1643 24518
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 9397 23354 9463 23357
rect 10225 23354 10291 23357
rect 11053 23354 11119 23357
rect 9397 23352 11119 23354
rect 9397 23296 9402 23352
rect 9458 23296 10230 23352
rect 10286 23296 11058 23352
rect 11114 23296 11119 23352
rect 9397 23294 11119 23296
rect 9397 23291 9463 23294
rect 10225 23291 10291 23294
rect 11053 23291 11119 23294
rect 7465 23218 7531 23221
rect 12157 23218 12223 23221
rect 7465 23216 12223 23218
rect 7465 23160 7470 23216
rect 7526 23160 12162 23216
rect 12218 23160 12223 23216
rect 7465 23158 12223 23160
rect 7465 23155 7531 23158
rect 12157 23155 12223 23158
rect 7097 23082 7163 23085
rect 9673 23082 9739 23085
rect 7097 23080 9739 23082
rect 7097 23024 7102 23080
rect 7158 23024 9678 23080
rect 9734 23024 9739 23080
rect 7097 23022 9739 23024
rect 7097 23019 7163 23022
rect 9673 23019 9739 23022
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 1669 22674 1735 22677
rect 5717 22674 5783 22677
rect 1669 22672 5783 22674
rect 1669 22616 1674 22672
rect 1730 22616 5722 22672
rect 5778 22616 5783 22672
rect 1669 22614 5783 22616
rect 1669 22611 1735 22614
rect 5717 22611 5783 22614
rect 2773 22538 2839 22541
rect 10869 22538 10935 22541
rect 2773 22536 10935 22538
rect 2773 22480 2778 22536
rect 2834 22480 10874 22536
rect 10930 22480 10935 22536
rect 2773 22478 10935 22480
rect 2773 22475 2839 22478
rect 10550 22405 10610 22478
rect 10869 22475 10935 22478
rect 9765 22404 9831 22405
rect 9765 22402 9812 22404
rect 9720 22400 9812 22402
rect 9720 22344 9770 22400
rect 9720 22342 9812 22344
rect 9765 22340 9812 22342
rect 9876 22340 9882 22404
rect 10501 22400 10610 22405
rect 10501 22344 10506 22400
rect 10562 22344 10610 22400
rect 10501 22342 10610 22344
rect 9765 22339 9831 22340
rect 10501 22339 10567 22342
rect 6277 22336 6597 22337
rect 0 22266 480 22296
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 0 22206 858 22266
rect 0 22176 480 22206
rect 798 22130 858 22206
rect 9397 22130 9463 22133
rect 9581 22130 9647 22133
rect 798 22070 1410 22130
rect 1350 21994 1410 22070
rect 9397 22128 9647 22130
rect 9397 22072 9402 22128
rect 9458 22072 9586 22128
rect 9642 22072 9647 22128
rect 9397 22070 9647 22072
rect 9397 22067 9463 22070
rect 9581 22067 9647 22070
rect 9765 22130 9831 22133
rect 10685 22130 10751 22133
rect 9765 22128 10751 22130
rect 9765 22072 9770 22128
rect 9826 22072 10690 22128
rect 10746 22072 10751 22128
rect 9765 22070 10751 22072
rect 9765 22067 9831 22070
rect 10685 22067 10751 22070
rect 1577 21994 1643 21997
rect 1350 21992 1643 21994
rect 1350 21936 1582 21992
rect 1638 21936 1643 21992
rect 1350 21934 1643 21936
rect 1577 21931 1643 21934
rect 8201 21994 8267 21997
rect 11881 21994 11947 21997
rect 8201 21992 11947 21994
rect 8201 21936 8206 21992
rect 8262 21936 11886 21992
rect 11942 21936 11947 21992
rect 8201 21934 11947 21936
rect 8201 21931 8267 21934
rect 11881 21931 11947 21934
rect 9673 21858 9739 21861
rect 9857 21858 9923 21861
rect 10133 21860 10199 21861
rect 10133 21858 10180 21860
rect 9673 21856 9923 21858
rect 9673 21800 9678 21856
rect 9734 21800 9862 21856
rect 9918 21800 9923 21856
rect 9673 21798 9923 21800
rect 10088 21856 10180 21858
rect 10088 21800 10138 21856
rect 10088 21798 10180 21800
rect 9673 21795 9739 21798
rect 9857 21795 9923 21798
rect 10133 21796 10180 21798
rect 10244 21796 10250 21860
rect 10133 21795 10199 21796
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 9857 21724 9923 21725
rect 9806 21722 9812 21724
rect 9766 21662 9812 21722
rect 9876 21720 9923 21724
rect 10593 21722 10659 21725
rect 9918 21664 9923 21720
rect 9806 21660 9812 21662
rect 9876 21660 9923 21664
rect 9857 21659 9923 21660
rect 10550 21720 10659 21722
rect 10550 21664 10598 21720
rect 10654 21664 10659 21720
rect 10550 21659 10659 21664
rect 4889 21586 4955 21589
rect 9765 21586 9831 21589
rect 4889 21584 9831 21586
rect 4889 21528 4894 21584
rect 4950 21528 9770 21584
rect 9826 21528 9831 21584
rect 4889 21526 9831 21528
rect 4889 21523 4955 21526
rect 9765 21523 9831 21526
rect 5533 21450 5599 21453
rect 9581 21452 9647 21453
rect 5533 21448 7666 21450
rect 5533 21392 5538 21448
rect 5594 21392 7666 21448
rect 5533 21390 7666 21392
rect 5533 21387 5599 21390
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 7606 21178 7666 21390
rect 9581 21448 9628 21452
rect 9692 21450 9698 21452
rect 9581 21392 9586 21448
rect 9581 21388 9628 21392
rect 9692 21390 9774 21450
rect 9692 21388 9698 21390
rect 9581 21387 9647 21388
rect 7741 21314 7807 21317
rect 10550 21314 10610 21659
rect 7741 21312 10610 21314
rect 7741 21256 7746 21312
rect 7802 21256 10610 21312
rect 7741 21254 10610 21256
rect 7741 21251 7807 21254
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 10961 21178 11027 21181
rect 7606 21176 11027 21178
rect 7606 21120 10966 21176
rect 11022 21120 11027 21176
rect 7606 21118 11027 21120
rect 10961 21115 11027 21118
rect 5901 21042 5967 21045
rect 9622 21042 9628 21044
rect 5901 21040 9628 21042
rect 5901 20984 5906 21040
rect 5962 20984 9628 21040
rect 5901 20982 9628 20984
rect 5901 20979 5967 20982
rect 9622 20980 9628 20982
rect 9692 21042 9698 21044
rect 10501 21042 10567 21045
rect 9692 21040 10567 21042
rect 9692 20984 10506 21040
rect 10562 20984 10567 21040
rect 9692 20982 10567 20984
rect 9692 20980 9698 20982
rect 10501 20979 10567 20982
rect 1669 20906 1735 20909
rect 9673 20906 9739 20909
rect 1669 20904 9739 20906
rect 1669 20848 1674 20904
rect 1730 20848 9678 20904
rect 9734 20848 9739 20904
rect 1669 20846 9739 20848
rect 1669 20843 1735 20846
rect 9673 20843 9739 20846
rect 10593 20906 10659 20909
rect 12433 20906 12499 20909
rect 10593 20904 12499 20906
rect 10593 20848 10598 20904
rect 10654 20848 12438 20904
rect 12494 20848 12499 20904
rect 10593 20846 12499 20848
rect 10593 20843 10659 20846
rect 12433 20843 12499 20846
rect 8661 20772 8727 20773
rect 8661 20770 8708 20772
rect 8616 20768 8708 20770
rect 8616 20712 8666 20768
rect 8616 20710 8708 20712
rect 8661 20708 8708 20710
rect 8772 20708 8778 20772
rect 8661 20707 8727 20708
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 10041 20362 10107 20365
rect 12893 20362 12959 20365
rect 10041 20360 12959 20362
rect 10041 20304 10046 20360
rect 10102 20304 12898 20360
rect 12954 20304 12959 20360
rect 10041 20302 12959 20304
rect 10041 20299 10107 20302
rect 12893 20299 12959 20302
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 13445 20090 13511 20093
rect 15520 20090 16000 20120
rect 13445 20088 16000 20090
rect 13445 20032 13450 20088
rect 13506 20032 16000 20088
rect 13445 20030 16000 20032
rect 13445 20027 13511 20030
rect 15520 20000 16000 20030
rect 0 19954 480 19984
rect 1577 19954 1643 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 480 19894
rect 1577 19891 1643 19894
rect 10501 19954 10567 19957
rect 13169 19954 13235 19957
rect 10501 19952 13235 19954
rect 10501 19896 10506 19952
rect 10562 19896 13174 19952
rect 13230 19896 13235 19952
rect 10501 19894 13235 19896
rect 10501 19891 10567 19894
rect 13169 19891 13235 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 9806 19076 9812 19140
rect 9876 19138 9882 19140
rect 10133 19138 10199 19141
rect 9876 19136 10199 19138
rect 9876 19080 10138 19136
rect 10194 19080 10199 19136
rect 9876 19078 10199 19080
rect 9876 19076 9882 19078
rect 10133 19075 10199 19078
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 9990 18940 9996 19004
rect 10060 19002 10066 19004
rect 10225 19002 10291 19005
rect 10060 19000 10291 19002
rect 10060 18944 10230 19000
rect 10286 18944 10291 19000
rect 10060 18942 10291 18944
rect 10060 18940 10066 18942
rect 10225 18939 10291 18942
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 1945 18322 2011 18325
rect 7833 18322 7899 18325
rect 1945 18320 7899 18322
rect 1945 18264 1950 18320
rect 2006 18264 7838 18320
rect 7894 18264 7899 18320
rect 1945 18262 7899 18264
rect 1945 18259 2011 18262
rect 7833 18259 7899 18262
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 7649 17914 7715 17917
rect 9857 17914 9923 17917
rect 7649 17912 9923 17914
rect 7649 17856 7654 17912
rect 7710 17856 9862 17912
rect 9918 17856 9923 17912
rect 7649 17854 9923 17856
rect 7649 17851 7715 17854
rect 9857 17851 9923 17854
rect 5533 17778 5599 17781
rect 11421 17778 11487 17781
rect 5533 17776 11487 17778
rect 5533 17720 5538 17776
rect 5594 17720 11426 17776
rect 11482 17720 11487 17776
rect 5533 17718 11487 17720
rect 5533 17715 5599 17718
rect 11421 17715 11487 17718
rect 0 17642 480 17672
rect 1577 17642 1643 17645
rect 0 17640 1643 17642
rect 0 17584 1582 17640
rect 1638 17584 1643 17640
rect 0 17582 1643 17584
rect 0 17552 480 17582
rect 1577 17579 1643 17582
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 9489 17098 9555 17101
rect 10961 17098 11027 17101
rect 9489 17096 11027 17098
rect 9489 17040 9494 17096
rect 9550 17040 10966 17096
rect 11022 17040 11027 17096
rect 9489 17038 11027 17040
rect 9489 17035 9555 17038
rect 10961 17035 11027 17038
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 8385 16690 8451 16693
rect 10225 16690 10291 16693
rect 8385 16688 10291 16690
rect 8385 16632 8390 16688
rect 8446 16632 10230 16688
rect 10286 16632 10291 16688
rect 8385 16630 10291 16632
rect 8385 16627 8451 16630
rect 10225 16627 10291 16630
rect 10777 16690 10843 16693
rect 13169 16690 13235 16693
rect 10777 16688 13235 16690
rect 10777 16632 10782 16688
rect 10838 16632 13174 16688
rect 13230 16632 13235 16688
rect 10777 16630 13235 16632
rect 10777 16627 10843 16630
rect 13169 16627 13235 16630
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 1945 16146 2011 16149
rect 10317 16146 10383 16149
rect 1945 16144 10383 16146
rect 1945 16088 1950 16144
rect 2006 16088 10322 16144
rect 10378 16088 10383 16144
rect 1945 16086 10383 16088
rect 1945 16083 2011 16086
rect 10317 16083 10383 16086
rect 4705 16010 4771 16013
rect 7649 16010 7715 16013
rect 4705 16008 7715 16010
rect 4705 15952 4710 16008
rect 4766 15952 7654 16008
rect 7710 15952 7715 16008
rect 4705 15950 7715 15952
rect 4705 15947 4771 15950
rect 7649 15947 7715 15950
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 7557 15602 7623 15605
rect 9806 15602 9812 15604
rect 7557 15600 9812 15602
rect 7557 15544 7562 15600
rect 7618 15544 9812 15600
rect 7557 15542 9812 15544
rect 7557 15539 7623 15542
rect 9806 15540 9812 15542
rect 9876 15540 9882 15604
rect 12249 15468 12315 15469
rect 12198 15404 12204 15468
rect 12268 15466 12315 15468
rect 12268 15464 12360 15466
rect 12310 15408 12360 15464
rect 12268 15406 12360 15408
rect 12268 15404 12315 15406
rect 12249 15403 12315 15404
rect 7925 15330 7991 15333
rect 8702 15330 8708 15332
rect 7925 15328 8708 15330
rect 7925 15272 7930 15328
rect 7986 15272 8708 15328
rect 7925 15270 8708 15272
rect 7925 15267 7991 15270
rect 8702 15268 8708 15270
rect 8772 15268 8778 15332
rect 3610 15264 3930 15265
rect 0 15194 480 15224
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 1577 15194 1643 15197
rect 0 15192 1643 15194
rect 0 15136 1582 15192
rect 1638 15136 1643 15192
rect 0 15134 1643 15136
rect 0 15104 480 15134
rect 1577 15131 1643 15134
rect 5349 15058 5415 15061
rect 9990 15058 9996 15060
rect 5349 15056 9996 15058
rect 5349 15000 5354 15056
rect 5410 15000 9996 15056
rect 5349 14998 9996 15000
rect 5349 14995 5415 14998
rect 2129 14922 2195 14925
rect 4613 14922 4679 14925
rect 2129 14920 4679 14922
rect 2129 14864 2134 14920
rect 2190 14864 4618 14920
rect 4674 14864 4679 14920
rect 2129 14862 4679 14864
rect 2129 14859 2195 14862
rect 4613 14859 4679 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 6545 14514 6611 14517
rect 6686 14514 6746 14998
rect 9990 14996 9996 14998
rect 10060 14996 10066 15060
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 6545 14512 6746 14514
rect 6545 14456 6550 14512
rect 6606 14456 6746 14512
rect 6545 14454 6746 14456
rect 6545 14451 6611 14454
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 4981 13834 5047 13837
rect 11237 13834 11303 13837
rect 4981 13832 11303 13834
rect 4981 13776 4986 13832
rect 5042 13776 11242 13832
rect 11298 13776 11303 13832
rect 4981 13774 11303 13776
rect 4981 13771 5047 13774
rect 11237 13771 11303 13774
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 0 12882 480 12912
rect 2773 12882 2839 12885
rect 0 12880 2839 12882
rect 0 12824 2778 12880
rect 2834 12824 2839 12880
rect 0 12822 2839 12824
rect 0 12792 480 12822
rect 2773 12819 2839 12822
rect 5441 12746 5507 12749
rect 5809 12746 5875 12749
rect 8477 12746 8543 12749
rect 9581 12746 9647 12749
rect 5441 12744 8543 12746
rect 5441 12688 5446 12744
rect 5502 12688 5814 12744
rect 5870 12688 8482 12744
rect 8538 12688 8543 12744
rect 5441 12686 8543 12688
rect 5441 12683 5507 12686
rect 5809 12683 5875 12686
rect 8477 12683 8543 12686
rect 9446 12744 9647 12746
rect 9446 12688 9586 12744
rect 9642 12688 9647 12744
rect 9446 12686 9647 12688
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 9446 12477 9506 12686
rect 9581 12683 9647 12686
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 1669 12474 1735 12477
rect 5165 12474 5231 12477
rect 1669 12472 5231 12474
rect 1669 12416 1674 12472
rect 1730 12416 5170 12472
rect 5226 12416 5231 12472
rect 1669 12414 5231 12416
rect 9446 12472 9555 12477
rect 9446 12416 9494 12472
rect 9550 12416 9555 12472
rect 9446 12414 9555 12416
rect 1669 12411 1735 12414
rect 5165 12411 5231 12414
rect 9489 12411 9555 12414
rect 5349 12338 5415 12341
rect 11053 12338 11119 12341
rect 12065 12338 12131 12341
rect 5349 12336 12131 12338
rect 5349 12280 5354 12336
rect 5410 12280 11058 12336
rect 11114 12280 12070 12336
rect 12126 12280 12131 12336
rect 5349 12278 12131 12280
rect 5349 12275 5415 12278
rect 11053 12275 11119 12278
rect 12065 12275 12131 12278
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 5441 11794 5507 11797
rect 10317 11794 10383 11797
rect 5441 11792 10383 11794
rect 5441 11736 5446 11792
rect 5502 11736 10322 11792
rect 10378 11736 10383 11792
rect 5441 11734 10383 11736
rect 5441 11731 5507 11734
rect 10317 11731 10383 11734
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 8109 10706 8175 10709
rect 12341 10706 12407 10709
rect 8109 10704 12407 10706
rect 8109 10648 8114 10704
rect 8170 10648 12346 10704
rect 12402 10648 12407 10704
rect 8109 10646 12407 10648
rect 8109 10643 8175 10646
rect 12341 10643 12407 10646
rect 0 10570 480 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 480 10510
rect 1577 10507 1643 10510
rect 6453 10570 6519 10573
rect 12249 10570 12315 10573
rect 6453 10568 12315 10570
rect 6453 10512 6458 10568
rect 6514 10512 12254 10568
rect 12310 10512 12315 10568
rect 6453 10510 12315 10512
rect 6453 10507 6519 10510
rect 12249 10507 12315 10510
rect 12249 10436 12315 10437
rect 12198 10434 12204 10436
rect 12158 10374 12204 10434
rect 12268 10432 12315 10436
rect 12310 10376 12315 10432
rect 12198 10372 12204 10374
rect 12268 10372 12315 10376
rect 12249 10371 12315 10372
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 8109 10298 8175 10301
rect 9489 10298 9555 10301
rect 8109 10296 9555 10298
rect 8109 10240 8114 10296
rect 8170 10240 9494 10296
rect 9550 10240 9555 10296
rect 8109 10238 9555 10240
rect 8109 10235 8175 10238
rect 9489 10235 9555 10238
rect 8702 10100 8708 10164
rect 8772 10162 8778 10164
rect 13721 10162 13787 10165
rect 8772 10160 13787 10162
rect 8772 10104 13726 10160
rect 13782 10104 13787 10160
rect 8772 10102 13787 10104
rect 8772 10100 8778 10102
rect 13721 10099 13787 10102
rect 8661 10026 8727 10029
rect 12065 10026 12131 10029
rect 8661 10024 12131 10026
rect 8661 9968 8666 10024
rect 8722 9968 12070 10024
rect 12126 9968 12131 10024
rect 8661 9966 12131 9968
rect 8661 9963 8727 9966
rect 12065 9963 12131 9966
rect 12341 10026 12407 10029
rect 12893 10026 12959 10029
rect 12341 10024 12959 10026
rect 12341 9968 12346 10024
rect 12402 9968 12898 10024
rect 12954 9968 12959 10024
rect 12341 9966 12959 9968
rect 12341 9963 12407 9966
rect 12893 9963 12959 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 3325 9482 3391 9485
rect 7925 9482 7991 9485
rect 3325 9480 7991 9482
rect 3325 9424 3330 9480
rect 3386 9424 7930 9480
rect 7986 9424 7991 9480
rect 3325 9422 7991 9424
rect 3325 9419 3391 9422
rect 7925 9419 7991 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 5625 8938 5691 8941
rect 11973 8938 12039 8941
rect 5625 8936 12039 8938
rect 5625 8880 5630 8936
rect 5686 8880 11978 8936
rect 12034 8880 12039 8936
rect 5625 8878 12039 8880
rect 5625 8875 5691 8878
rect 11973 8875 12039 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 2773 8530 2839 8533
rect 7649 8530 7715 8533
rect 8109 8530 8175 8533
rect 2773 8528 8175 8530
rect 2773 8472 2778 8528
rect 2834 8472 7654 8528
rect 7710 8472 8114 8528
rect 8170 8472 8175 8528
rect 2773 8470 8175 8472
rect 2773 8467 2839 8470
rect 7649 8467 7715 8470
rect 8109 8467 8175 8470
rect 9438 8468 9444 8532
rect 9508 8530 9514 8532
rect 9581 8530 9647 8533
rect 9508 8528 9647 8530
rect 9508 8472 9586 8528
rect 9642 8472 9647 8528
rect 9508 8470 9647 8472
rect 9508 8468 9514 8470
rect 9581 8467 9647 8470
rect 3785 8394 3851 8397
rect 9305 8394 9371 8397
rect 3785 8392 9371 8394
rect 3785 8336 3790 8392
rect 3846 8336 9310 8392
rect 9366 8336 9371 8392
rect 3785 8334 9371 8336
rect 3785 8331 3851 8334
rect 9305 8331 9371 8334
rect 6277 8192 6597 8193
rect 0 8122 480 8152
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 2773 8122 2839 8125
rect 0 8120 2839 8122
rect 0 8064 2778 8120
rect 2834 8064 2839 8120
rect 0 8062 2839 8064
rect 0 8032 480 8062
rect 2773 8059 2839 8062
rect 7097 8122 7163 8125
rect 10133 8122 10199 8125
rect 7097 8120 10199 8122
rect 7097 8064 7102 8120
rect 7158 8064 10138 8120
rect 10194 8064 10199 8120
rect 7097 8062 10199 8064
rect 7097 8059 7163 8062
rect 10133 8059 10199 8062
rect 7373 7986 7439 7989
rect 7925 7986 7991 7989
rect 8385 7986 8451 7989
rect 7373 7984 8451 7986
rect 7373 7928 7378 7984
rect 7434 7928 7930 7984
rect 7986 7928 8390 7984
rect 8446 7928 8451 7984
rect 7373 7926 8451 7928
rect 7373 7923 7439 7926
rect 7925 7923 7991 7926
rect 8385 7923 8451 7926
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 3049 7306 3115 7309
rect 8753 7306 8819 7309
rect 3049 7304 8819 7306
rect 3049 7248 3054 7304
rect 3110 7248 8758 7304
rect 8814 7248 8819 7304
rect 3049 7246 8819 7248
rect 3049 7243 3115 7246
rect 8753 7243 8819 7246
rect 1945 7170 2011 7173
rect 5533 7170 5599 7173
rect 1945 7168 5599 7170
rect 1945 7112 1950 7168
rect 2006 7112 5538 7168
rect 5594 7112 5599 7168
rect 1945 7110 5599 7112
rect 1945 7107 2011 7110
rect 5533 7107 5599 7110
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 2865 6898 2931 6901
rect 4061 6898 4127 6901
rect 8845 6898 8911 6901
rect 2865 6896 8911 6898
rect 2865 6840 2870 6896
rect 2926 6840 4066 6896
rect 4122 6840 8850 6896
rect 8906 6840 8911 6896
rect 2865 6838 8911 6840
rect 2865 6835 2931 6838
rect 4061 6835 4127 6838
rect 8845 6835 8911 6838
rect 11973 6898 12039 6901
rect 11973 6896 15394 6898
rect 11973 6840 11978 6896
rect 12034 6840 15394 6896
rect 11973 6838 15394 6840
rect 11973 6835 12039 6838
rect 7097 6762 7163 6765
rect 12249 6762 12315 6765
rect 7097 6760 12315 6762
rect 7097 6704 7102 6760
rect 7158 6704 12254 6760
rect 12310 6704 12315 6760
rect 7097 6702 12315 6704
rect 15334 6762 15394 6838
rect 15520 6762 16000 6792
rect 15334 6702 16000 6762
rect 7097 6699 7163 6702
rect 12249 6699 12315 6702
rect 15520 6672 16000 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 8293 6354 8359 6357
rect 10041 6354 10107 6357
rect 8293 6352 10107 6354
rect 8293 6296 8298 6352
rect 8354 6296 10046 6352
rect 10102 6296 10107 6352
rect 8293 6294 10107 6296
rect 8293 6291 8359 6294
rect 10041 6291 10107 6294
rect 4613 6218 4679 6221
rect 9765 6218 9831 6221
rect 4613 6216 9831 6218
rect 4613 6160 4618 6216
rect 4674 6160 9770 6216
rect 9826 6160 9831 6216
rect 4613 6158 9831 6160
rect 4613 6155 4679 6158
rect 9765 6155 9831 6158
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 0 5810 480 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 480 5750
rect 1577 5747 1643 5750
rect 5441 5674 5507 5677
rect 6821 5674 6887 5677
rect 5441 5672 6887 5674
rect 5441 5616 5446 5672
rect 5502 5616 6826 5672
rect 6882 5616 6887 5672
rect 5441 5614 6887 5616
rect 5441 5611 5507 5614
rect 6821 5611 6887 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 8201 5402 8267 5405
rect 7928 5400 8267 5402
rect 7928 5344 8206 5400
rect 8262 5344 8267 5400
rect 7928 5342 8267 5344
rect 7741 5266 7807 5269
rect 7928 5266 7988 5342
rect 8201 5339 8267 5342
rect 7741 5264 7988 5266
rect 7741 5208 7746 5264
rect 7802 5208 7988 5264
rect 7741 5206 7988 5208
rect 8201 5266 8267 5269
rect 8937 5266 9003 5269
rect 11053 5266 11119 5269
rect 11605 5266 11671 5269
rect 8201 5264 11671 5266
rect 8201 5208 8206 5264
rect 8262 5208 8942 5264
rect 8998 5208 11058 5264
rect 11114 5208 11610 5264
rect 11666 5208 11671 5264
rect 8201 5206 11671 5208
rect 7741 5203 7807 5206
rect 8201 5203 8267 5206
rect 8937 5203 9003 5206
rect 11053 5203 11119 5206
rect 11605 5203 11671 5206
rect 8661 5130 8727 5133
rect 10317 5130 10383 5133
rect 8661 5128 10383 5130
rect 8661 5072 8666 5128
rect 8722 5072 10322 5128
rect 10378 5072 10383 5128
rect 8661 5070 10383 5072
rect 8661 5067 8727 5070
rect 10317 5067 10383 5070
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 1761 4722 1827 4725
rect 8385 4722 8451 4725
rect 1761 4720 8451 4722
rect 1761 4664 1766 4720
rect 1822 4664 8390 4720
rect 8446 4664 8451 4720
rect 1761 4662 8451 4664
rect 1761 4659 1827 4662
rect 8385 4659 8451 4662
rect 1393 4586 1459 4589
rect 6177 4586 6243 4589
rect 1393 4584 6243 4586
rect 1393 4528 1398 4584
rect 1454 4528 6182 4584
rect 6238 4528 6243 4584
rect 1393 4526 6243 4528
rect 1393 4523 1459 4526
rect 6177 4523 6243 4526
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 565 4314 631 4317
rect 3049 4314 3115 4317
rect 565 4312 3115 4314
rect 565 4256 570 4312
rect 626 4256 3054 4312
rect 3110 4256 3115 4312
rect 565 4254 3115 4256
rect 565 4251 631 4254
rect 3049 4251 3115 4254
rect 2313 4178 2379 4181
rect 4797 4178 4863 4181
rect 7281 4178 7347 4181
rect 2313 4176 7347 4178
rect 2313 4120 2318 4176
rect 2374 4120 4802 4176
rect 4858 4120 7286 4176
rect 7342 4120 7347 4176
rect 2313 4118 7347 4120
rect 2313 4115 2379 4118
rect 4797 4115 4863 4118
rect 7281 4115 7347 4118
rect 10409 4178 10475 4181
rect 12893 4178 12959 4181
rect 10409 4176 12959 4178
rect 10409 4120 10414 4176
rect 10470 4120 12898 4176
rect 12954 4120 12959 4176
rect 10409 4118 12959 4120
rect 10409 4115 10475 4118
rect 12893 4115 12959 4118
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 3601 3770 3667 3773
rect 5533 3770 5599 3773
rect 3601 3768 5599 3770
rect 3601 3712 3606 3768
rect 3662 3712 5538 3768
rect 5594 3712 5599 3768
rect 3601 3710 5599 3712
rect 3601 3707 3667 3710
rect 5533 3707 5599 3710
rect 7281 3770 7347 3773
rect 8753 3770 8819 3773
rect 10777 3770 10843 3773
rect 7281 3768 8819 3770
rect 7281 3712 7286 3768
rect 7342 3712 8758 3768
rect 8814 3712 8819 3768
rect 7281 3710 8819 3712
rect 7281 3707 7347 3710
rect 8753 3707 8819 3710
rect 8894 3768 10843 3770
rect 8894 3712 10782 3768
rect 10838 3712 10843 3768
rect 8894 3710 10843 3712
rect 5257 3634 5323 3637
rect 8894 3634 8954 3710
rect 10777 3707 10843 3710
rect 5257 3632 8954 3634
rect 5257 3576 5262 3632
rect 5318 3576 8954 3632
rect 5257 3574 8954 3576
rect 9397 3634 9463 3637
rect 15377 3634 15443 3637
rect 9397 3632 15443 3634
rect 9397 3576 9402 3632
rect 9458 3576 15382 3632
rect 15438 3576 15443 3632
rect 9397 3574 15443 3576
rect 5257 3571 5323 3574
rect 9397 3571 9463 3574
rect 15377 3571 15443 3574
rect 0 3498 480 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 480 3438
rect 1485 3435 1551 3438
rect 2313 3498 2379 3501
rect 5625 3498 5691 3501
rect 2313 3496 5691 3498
rect 2313 3440 2318 3496
rect 2374 3440 5630 3496
rect 5686 3440 5691 3496
rect 2313 3438 5691 3440
rect 2313 3435 2379 3438
rect 5625 3435 5691 3438
rect 7097 3498 7163 3501
rect 10501 3498 10567 3501
rect 7097 3496 10567 3498
rect 7097 3440 7102 3496
rect 7158 3440 10506 3496
rect 10562 3440 10567 3496
rect 7097 3438 10567 3440
rect 7097 3435 7163 3438
rect 10501 3435 10567 3438
rect 10777 3498 10843 3501
rect 13997 3498 14063 3501
rect 10777 3496 14063 3498
rect 10777 3440 10782 3496
rect 10838 3440 14002 3496
rect 14058 3440 14063 3496
rect 10777 3438 14063 3440
rect 10777 3435 10843 3438
rect 13997 3435 14063 3438
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 9438 3164 9444 3228
rect 9508 3226 9514 3228
rect 10685 3226 10751 3229
rect 12801 3226 12867 3229
rect 9508 3166 9874 3226
rect 9508 3164 9514 3166
rect 3049 3090 3115 3093
rect 6637 3090 6703 3093
rect 3049 3088 6703 3090
rect 3049 3032 3054 3088
rect 3110 3032 6642 3088
rect 6698 3032 6703 3088
rect 3049 3030 6703 3032
rect 3049 3027 3115 3030
rect 6637 3027 6703 3030
rect 6913 3090 6979 3093
rect 9673 3090 9739 3093
rect 6913 3088 9739 3090
rect 6913 3032 6918 3088
rect 6974 3032 9678 3088
rect 9734 3032 9739 3088
rect 6913 3030 9739 3032
rect 9814 3090 9874 3166
rect 10685 3224 12867 3226
rect 10685 3168 10690 3224
rect 10746 3168 12806 3224
rect 12862 3168 12867 3224
rect 10685 3166 12867 3168
rect 10685 3163 10751 3166
rect 12801 3163 12867 3166
rect 11329 3090 11395 3093
rect 9814 3088 11395 3090
rect 9814 3032 11334 3088
rect 11390 3032 11395 3088
rect 9814 3030 11395 3032
rect 6913 3027 6979 3030
rect 9673 3027 9739 3030
rect 11329 3027 11395 3030
rect 4521 2954 4587 2957
rect 11145 2954 11211 2957
rect 4521 2952 11211 2954
rect 4521 2896 4526 2952
rect 4582 2896 11150 2952
rect 11206 2896 11211 2952
rect 4521 2894 11211 2896
rect 4521 2891 4587 2894
rect 11145 2891 11211 2894
rect 1945 2818 2011 2821
rect 5349 2818 5415 2821
rect 1945 2816 5415 2818
rect 1945 2760 1950 2816
rect 2006 2760 5354 2816
rect 5410 2760 5415 2816
rect 1945 2758 5415 2760
rect 1945 2755 2011 2758
rect 5349 2755 5415 2758
rect 6729 2818 6795 2821
rect 7557 2818 7623 2821
rect 6729 2816 7623 2818
rect 6729 2760 6734 2816
rect 6790 2760 7562 2816
rect 7618 2760 7623 2816
rect 6729 2758 7623 2760
rect 6729 2755 6795 2758
rect 7557 2755 7623 2758
rect 7925 2818 7991 2821
rect 10961 2818 11027 2821
rect 7925 2816 11027 2818
rect 7925 2760 7930 2816
rect 7986 2760 10966 2816
rect 11022 2760 11027 2816
rect 7925 2758 11027 2760
rect 7925 2755 7991 2758
rect 10961 2755 11027 2758
rect 12801 2818 12867 2821
rect 14917 2818 14983 2821
rect 12801 2816 14983 2818
rect 12801 2760 12806 2816
rect 12862 2760 14922 2816
rect 14978 2760 14983 2816
rect 12801 2758 14983 2760
rect 12801 2755 12867 2758
rect 14917 2755 14983 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 8477 2682 8543 2685
rect 11237 2682 11303 2685
rect 8477 2680 11303 2682
rect 8477 2624 8482 2680
rect 8538 2624 11242 2680
rect 11298 2624 11303 2680
rect 8477 2622 11303 2624
rect 8477 2619 8543 2622
rect 11237 2619 11303 2622
rect 2497 2546 2563 2549
rect 8109 2546 8175 2549
rect 12525 2546 12591 2549
rect 2497 2544 8175 2546
rect 2497 2488 2502 2544
rect 2558 2488 8114 2544
rect 8170 2488 8175 2544
rect 2497 2486 8175 2488
rect 2497 2483 2563 2486
rect 8109 2483 8175 2486
rect 8526 2544 12591 2546
rect 8526 2488 12530 2544
rect 12586 2488 12591 2544
rect 8526 2486 12591 2488
rect 8526 2413 8586 2486
rect 12525 2483 12591 2486
rect 2773 2410 2839 2413
rect 8477 2410 8586 2413
rect 12893 2410 12959 2413
rect 2773 2408 8586 2410
rect 2773 2352 2778 2408
rect 2834 2352 8482 2408
rect 8538 2352 8586 2408
rect 2773 2350 8586 2352
rect 8710 2408 12959 2410
rect 8710 2352 12898 2408
rect 12954 2352 12959 2408
rect 8710 2350 12959 2352
rect 2773 2347 2839 2350
rect 8477 2347 8543 2350
rect 8710 2277 8770 2350
rect 12893 2347 12959 2350
rect 5257 2274 5323 2277
rect 8710 2274 8819 2277
rect 5257 2272 8819 2274
rect 5257 2216 5262 2272
rect 5318 2216 8758 2272
rect 8814 2216 8819 2272
rect 5257 2214 8819 2216
rect 5257 2211 5323 2214
rect 8753 2211 8819 2214
rect 11237 2274 11303 2277
rect 14089 2274 14155 2277
rect 11237 2272 14155 2274
rect 11237 2216 11242 2272
rect 11298 2216 14094 2272
rect 14150 2216 14155 2272
rect 11237 2214 14155 2216
rect 11237 2211 11303 2214
rect 14089 2211 14155 2214
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 8293 2002 8359 2005
rect 12985 2002 13051 2005
rect 8293 2000 13051 2002
rect 8293 1944 8298 2000
rect 8354 1944 12990 2000
rect 13046 1944 13051 2000
rect 8293 1942 13051 1944
rect 8293 1939 8359 1942
rect 12985 1939 13051 1942
rect 2405 1730 2471 1733
rect 13077 1730 13143 1733
rect 2405 1728 13143 1730
rect 2405 1672 2410 1728
rect 2466 1672 13082 1728
rect 13138 1672 13143 1728
rect 2405 1670 13143 1672
rect 2405 1667 2471 1670
rect 13077 1667 13143 1670
rect 4153 1458 4219 1461
rect 7097 1458 7163 1461
rect 4153 1456 7163 1458
rect 4153 1400 4158 1456
rect 4214 1400 7102 1456
rect 7158 1400 7163 1456
rect 4153 1398 7163 1400
rect 4153 1395 4219 1398
rect 7097 1395 7163 1398
rect 0 1186 480 1216
rect 1853 1186 1919 1189
rect 0 1184 1919 1186
rect 0 1128 1858 1184
rect 1914 1128 1919 1184
rect 0 1126 1919 1128
rect 0 1096 480 1126
rect 1853 1123 1919 1126
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 8708 27644 8772 27708
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 10180 26556 10244 26620
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 9812 22400 9876 22404
rect 9812 22344 9826 22400
rect 9826 22344 9876 22400
rect 9812 22340 9876 22344
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 10180 21856 10244 21860
rect 10180 21800 10194 21856
rect 10194 21800 10244 21856
rect 10180 21796 10244 21800
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 9812 21720 9876 21724
rect 9812 21664 9862 21720
rect 9862 21664 9876 21720
rect 9812 21660 9876 21664
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 9628 21448 9692 21452
rect 9628 21392 9642 21448
rect 9642 21392 9692 21448
rect 9628 21388 9692 21392
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 9628 20980 9692 21044
rect 8708 20768 8772 20772
rect 8708 20712 8722 20768
rect 8722 20712 8772 20768
rect 8708 20708 8772 20712
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 9812 19076 9876 19140
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 9996 18940 10060 19004
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 9812 15540 9876 15604
rect 12204 15464 12268 15468
rect 12204 15408 12254 15464
rect 12254 15408 12268 15464
rect 12204 15404 12268 15408
rect 8708 15268 8772 15332
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 9996 14996 10060 15060
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 12204 10432 12268 10436
rect 12204 10376 12254 10432
rect 12254 10376 12268 10432
rect 12204 10372 12268 10376
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 8708 10100 8772 10164
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 9444 8468 9508 8532
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 9444 3164 9508 3228
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8707 27708 8773 27709
rect 8707 27644 8708 27708
rect 8772 27644 8773 27708
rect 8707 27643 8773 27644
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 8710 20773 8770 27643
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 10179 26620 10245 26621
rect 10179 26556 10180 26620
rect 10244 26556 10245 26620
rect 10179 26555 10245 26556
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 9811 22404 9877 22405
rect 9811 22340 9812 22404
rect 9876 22340 9877 22404
rect 9811 22339 9877 22340
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8707 20772 8773 20773
rect 8707 20708 8708 20772
rect 8772 20708 8773 20772
rect 8707 20707 8773 20708
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 8944 20704 9264 21728
rect 9814 21725 9874 22339
rect 10182 21861 10242 26555
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 10179 21860 10245 21861
rect 10179 21796 10180 21860
rect 10244 21796 10245 21860
rect 10179 21795 10245 21796
rect 9811 21724 9877 21725
rect 9811 21660 9812 21724
rect 9876 21660 9877 21724
rect 9811 21659 9877 21660
rect 9627 21452 9693 21453
rect 9627 21388 9628 21452
rect 9692 21388 9693 21452
rect 9627 21387 9693 21388
rect 9630 21045 9690 21387
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 9627 21044 9693 21045
rect 9627 20980 9628 21044
rect 9692 20980 9693 21044
rect 9627 20979 9693 20980
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 9811 19140 9877 19141
rect 9811 19076 9812 19140
rect 9876 19076 9877 19140
rect 9811 19075 9877 19076
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8707 15332 8773 15333
rect 8707 15268 8708 15332
rect 8772 15268 8773 15332
rect 8707 15267 8773 15268
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 8710 10165 8770 15267
rect 8944 15264 9264 16288
rect 9814 15605 9874 19075
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 9995 19004 10061 19005
rect 9995 18940 9996 19004
rect 10060 18940 10061 19004
rect 9995 18939 10061 18940
rect 9811 15604 9877 15605
rect 9811 15540 9812 15604
rect 9876 15540 9877 15604
rect 9811 15539 9877 15540
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 9998 15061 10058 18939
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 9995 15060 10061 15061
rect 9995 14996 9996 15060
rect 10060 14996 10061 15060
rect 9995 14995 10061 14996
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8707 10164 8773 10165
rect 8707 10100 8708 10164
rect 8772 10100 8773 10164
rect 8707 10099 8773 10100
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 11610 14720 11930 15744
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 12203 15468 12269 15469
rect 12203 15404 12204 15468
rect 12268 15404 12269 15468
rect 12203 15403 12269 15404
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 12206 10437 12266 15403
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 12203 10436 12269 10437
rect 12203 10372 12204 10436
rect 12268 10372 12269 10436
rect 12203 10371 12269 10372
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 9443 8532 9509 8533
rect 9443 8468 9444 8532
rect 9508 8468 9509 8532
rect 9443 8467 9509 8468
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 9446 3229 9506 8467
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 9443 3228 9509 3229
rect 9443 3164 9444 3228
rect 9508 3164 9509 3228
rect 9443 3163 9509 3164
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _40_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_14
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_18
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_36
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_2_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_40
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l1_in_2_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_78
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_121
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_decap_8  FILLER_1_136 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_142
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_54
timestamp 1586364061
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 406 592
use scs8hd_conb_1  _22_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_9
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_13
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_37
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_41
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_45
timestamp 1586364061
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_96
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_144
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_47
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_99
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_127
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_131 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 1786 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_120
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_5_139 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_145
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_7_25
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_33
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_70
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _35_
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_78
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_145
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  mux_right_ipin_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_17
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_42
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_99
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_11
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_63
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_44
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_9
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_6
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_64
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_103
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_50
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_16_9
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_53
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_77
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 1786 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_32
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_14
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_42
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_57
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_18_100
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_8
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_3.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_31
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_40
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_124
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_19_139
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_145
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_43
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_69
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _17_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_72
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_135
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_143
timestamp 1586364061
transform 1 0 14260 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_21
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_24
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_82
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_24_57
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_75
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_96
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_114
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  mux_right_ipin_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_6
timestamp 1586364061
transform 1 0 1656 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_10
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_17
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 590 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 5244 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_43
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_55
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_29
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_38
timestamp 1586364061
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_23
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_42
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_54
timestamp 1586364061
transform 1 0 6072 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_decap_8  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_75
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_85
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_90
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_29
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_72
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_6.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_114
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_4.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_ipin_7.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_60
timestamp 1586364061
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_68
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_72
timestamp 1586364061
transform 1 0 7728 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_103
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_107
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_ipin_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_63
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_82
timestamp 1586364061
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_90
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_110
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_116
timestamp 1586364061
transform 1 0 11776 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_75
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_81
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_85
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_32_106
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_133
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_19
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2668 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_45
timestamp 1586364061
transform 1 0 5244 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_42
timestamp 1586364061
transform 1 0 4968 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_65
timestamp 1586364061
transform 1 0 7084 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_79
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_75
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_86
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_82
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_83
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_97
timestamp 1586364061
transform 1 0 10028 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10120 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_34_104
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_100
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 10948 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_118
timestamp 1586364061
transform 1 0 11960 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_115
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_122
timestamp 1586364061
transform 1 0 12328 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_133
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 1786 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_8
timestamp 1586364061
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_16
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_36
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_40
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_81
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_91
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_144
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_buf_1  mux_right_ipin_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_36_59
timestamp 1586364061
transform 1 0 6532 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6992 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_63
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_66
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_76
timestamp 1586364061
transform 1 0 8096 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_119
timestamp 1586364061
transform 1 0 12052 0 -1 22304
box -38 -48 406 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_130
timestamp 1586364061
transform 1 0 13064 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_142
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2668 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_13
timestamp 1586364061
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_26
timestamp 1586364061
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_30
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_73
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_77
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_90
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_94
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_107
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_111
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_115
timestamp 1586364061
transform 1 0 11684 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_136
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_37_140
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 590 592
use scs8hd_buf_1  mux_right_ipin_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 2668 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_14
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5704 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 5520 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_41
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_47
timestamp 1586364061
transform 1 0 5428 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_59
timestamp 1586364061
transform 1 0 6532 0 -1 23392
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_63
timestamp 1586364061
transform 1 0 6900 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_66
timestamp 1586364061
transform 1 0 7176 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_70
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9108 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_82
timestamp 1586364061
transform 1 0 8648 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_86
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_89
timestamp 1586364061
transform 1 0 9292 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_112
timestamp 1586364061
transform 1 0 11408 0 -1 23392
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12144 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 13156 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_133
timestamp 1586364061
transform 1 0 13340 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_11
timestamp 1586364061
transform 1 0 2116 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 2668 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2300 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_31
timestamp 1586364061
transform 1 0 3956 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_42
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_52
timestamp 1586364061
transform 1 0 5888 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_53
timestamp 1586364061
transform 1 0 5980 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_64
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_61
timestamp 1586364061
transform 1 0 6716 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_77
timestamp 1586364061
transform 1 0 8188 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_79
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8372 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_ipin_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9108 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_83
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_81
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_3  FILLER_40_89
timestamp 1586364061
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_106
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 11040 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_110
timestamp 1586364061
transform 1 0 11224 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11316 0 -1 24480
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_130
timestamp 1586364061
transform 1 0 13064 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_142
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_10.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 2116 0 1 24480
box -38 -48 1786 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_7
timestamp 1586364061
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4600 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_30
timestamp 1586364061
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_34
timestamp 1586364061
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5612 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_47
timestamp 1586364061
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_55
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_ipin_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_41_70
timestamp 1586364061
transform 1 0 7544 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_92
timestamp 1586364061
transform 1 0 9568 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_104
timestamp 1586364061
transform 1 0 10672 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_41_116
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2300 0 -1 25568
box -38 -48 866 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_10.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 2116 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 774 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 4140 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 4600 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_22
timestamp 1586364061
transform 1 0 3128 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_30
timestamp 1586364061
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_36
timestamp 1586364061
transform 1 0 4416 0 -1 25568
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_42_40
timestamp 1586364061
transform 1 0 4784 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7820 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_71
timestamp 1586364061
transform 1 0 7636 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 10120 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_83
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_97
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_100
timestamp 1586364061
transform 1 0 10304 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_112
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_124
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_136
timestamp 1586364061
transform 1 0 13616 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_144
timestamp 1586364061
transform 1 0 14352 0 -1 25568
box -38 -48 222 592
use scs8hd_buf_1  mux_right_ipin_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_6
timestamp 1586364061
transform 1 0 1656 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_10
timestamp 1586364061
transform 1 0 2024 0 1 25568
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4508 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4324 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 3956 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_22
timestamp 1586364061
transform 1 0 3128 0 1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_43_30
timestamp 1586364061
transform 1 0 3864 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_33
timestamp 1586364061
transform 1 0 4140 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_46
timestamp 1586364061
transform 1 0 5336 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_50
timestamp 1586364061
transform 1 0 5704 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_53
timestamp 1586364061
transform 1 0 5980 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_57
timestamp 1586364061
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8372 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_71
timestamp 1586364061
transform 1 0 7636 0 1 25568
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1586364061
transform 1 0 8556 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 9936 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9568 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_90
timestamp 1586364061
transform 1 0 9384 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_94
timestamp 1586364061
transform 1 0 9752 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11132 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11500 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_107
timestamp 1586364061
transform 1 0 10948 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_111
timestamp 1586364061
transform 1 0 11316 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_115
timestamp 1586364061
transform 1 0 11684 0 1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_43_121
timestamp 1586364061
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2576 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_18
timestamp 1586364061
transform 1 0 2760 0 -1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4508 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2944 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_22
timestamp 1586364061
transform 1 0 3128 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_30
timestamp 1586364061
transform 1 0 3864 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_36
timestamp 1586364061
transform 1 0 4416 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_6  FILLER_44_39
timestamp 1586364061
transform 1 0 4692 0 -1 26656
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1586364061
transform 1 0 5888 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 5704 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 5336 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_45
timestamp 1586364061
transform 1 0 5244 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_48
timestamp 1586364061
transform 1 0 5520 0 -1 26656
box -38 -48 222 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 7452 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 6900 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7912 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_61
timestamp 1586364061
transform 1 0 6716 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_65
timestamp 1586364061
transform 1 0 7084 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_44_72
timestamp 1586364061
transform 1 0 7728 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_76
timestamp 1586364061
transform 1 0 8096 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_4  FILLER_44_83
timestamp 1586364061
transform 1 0 8740 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_87
timestamp 1586364061
transform 1 0 9108 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_90
timestamp 1586364061
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 9936 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_99
timestamp 1586364061
transform 1 0 10212 0 -1 26656
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10948 0 -1 26656
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 10396 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_103
timestamp 1586364061
transform 1 0 10580 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 12880 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_126
timestamp 1586364061
transform 1 0 12696 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_130
timestamp 1586364061
transform 1 0 13064 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_44_142
timestamp 1586364061
transform 1 0 14168 0 -1 26656
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2576 0 1 26656
box -38 -48 1786 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2392 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2024 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 1656 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_8
timestamp 1586364061
transform 1 0 1840 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_12
timestamp 1586364061
transform 1 0 2208 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4508 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_35
timestamp 1586364061
transform 1 0 4324 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4876 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_43
timestamp 1586364061
transform 1 0 5060 0 1 26656
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_71
timestamp 1586364061
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_75
timestamp 1586364061
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_79
timestamp 1586364061
transform 1 0 8372 0 1 26656
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8648 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_84
timestamp 1586364061
transform 1 0 8832 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_97
timestamp 1586364061
transform 1 0 10028 0 1 26656
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1586364061
transform 1 0 10764 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 10580 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_101
timestamp 1586364061
transform 1 0 10396 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_114
timestamp 1586364061
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_118
timestamp 1586364061
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 13432 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_132
timestamp 1586364061
transform 1 0 13248 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_136
timestamp 1586364061
transform 1 0 13616 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_144
timestamp 1586364061
transform 1 0 14352 0 1 26656
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2852 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_3  FILLER_46_11
timestamp 1586364061
transform 1 0 2116 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_17
timestamp 1586364061
transform 1 0 2668 0 1 27744
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3036 0 1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 4508 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_23
timestamp 1586364061
transform 1 0 3220 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_6  FILLER_47_30
timestamp 1586364061
transform 1 0 3864 0 1 27744
box -38 -48 590 592
use scs8hd_fill_1  FILLER_47_36
timestamp 1586364061
transform 1 0 4416 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_47
timestamp 1586364061
transform 1 0 5428 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_43
timestamp 1586364061
transform 1 0 5060 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 5244 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 4876 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_54
timestamp 1586364061
transform 1 0 6072 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_46_51
timestamp 1586364061
transform 1 0 5796 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5888 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6256 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_58
timestamp 1586364061
transform 1 0 6440 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_46_59
timestamp 1586364061
transform 1 0 6532 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_69
timestamp 1586364061
transform 1 0 7452 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_66
timestamp 1586364061
transform 1 0 7176 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 406 592
use scs8hd_decap_6  FILLER_46_64
timestamp 1586364061
transform 1 0 6992 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 6808 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7268 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_6  FILLER_46_79
timestamp 1586364061
transform 1 0 8372 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7636 0 1 27744
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7544 0 -1 27744
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7820 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_82
timestamp 1586364061
transform 1 0 8648 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_88
timestamp 1586364061
transform 1 0 9200 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_85
timestamp 1586364061
transform 1 0 8924 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8832 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 9200 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_47_99
timestamp 1586364061
transform 1 0 10212 0 1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9384 0 1 27744
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10948 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11316 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11684 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_107
timestamp 1586364061
transform 1 0 10948 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_109
timestamp 1586364061
transform 1 0 11132 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_47_113
timestamp 1586364061
transform 1 0 11500 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_46_136
timestamp 1586364061
transform 1 0 13616 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_1  FILLER_47_121
timestamp 1586364061
transform 1 0 12236 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_46_144
timestamp 1586364061
transform 1 0 14352 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1586364061
transform 1 0 4508 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3036 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_23
timestamp 1586364061
transform 1 0 3220 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_4  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_36
timestamp 1586364061
transform 1 0 4416 0 -1 28832
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 5520 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_46
timestamp 1586364061
transform 1 0 5336 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_50
timestamp 1586364061
transform 1 0 5704 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_54
timestamp 1586364061
transform 1 0 6072 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8280 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_75
timestamp 1586364061
transform 1 0 8004 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8648 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10212 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_48_84
timestamp 1586364061
transform 1 0 8832 0 -1 28832
box -38 -48 590 592
use scs8hd_decap_6  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10948 0 -1 28832
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_101
timestamp 1586364061
transform 1 0 10396 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_126
timestamp 1586364061
transform 1 0 12696 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_138
timestamp 1586364061
transform 1 0 13800 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2208 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_6
timestamp 1586364061
transform 1 0 1656 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_10
timestamp 1586364061
transform 1 0 2024 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_14
timestamp 1586364061
transform 1 0 2392 0 1 28832
box -38 -48 1142 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 4048 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 4508 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_26
timestamp 1586364061
transform 1 0 3496 0 1 28832
box -38 -48 590 592
use scs8hd_fill_2  FILLER_49_35
timestamp 1586364061
transform 1 0 4324 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1586364061
transform 1 0 5060 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 4876 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6072 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_52
timestamp 1586364061
transform 1 0 5888 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_56
timestamp 1586364061
transform 1 0 6256 0 1 28832
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8280 0 1 28832
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7728 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8096 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7360 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_60
timestamp 1586364061
transform 1 0 6624 0 1 28832
box -38 -48 130 592
use scs8hd_decap_6  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 590 592
use scs8hd_fill_2  FILLER_49_70
timestamp 1586364061
transform 1 0 7544 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10212 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_97
timestamp 1586364061
transform 1 0 10028 0 1 28832
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_101
timestamp 1586364061
transform 1 0 10396 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_114
timestamp 1586364061
transform 1 0 11592 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_118
timestamp 1586364061
transform 1 0 11960 0 1 28832
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 2852 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2392 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_6
timestamp 1586364061
transform 1 0 1656 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  FILLER_50_16
timestamp 1586364061
transform 1 0 2576 0 -1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 4232 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 3220 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_21
timestamp 1586364061
transform 1 0 3036 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_25
timestamp 1586364061
transform 1 0 3404 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_2  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_36
timestamp 1586364061
transform 1 0 4416 0 -1 29920
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 4876 0 -1 29920
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_50_40
timestamp 1586364061
transform 1 0 4784 0 -1 29920
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7728 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6808 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7176 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 7544 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_60
timestamp 1586364061
transform 1 0 6624 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_64
timestamp 1586364061
transform 1 0 6992 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_ipin_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10212 0 -1 29920
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8740 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_81
timestamp 1586364061
transform 1 0 8556 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_85
timestamp 1586364061
transform 1 0 8924 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_91
timestamp 1586364061
transform 1 0 9476 0 -1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_97
timestamp 1586364061
transform 1 0 10028 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_118
timestamp 1586364061
transform 1 0 11960 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_130
timestamp 1586364061
transform 1 0 13064 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_50_142
timestamp 1586364061
transform 1 0 14168 0 -1 29920
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1586364061
transform 1 0 2852 0 1 29920
box -38 -48 866 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2392 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2024 0 1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_51_9
timestamp 1586364061
transform 1 0 1932 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_12
timestamp 1586364061
transform 1 0 2208 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_16
timestamp 1586364061
transform 1 0 2576 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 4048 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 4416 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_28
timestamp 1586364061
transform 1 0 3680 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_34
timestamp 1586364061
transform 1 0 4232 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_38
timestamp 1586364061
transform 1 0 4600 0 1 29920
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_53
timestamp 1586364061
transform 1 0 5980 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_57
timestamp 1586364061
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8280 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_71
timestamp 1586364061
transform 1 0 7636 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_76
timestamp 1586364061
transform 1 0 8096 0 1 29920
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9568 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8648 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_80
timestamp 1586364061
transform 1 0 8464 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_84
timestamp 1586364061
transform 1 0 8832 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_88
timestamp 1586364061
transform 1 0 9200 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 10580 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 11500 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 10948 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 11868 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_101
timestamp 1586364061
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_105
timestamp 1586364061
transform 1 0 10764 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_109
timestamp 1586364061
transform 1 0 11132 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_115
timestamp 1586364061
transform 1 0 11684 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_119
timestamp 1586364061
transform 1 0 12052 0 1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_8  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 774 592
use scs8hd_decap_8  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_16
timestamp 1586364061
transform 1 0 2576 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_11
timestamp 1586364061
transform 1 0 2116 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_52_11
timestamp 1586364061
transform 1 0 2116 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2760 0 1 31008
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_29
timestamp 1586364061
transform 1 0 3772 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_23
timestamp 1586364061
transform 1 0 3220 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2944 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_33
timestamp 1586364061
transform 1 0 4140 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3956 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1586364061
transform 1 0 4508 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_46
timestamp 1586364061
transform 1 0 5336 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_49
timestamp 1586364061
transform 1 0 5612 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_45
timestamp 1586364061
transform 1 0 5244 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_41
timestamp 1586364061
transform 1 0 4876 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 5060 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 5520 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_58
timestamp 1586364061
transform 1 0 6440 0 1 31008
box -38 -48 314 592
use scs8hd_decap_8  FILLER_53_50
timestamp 1586364061
transform 1 0 5704 0 1 31008
box -38 -48 774 592
use scs8hd_decap_4  FILLER_52_53
timestamp 1586364061
transform 1 0 5980 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5796 0 -1 31008
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6348 0 -1 31008
box -38 -48 866 592
use scs8hd_decap_6  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 590 592
use scs8hd_fill_2  FILLER_52_66
timestamp 1586364061
transform 1 0 7176 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_6  FILLER_53_78
timestamp 1586364061
transform 1 0 8280 0 1 31008
box -38 -48 590 592
use scs8hd_fill_2  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_70
timestamp 1586364061
transform 1 0 7544 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_70
timestamp 1586364061
transform 1 0 7544 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8096 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 7728 0 1 31008
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7912 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_1  FILLER_53_84
timestamp 1586364061
transform 1 0 8832 0 1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_52_89
timestamp 1586364061
transform 1 0 9292 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_52_83
timestamp 1586364061
transform 1 0 8740 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 9108 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 8924 0 1 31008
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1586364061
transform 1 0 9108 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_96
timestamp 1586364061
transform 1 0 9936 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 11500 0 -1 31008
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10856 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_102
timestamp 1586364061
transform 1 0 10488 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_3  FILLER_52_110
timestamp 1586364061
transform 1 0 11224 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_100
timestamp 1586364061
transform 1 0 10304 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_104
timestamp 1586364061
transform 1 0 10672 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_108
timestamp 1586364061
transform 1 0 11040 0 1 31008
box -38 -48 1142 592
use scs8hd_buf_1  mux_left_ipin_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_132
timestamp 1586364061
transform 1 0 13248 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_120
timestamp 1586364061
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_138
timestamp 1586364061
transform 1 0 13800 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13984 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_144
timestamp 1586364061
transform 1 0 14352 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_142
timestamp 1586364061
transform 1 0 14168 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_19
timestamp 1586364061
transform 1 0 2852 0 -1 32096
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 2944 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_22
timestamp 1586364061
transform 1 0 3128 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_1  FILLER_54_30
timestamp 1586364061
transform 1 0 3864 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5980 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6348 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_51
timestamp 1586364061
transform 1 0 5796 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_55
timestamp 1586364061
transform 1 0 6164 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_59
timestamp 1586364061
transform 1 0 6532 0 -1 32096
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7084 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 6716 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_63
timestamp 1586364061
transform 1 0 6900 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_67
timestamp 1586364061
transform 1 0 7268 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_77
timestamp 1586364061
transform 1 0 8188 0 -1 32096
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10120 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 9108 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 9936 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_85
timestamp 1586364061
transform 1 0 8924 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_89
timestamp 1586364061
transform 1 0 9292 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 11132 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_107
timestamp 1586364061
transform 1 0 10948 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_111
timestamp 1586364061
transform 1 0 11316 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_115
timestamp 1586364061
transform 1 0 11684 0 -1 32096
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 12328 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_121
timestamp 1586364061
transform 1 0 12236 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_124
timestamp 1586364061
transform 1 0 12512 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_54_136
timestamp 1586364061
transform 1 0 13616 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_54_144
timestamp 1586364061
transform 1 0 14352 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_7
timestamp 1586364061
transform 1 0 1748 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_19
timestamp 1586364061
transform 1 0 2852 0 1 32096
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4232 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_31
timestamp 1586364061
transform 1 0 3956 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_36
timestamp 1586364061
transform 1 0 4416 0 1 32096
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_40
timestamp 1586364061
transform 1 0 4784 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1586364061
transform 1 0 7452 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7084 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_67
timestamp 1586364061
transform 1 0 7268 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_78
timestamp 1586364061
transform 1 0 8280 0 1 32096
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10212 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 8464 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 8832 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_82
timestamp 1586364061
transform 1 0 8648 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_95
timestamp 1586364061
transform 1 0 9844 0 1 32096
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 10580 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_101
timestamp 1586364061
transform 1 0 10396 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_114
timestamp 1586364061
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_118
timestamp 1586364061
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 12880 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_126
timestamp 1586364061
transform 1 0 12696 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_130
timestamp 1586364061
transform 1 0 13064 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_55_142
timestamp 1586364061
transform 1 0 14168 0 1 32096
box -38 -48 406 592
use scs8hd_buf_1  mux_right_ipin_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_6
timestamp 1586364061
transform 1 0 1656 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_18
timestamp 1586364061
transform 1 0 2760 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_30
timestamp 1586364061
transform 1 0 3864 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_36
timestamp 1586364061
transform 1 0 4416 0 -1 33184
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5520 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_46
timestamp 1586364061
transform 1 0 5336 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_57
timestamp 1586364061
transform 1 0 6348 0 -1 33184
box -38 -48 590 592
use scs8hd_mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7084 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8096 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 6900 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_74
timestamp 1586364061
transform 1 0 7912 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_78
timestamp 1586364061
transform 1 0 8280 0 -1 33184
box -38 -48 774 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 9016 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_88
timestamp 1586364061
transform 1 0 9200 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_96
timestamp 1586364061
transform 1 0 9936 0 -1 33184
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10304 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_102
timestamp 1586364061
transform 1 0 10488 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_114
timestamp 1586364061
transform 1 0 11592 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_119
timestamp 1586364061
transform 1 0 12052 0 -1 33184
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1586364061
transform 1 0 12328 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_12  FILLER_56_131
timestamp 1586364061
transform 1 0 13156 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_143
timestamp 1586364061
transform 1 0 14260 0 -1 33184
box -38 -48 314 592
use scs8hd_buf_1  mux_right_ipin_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 1840 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 2852 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2208 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_6
timestamp 1586364061
transform 1 0 1656 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_10
timestamp 1586364061
transform 1 0 2024 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_14
timestamp 1586364061
transform 1 0 2392 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_18
timestamp 1586364061
transform 1 0 2760 0 1 33184
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 33184
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 4048 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3680 0 1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_57_21
timestamp 1586364061
transform 1 0 3036 0 1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_30
timestamp 1586364061
transform 1 0 3864 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6256 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_53
timestamp 1586364061
transform 1 0 5980 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_58
timestamp 1586364061
transform 1 0 6440 0 1 33184
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7636 0 1 33184
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7452 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_66
timestamp 1586364061
transform 1 0 7176 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_90
timestamp 1586364061
transform 1 0 9384 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_96
timestamp 1586364061
transform 1 0 9936 0 1 33184
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11868 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_100
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_113
timestamp 1586364061
transform 1 0 11500 0 1 33184
box -38 -48 406 592
use scs8hd_decap_3  FILLER_57_119
timestamp 1586364061
transform 1 0 12052 0 1 33184
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 13800 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_132
timestamp 1586364061
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_136
timestamp 1586364061
transform 1 0 13616 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 14168 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_140
timestamp 1586364061
transform 1 0 13984 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_144
timestamp 1586364061
transform 1 0 14352 0 1 33184
box -38 -48 222 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 2852 0 -1 34272
box -38 -48 406 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 1748 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 1564 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_11
timestamp 1586364061
transform 1 0 2116 0 -1 34272
box -38 -48 774 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 4600 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 3404 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_23
timestamp 1586364061
transform 1 0 3220 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_36
timestamp 1586364061
transform 1 0 4416 0 -1 34272
box -38 -48 222 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_58_40
timestamp 1586364061
transform 1 0 4784 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_58_48
timestamp 1586364061
transform 1 0 5520 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_58_75
timestamp 1586364061
transform 1 0 8004 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9844 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_87
timestamp 1586364061
transform 1 0 9108 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_97
timestamp 1586364061
transform 1 0 10028 0 -1 34272
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10304 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11316 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_109
timestamp 1586364061
transform 1 0 11132 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_113
timestamp 1586364061
transform 1 0 11500 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_136
timestamp 1586364061
transform 1 0 13616 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_144
timestamp 1586364061
transform 1 0 14352 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_7
timestamp 1586364061
transform 1 0 1748 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_7
timestamp 1586364061
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_6  FILLER_59_17
timestamp 1586364061
transform 1 0 2668 0 1 34272
box -38 -48 590 592
use scs8hd_decap_4  FILLER_59_11
timestamp 1586364061
transform 1 0 2116 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 222 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_19
timestamp 1586364061
transform 1 0 2852 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 4508 0 -1 35360
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_11.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 3404 0 1 34272
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_11.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 3220 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_36
timestamp 1586364061
transform 1 0 4416 0 -1 35360
box -38 -48 130 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 5612 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 5612 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_44
timestamp 1586364061
transform 1 0 5152 0 1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_59_48
timestamp 1586364061
transform 1 0 5520 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_decap_8  FILLER_60_41
timestamp 1586364061
transform 1 0 4876 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_53
timestamp 1586364061
transform 1 0 5980 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_ipin_13.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 7360 0 1 34272
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_13.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 7912 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 406 592
use scs8hd_decap_3  FILLER_60_65
timestamp 1586364061
transform 1 0 7084 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_72
timestamp 1586364061
transform 1 0 7728 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_76
timestamp 1586364061
transform 1 0 8096 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_6  FILLER_60_84
timestamp 1586364061
transform 1 0 8832 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_87
timestamp 1586364061
transform 1 0 9108 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 9292 0 1 34272
box -38 -48 222 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_91
timestamp 1586364061
transform 1 0 9476 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9384 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_ipin_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_114
timestamp 1586364061
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_118
timestamp 1586364061
transform 1 0 11960 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_112
timestamp 1586364061
transform 1 0 11408 0 -1 35360
box -38 -48 774 592
use scs8hd_mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 12420 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_132
timestamp 1586364061
transform 1 0 13248 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_60_120
timestamp 1586364061
transform 1 0 12144 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_60_125
timestamp 1586364061
transform 1 0 12604 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_60_137
timestamp 1586364061
transform 1 0 13708 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_144
timestamp 1586364061
transform 1 0 14352 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_buf_1  mux_right_ipin_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1840 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_6
timestamp 1586364061
transform 1 0 1656 0 1 35360
box -38 -48 222 592
use scs8hd_decap_8  FILLER_61_10
timestamp 1586364061
transform 1 0 2024 0 1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_61_18
timestamp 1586364061
transform 1 0 2760 0 1 35360
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 4048 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 2944 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 3496 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 4600 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_24
timestamp 1586364061
transform 1 0 3312 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_28
timestamp 1586364061
transform 1 0 3680 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_36
timestamp 1586364061
transform 1 0 4416 0 1 35360
box -38 -48 222 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 5612 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 5428 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 6164 0 1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_61_40
timestamp 1586364061
transform 1 0 4784 0 1 35360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_61_46
timestamp 1586364061
transform 1 0 5336 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_53
timestamp 1586364061
transform 1 0 5980 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_57
timestamp 1586364061
transform 1 0 6348 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 7360 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_66
timestamp 1586364061
transform 1 0 7176 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_70
timestamp 1586364061
transform 1 0 7544 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_78
timestamp 1586364061
transform 1 0 8280 0 1 35360
box -38 -48 222 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 9660 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 8464 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 9476 0 1 35360
box -38 -48 222 592
use scs8hd_decap_8  FILLER_61_82
timestamp 1586364061
transform 1 0 8648 0 1 35360
box -38 -48 774 592
use scs8hd_fill_1  FILLER_61_90
timestamp 1586364061
transform 1 0 9384 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_97
timestamp 1586364061
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_101
timestamp 1586364061
transform 1 0 10396 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_113
timestamp 1586364061
transform 1 0 11500 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_fill_1  FILLER_61_121
timestamp 1586364061
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 5428 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_3  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_51
timestamp 1586364061
transform 1 0 5796 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_63
timestamp 1586364061
transform 1 0 6900 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_75
timestamp 1586364061
transform 1 0 8004 0 -1 36448
box -38 -48 1142 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_87
timestamp 1586364061
transform 1 0 9108 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_91
timestamp 1586364061
transform 1 0 9476 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_97
timestamp 1586364061
transform 1 0 10028 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_109
timestamp 1586364061
transform 1 0 11132 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_121
timestamp 1586364061
transform 1 0 12236 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_133
timestamp 1586364061
transform 1 0 13340 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 590 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 5244 0 1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_49
timestamp 1586364061
transform 1 0 5612 0 1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_63_53
timestamp 1586364061
transform 1 0 5980 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 1096 480 1216 6 ccff_head
port 0 nsew default input
rlabel metal3 s 15520 20000 16000 20120 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 left_grid_pin_0_
port 82 nsew default tristate
rlabel metal3 s 0 26936 480 27056 6 left_grid_pin_10_
port 83 nsew default tristate
rlabel metal3 s 0 29248 480 29368 6 left_grid_pin_11_
port 84 nsew default tristate
rlabel metal3 s 0 31560 480 31680 6 left_grid_pin_12_
port 85 nsew default tristate
rlabel metal3 s 0 34008 480 34128 6 left_grid_pin_13_
port 86 nsew default tristate
rlabel metal3 s 0 36320 480 36440 6 left_grid_pin_14_
port 87 nsew default tristate
rlabel metal3 s 0 38632 480 38752 6 left_grid_pin_15_
port 88 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 left_grid_pin_1_
port 89 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 left_grid_pin_2_
port 90 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 left_grid_pin_3_
port 91 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 left_grid_pin_4_
port 92 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 left_grid_pin_5_
port 93 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 left_grid_pin_6_
port 94 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 left_grid_pin_7_
port 95 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 left_grid_pin_8_
port 96 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 left_grid_pin_9_
port 97 nsew default tristate
rlabel metal3 s 15520 6672 16000 6792 6 prog_clk
port 98 nsew default input
rlabel metal3 s 15520 33328 16000 33448 6 right_grid_pin_52_
port 99 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 100 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
