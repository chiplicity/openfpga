magic
tech EFS8A
magscale 1 2
timestamp 1602873894
<< locali >>
rect 6187 34153 6193 34187
rect 10051 34153 10057 34187
rect 6187 34085 6221 34153
rect 10051 34085 10085 34153
rect 4019 31841 4146 31875
rect 8527 31841 8654 31875
rect 11287 31841 11322 31875
rect 10051 30889 10057 30923
rect 10051 30821 10085 30889
rect 8815 30345 8953 30379
rect 7147 30073 7192 30107
rect 2881 29665 3042 29699
rect 12299 29665 12334 29699
rect 2881 29631 2915 29665
rect 13311 28577 13346 28611
rect 13127 27489 13162 27523
rect 9045 25687 9079 25993
rect 10051 25449 10057 25483
rect 10051 25381 10085 25449
rect 12391 22525 12518 22559
rect 9407 22423 9441 22491
rect 9407 22389 9413 22423
rect 5359 22185 5365 22219
rect 5359 22117 5393 22185
rect 10051 21097 10057 21131
rect 10051 21029 10085 21097
rect 12391 20349 12518 20383
rect 7113 19771 7147 19873
rect 7573 18071 7607 18173
rect 9775 18071 9809 18139
rect 9775 18037 9781 18071
rect 5267 17833 5273 17867
rect 5267 17765 5301 17833
rect 10051 15657 10057 15691
rect 10051 15589 10085 15657
rect 13035 15521 13070 15555
rect 4939 14433 5066 14467
rect 5267 13719 5301 13787
rect 5267 13685 5273 13719
rect 7975 13413 8020 13447
rect 4813 12257 4974 12291
rect 4813 12087 4847 12257
rect 4387 8993 4422 9027
rect 9505 8415 9539 8585
rect 8119 6953 8125 6987
rect 8119 6885 8153 6953
rect 6377 5151 6411 5321
rect 8493 5083 8527 5253
rect 11161 2907 11195 3077
rect 4399 2601 4537 2635
<< viali >>
rect 8125 37077 8159 37111
rect 10977 36873 11011 36907
rect 6964 36669 6998 36703
rect 7941 36669 7975 36703
rect 8033 36669 8067 36703
rect 8585 36669 8619 36703
rect 10793 36669 10827 36703
rect 7389 36601 7423 36635
rect 7067 36533 7101 36567
rect 8309 36533 8343 36567
rect 11345 36533 11379 36567
rect 9873 36329 9907 36363
rect 11437 36329 11471 36363
rect 7297 36261 7331 36295
rect 9689 36193 9723 36227
rect 11253 36193 11287 36227
rect 7205 36125 7239 36159
rect 7757 36057 7791 36091
rect 8769 35989 8803 36023
rect 8125 35785 8159 35819
rect 10425 35785 10459 35819
rect 11483 35785 11517 35819
rect 12633 35785 12667 35819
rect 7757 35717 7791 35751
rect 8585 35581 8619 35615
rect 8677 35581 8711 35615
rect 9229 35581 9263 35615
rect 10241 35581 10275 35615
rect 10793 35581 10827 35615
rect 11412 35581 11446 35615
rect 12449 35581 12483 35615
rect 13001 35581 13035 35615
rect 6285 35513 6319 35547
rect 7205 35513 7239 35547
rect 7297 35513 7331 35547
rect 6653 35445 6687 35479
rect 8769 35445 8803 35479
rect 9781 35445 9815 35479
rect 11805 35445 11839 35479
rect 12173 35445 12207 35479
rect 11713 35241 11747 35275
rect 12909 35241 12943 35275
rect 7021 35173 7055 35207
rect 9965 35173 9999 35207
rect 5892 35105 5926 35139
rect 8620 35105 8654 35139
rect 11529 35105 11563 35139
rect 12725 35105 12759 35139
rect 6929 35037 6963 35071
rect 7573 35037 7607 35071
rect 8723 35037 8757 35071
rect 9873 35037 9907 35071
rect 10517 35037 10551 35071
rect 5963 34969 5997 35003
rect 6653 34969 6687 35003
rect 5273 34901 5307 34935
rect 7849 34901 7883 34935
rect 10885 34901 10919 34935
rect 6193 34697 6227 34731
rect 7757 34697 7791 34731
rect 8585 34697 8619 34731
rect 13645 34697 13679 34731
rect 4307 34629 4341 34663
rect 5089 34561 5123 34595
rect 8217 34561 8251 34595
rect 8677 34561 8711 34595
rect 10517 34561 10551 34595
rect 10977 34561 11011 34595
rect 12909 34561 12943 34595
rect 13277 34561 13311 34595
rect 4236 34493 4270 34527
rect 4629 34493 4663 34527
rect 5181 34493 5215 34527
rect 5641 34493 5675 34527
rect 5917 34493 5951 34527
rect 6837 34493 6871 34527
rect 12484 34493 12518 34527
rect 13461 34493 13495 34527
rect 14013 34493 14047 34527
rect 6653 34425 6687 34459
rect 7199 34425 7233 34459
rect 9039 34425 9073 34459
rect 10609 34425 10643 34459
rect 11621 34425 11655 34459
rect 9597 34357 9631 34391
rect 9873 34357 9907 34391
rect 10333 34357 10367 34391
rect 12587 34357 12621 34391
rect 5365 34153 5399 34187
rect 6193 34153 6227 34187
rect 6745 34153 6779 34187
rect 7021 34153 7055 34187
rect 7389 34153 7423 34187
rect 9413 34153 9447 34187
rect 10057 34153 10091 34187
rect 10609 34153 10643 34187
rect 13553 34153 13587 34187
rect 7757 34085 7791 34119
rect 11529 34085 11563 34119
rect 11621 34085 11655 34119
rect 4848 34017 4882 34051
rect 13369 34017 13403 34051
rect 5825 33949 5859 33983
rect 7665 33949 7699 33983
rect 7941 33949 7975 33983
rect 9689 33949 9723 33983
rect 4951 33881 4985 33915
rect 12081 33881 12115 33915
rect 5641 33813 5675 33847
rect 8677 33813 8711 33847
rect 10885 33813 10919 33847
rect 12541 33813 12575 33847
rect 6285 33609 6319 33643
rect 7849 33609 7883 33643
rect 8309 33609 8343 33643
rect 10057 33609 10091 33643
rect 10425 33609 10459 33643
rect 11713 33609 11747 33643
rect 9689 33541 9723 33575
rect 4353 33473 4387 33507
rect 5917 33473 5951 33507
rect 6561 33473 6595 33507
rect 7573 33473 7607 33507
rect 8769 33473 8803 33507
rect 12541 33473 12575 33507
rect 12817 33473 12851 33507
rect 3525 33405 3559 33439
rect 3617 33405 3651 33439
rect 4077 33405 4111 33439
rect 5181 33405 5215 33439
rect 5641 33405 5675 33439
rect 10517 33405 10551 33439
rect 6929 33337 6963 33371
rect 7021 33337 7055 33371
rect 8677 33337 8711 33371
rect 9131 33337 9165 33371
rect 10838 33337 10872 33371
rect 12265 33337 12299 33371
rect 12633 33337 12667 33371
rect 4813 33269 4847 33303
rect 11437 33269 11471 33303
rect 13553 33269 13587 33303
rect 3709 33065 3743 33099
rect 4859 33065 4893 33099
rect 8861 33065 8895 33099
rect 11529 33065 11563 33099
rect 6095 32997 6129 33031
rect 8033 32997 8067 33031
rect 10333 32997 10367 33031
rect 10885 32997 10919 33031
rect 11897 32997 11931 33031
rect 12449 32997 12483 33031
rect 4788 32929 4822 32963
rect 13344 32929 13378 32963
rect 5273 32861 5307 32895
rect 5733 32861 5767 32895
rect 7941 32861 7975 32895
rect 8217 32861 8251 32895
rect 10241 32861 10275 32895
rect 11805 32861 11839 32895
rect 5641 32725 5675 32759
rect 6653 32725 6687 32759
rect 7021 32725 7055 32759
rect 7389 32725 7423 32759
rect 9965 32725 9999 32759
rect 13415 32725 13449 32759
rect 8309 32521 8343 32555
rect 8585 32521 8619 32555
rect 9873 32521 9907 32555
rect 10977 32521 11011 32555
rect 11713 32521 11747 32555
rect 12081 32521 12115 32555
rect 12587 32521 12621 32555
rect 5089 32453 5123 32487
rect 11345 32453 11379 32487
rect 6561 32385 6595 32419
rect 9505 32385 9539 32419
rect 10057 32385 10091 32419
rect 10701 32385 10735 32419
rect 4236 32317 4270 32351
rect 4629 32317 4663 32351
rect 5457 32317 5491 32351
rect 5733 32317 5767 32351
rect 7389 32317 7423 32351
rect 12484 32317 12518 32351
rect 12909 32317 12943 32351
rect 5917 32249 5951 32283
rect 7710 32249 7744 32283
rect 10149 32249 10183 32283
rect 4307 32181 4341 32215
rect 6285 32181 6319 32215
rect 7205 32181 7239 32215
rect 13369 32181 13403 32215
rect 6285 31977 6319 32011
rect 8217 31977 8251 32011
rect 8723 31977 8757 32011
rect 9965 31977 9999 32011
rect 11391 31977 11425 32011
rect 4215 31909 4249 31943
rect 6009 31909 6043 31943
rect 7021 31909 7055 31943
rect 7573 31909 7607 31943
rect 7849 31909 7883 31943
rect 3985 31841 4019 31875
rect 5549 31841 5583 31875
rect 5825 31841 5859 31875
rect 8493 31841 8527 31875
rect 9689 31841 9723 31875
rect 10149 31841 10183 31875
rect 11253 31841 11287 31875
rect 6929 31773 6963 31807
rect 9045 31637 9079 31671
rect 10793 31637 10827 31671
rect 6561 31433 6595 31467
rect 7021 31433 7055 31467
rect 10425 31433 10459 31467
rect 7573 31297 7607 31331
rect 8217 31297 8251 31331
rect 10793 31297 10827 31331
rect 11437 31297 11471 31331
rect 4537 31229 4571 31263
rect 5273 31229 5307 31263
rect 9045 31229 9079 31263
rect 9505 31229 9539 31263
rect 10057 31229 10091 31263
rect 4169 31161 4203 31195
rect 5733 31161 5767 31195
rect 7665 31161 7699 31195
rect 9781 31161 9815 31195
rect 10885 31161 10919 31195
rect 4905 31093 4939 31127
rect 6101 31093 6135 31127
rect 8677 31093 8711 31127
rect 11713 31093 11747 31127
rect 10057 30889 10091 30923
rect 10609 30889 10643 30923
rect 10977 30889 11011 30923
rect 4813 30821 4847 30855
rect 7849 30821 7883 30855
rect 11621 30821 11655 30855
rect 12173 30821 12207 30855
rect 6285 30753 6319 30787
rect 6469 30753 6503 30787
rect 4721 30685 4755 30719
rect 5365 30685 5399 30719
rect 7757 30685 7791 30719
rect 8217 30685 8251 30719
rect 8677 30685 8711 30719
rect 9689 30685 9723 30719
rect 11529 30685 11563 30719
rect 9045 30617 9079 30651
rect 5733 30549 5767 30583
rect 6561 30549 6595 30583
rect 7113 30549 7147 30583
rect 7573 30549 7607 30583
rect 3893 30345 3927 30379
rect 4721 30345 4755 30379
rect 7757 30345 7791 30379
rect 8033 30345 8067 30379
rect 8953 30345 8987 30379
rect 10885 30345 10919 30379
rect 11529 30345 11563 30379
rect 10609 30277 10643 30311
rect 11805 30277 11839 30311
rect 3985 30209 4019 30243
rect 5365 30209 5399 30243
rect 9689 30209 9723 30243
rect 6837 30141 6871 30175
rect 8401 30141 8435 30175
rect 8712 30141 8746 30175
rect 5089 30073 5123 30107
rect 5181 30073 5215 30107
rect 7113 30073 7147 30107
rect 10010 30073 10044 30107
rect 6377 30005 6411 30039
rect 9137 30005 9171 30039
rect 9505 30005 9539 30039
rect 4629 29801 4663 29835
rect 7573 29801 7607 29835
rect 7849 29801 7883 29835
rect 8401 29801 8435 29835
rect 9505 29801 9539 29835
rect 11253 29801 11287 29835
rect 4905 29733 4939 29767
rect 6974 29733 7008 29767
rect 9873 29733 9907 29767
rect 12265 29665 12299 29699
rect 2881 29597 2915 29631
rect 4813 29597 4847 29631
rect 6653 29597 6687 29631
rect 9781 29597 9815 29631
rect 10425 29597 10459 29631
rect 5365 29529 5399 29563
rect 3111 29461 3145 29495
rect 5733 29461 5767 29495
rect 6285 29461 6319 29495
rect 10701 29461 10735 29495
rect 12403 29461 12437 29495
rect 12909 29257 12943 29291
rect 4031 29189 4065 29223
rect 6561 29189 6595 29223
rect 8401 29189 8435 29223
rect 4997 29121 5031 29155
rect 5365 29121 5399 29155
rect 10885 29121 10919 29155
rect 3960 29053 3994 29087
rect 6837 29053 6871 29087
rect 7297 29053 7331 29087
rect 8585 29053 8619 29087
rect 9505 29053 9539 29087
rect 12449 29053 12483 29087
rect 13277 29053 13311 29087
rect 13528 29053 13562 29087
rect 13921 29053 13955 29087
rect 5089 28985 5123 29019
rect 8906 28985 8940 29019
rect 10425 28985 10459 29019
rect 10517 28985 10551 29019
rect 3065 28917 3099 28951
rect 4445 28917 4479 28951
rect 4721 28917 4755 28951
rect 6193 28917 6227 28951
rect 6929 28917 6963 28951
rect 8033 28917 8067 28951
rect 9873 28917 9907 28951
rect 10241 28917 10275 28951
rect 12633 28917 12667 28951
rect 13599 28917 13633 28951
rect 4629 28713 4663 28747
rect 6193 28713 6227 28747
rect 9965 28713 9999 28747
rect 4721 28645 4755 28679
rect 7021 28645 7055 28679
rect 8769 28645 8803 28679
rect 10333 28645 10367 28679
rect 11897 28645 11931 28679
rect 12449 28645 12483 28679
rect 4813 28577 4847 28611
rect 5733 28577 5767 28611
rect 6561 28577 6595 28611
rect 6745 28577 6779 28611
rect 7297 28577 7331 28611
rect 8125 28577 8159 28611
rect 8493 28577 8527 28611
rect 10885 28577 10919 28611
rect 13277 28577 13311 28611
rect 10241 28509 10275 28543
rect 11805 28509 11839 28543
rect 13415 28373 13449 28407
rect 4537 28169 4571 28203
rect 5917 28169 5951 28203
rect 6285 28169 6319 28203
rect 8309 28169 8343 28203
rect 9689 28169 9723 28203
rect 11161 28169 11195 28203
rect 11437 28169 11471 28203
rect 11805 28169 11839 28203
rect 13645 28169 13679 28203
rect 6561 28033 6595 28067
rect 8033 28033 8067 28067
rect 3709 27965 3743 27999
rect 3801 27965 3835 27999
rect 4169 27965 4203 27999
rect 4997 27965 5031 27999
rect 6929 27965 6963 27999
rect 7481 27965 7515 27999
rect 7665 27965 7699 27999
rect 8493 27965 8527 27999
rect 9413 27965 9447 27999
rect 10241 27965 10275 27999
rect 12633 27965 12667 27999
rect 13369 27965 13403 27999
rect 3341 27897 3375 27931
rect 5318 27897 5352 27931
rect 8815 27897 8849 27931
rect 10603 27897 10637 27931
rect 12449 27897 12483 27931
rect 4905 27829 4939 27863
rect 10057 27829 10091 27863
rect 12173 27829 12207 27863
rect 12725 27829 12759 27863
rect 4721 27625 4755 27659
rect 5273 27625 5307 27659
rect 7021 27625 7055 27659
rect 8033 27625 8067 27659
rect 8953 27625 8987 27659
rect 12633 27625 12667 27659
rect 10149 27557 10183 27591
rect 10701 27557 10735 27591
rect 11345 27557 11379 27591
rect 11713 27557 11747 27591
rect 13231 27557 13265 27591
rect 3525 27489 3559 27523
rect 4169 27489 4203 27523
rect 5457 27489 5491 27523
rect 5641 27489 5675 27523
rect 6009 27489 6043 27523
rect 7941 27489 7975 27523
rect 8493 27489 8527 27523
rect 12265 27489 12299 27523
rect 13093 27489 13127 27523
rect 10057 27421 10091 27455
rect 11621 27421 11655 27455
rect 4353 27353 4387 27387
rect 10977 27353 11011 27387
rect 5089 27285 5123 27319
rect 6653 27285 6687 27319
rect 9505 27285 9539 27319
rect 4169 27081 4203 27115
rect 5917 27081 5951 27115
rect 6193 27081 6227 27115
rect 7021 27081 7055 27115
rect 10057 27081 10091 27115
rect 11621 27081 11655 27115
rect 12587 27081 12621 27115
rect 13093 27081 13127 27115
rect 7389 27013 7423 27047
rect 4905 26945 4939 26979
rect 8677 26945 8711 26979
rect 10517 26945 10551 26979
rect 12173 26945 12207 26979
rect 4997 26877 5031 26911
rect 6837 26877 6871 26911
rect 7941 26877 7975 26911
rect 8493 26877 8527 26911
rect 12484 26877 12518 26911
rect 5318 26809 5352 26843
rect 6561 26809 6595 26843
rect 10609 26809 10643 26843
rect 11161 26809 11195 26843
rect 7849 26741 7883 26775
rect 8953 26741 8987 26775
rect 9321 26741 9355 26775
rect 10057 26537 10091 26571
rect 10425 26537 10459 26571
rect 11529 26537 11563 26571
rect 12219 26537 12253 26571
rect 4813 26469 4847 26503
rect 10701 26469 10735 26503
rect 11253 26469 11287 26503
rect 4905 26401 4939 26435
rect 7021 26401 7055 26435
rect 8033 26401 8067 26435
rect 8585 26401 8619 26435
rect 12116 26401 12150 26435
rect 7113 26333 7147 26367
rect 7849 26333 7883 26367
rect 8769 26333 8803 26367
rect 10609 26333 10643 26367
rect 4721 26197 4755 26231
rect 5825 26197 5859 26231
rect 9321 26197 9355 26231
rect 4905 25993 4939 26027
rect 6469 25993 6503 26027
rect 9045 25993 9079 26027
rect 9137 25993 9171 26027
rect 10241 25993 10275 26027
rect 10885 25993 10919 26027
rect 11483 25993 11517 26027
rect 12081 25993 12115 26027
rect 5917 25857 5951 25891
rect 4537 25789 4571 25823
rect 5549 25789 5583 25823
rect 7757 25789 7791 25823
rect 8309 25789 8343 25823
rect 5365 25721 5399 25755
rect 7573 25721 7607 25755
rect 8493 25721 8527 25755
rect 9321 25789 9355 25823
rect 11380 25789 11414 25823
rect 9643 25721 9677 25755
rect 5181 25653 5215 25687
rect 8769 25653 8803 25687
rect 9045 25653 9079 25687
rect 10609 25653 10643 25687
rect 5365 25449 5399 25483
rect 6653 25449 6687 25483
rect 7113 25449 7147 25483
rect 9045 25449 9079 25483
rect 9413 25449 9447 25483
rect 10057 25449 10091 25483
rect 10609 25449 10643 25483
rect 11437 25449 11471 25483
rect 5181 25381 5215 25415
rect 11897 25381 11931 25415
rect 5549 25313 5583 25347
rect 6101 25313 6135 25347
rect 7205 25313 7239 25347
rect 7297 25313 7331 25347
rect 9689 25313 9723 25347
rect 10977 25313 11011 25347
rect 6193 25245 6227 25279
rect 4445 25109 4479 25143
rect 4813 25109 4847 25143
rect 8217 25109 8251 25143
rect 5457 24905 5491 24939
rect 7665 24905 7699 24939
rect 7159 24837 7193 24871
rect 7297 24837 7331 24871
rect 8861 24837 8895 24871
rect 5089 24769 5123 24803
rect 5549 24769 5583 24803
rect 6653 24769 6687 24803
rect 7389 24769 7423 24803
rect 9045 24769 9079 24803
rect 10885 24769 10919 24803
rect 11253 24769 11287 24803
rect 3985 24701 4019 24735
rect 5328 24701 5362 24735
rect 8033 24701 8067 24735
rect 9965 24701 9999 24735
rect 10609 24701 10643 24735
rect 3801 24633 3835 24667
rect 4353 24633 4387 24667
rect 5181 24633 5215 24667
rect 5917 24633 5951 24667
rect 6285 24633 6319 24667
rect 7021 24633 7055 24667
rect 9407 24633 9441 24667
rect 10241 24633 10275 24667
rect 10977 24633 11011 24667
rect 3617 24565 3651 24599
rect 4721 24565 4755 24599
rect 8493 24565 8527 24599
rect 7205 24361 7239 24395
rect 7849 24361 7883 24395
rect 9781 24361 9815 24395
rect 5273 24293 5307 24327
rect 6653 24293 6687 24327
rect 11253 24293 11287 24327
rect 2973 24225 3007 24259
rect 4261 24225 4295 24259
rect 5733 24225 5767 24259
rect 6193 24225 6227 24259
rect 6745 24225 6779 24259
rect 7021 24225 7055 24259
rect 8309 24225 8343 24259
rect 8769 24225 8803 24259
rect 9689 24225 9723 24259
rect 10149 24225 10183 24259
rect 11345 24225 11379 24259
rect 12541 24225 12575 24259
rect 4169 24157 4203 24191
rect 3525 24089 3559 24123
rect 5641 24089 5675 24123
rect 6837 24089 6871 24123
rect 8493 24089 8527 24123
rect 3157 24021 3191 24055
rect 5917 24021 5951 24055
rect 9137 24021 9171 24055
rect 10701 24021 10735 24055
rect 11161 24021 11195 24055
rect 2789 23817 2823 23851
rect 4353 23817 4387 23851
rect 4721 23817 4755 23851
rect 6653 23817 6687 23851
rect 7573 23817 7607 23851
rect 8217 23817 8251 23851
rect 8953 23817 8987 23851
rect 10149 23817 10183 23851
rect 11529 23817 11563 23851
rect 12725 23817 12759 23851
rect 3341 23749 3375 23783
rect 7251 23749 7285 23783
rect 7389 23749 7423 23783
rect 8585 23749 8619 23783
rect 8815 23749 8849 23783
rect 12265 23749 12299 23783
rect 12587 23749 12621 23783
rect 3985 23681 4019 23715
rect 6285 23681 6319 23715
rect 7481 23681 7515 23715
rect 9045 23681 9079 23715
rect 10517 23681 10551 23715
rect 11897 23681 11931 23715
rect 12817 23681 12851 23715
rect 3157 23613 3191 23647
rect 3249 23613 3283 23647
rect 3525 23613 3559 23647
rect 4813 23613 4847 23647
rect 5641 23613 5675 23647
rect 5825 23613 5859 23647
rect 9413 23613 9447 23647
rect 7113 23545 7147 23579
rect 8677 23545 8711 23579
rect 10609 23545 10643 23579
rect 11161 23545 11195 23579
rect 12449 23545 12483 23579
rect 4905 23477 4939 23511
rect 9689 23477 9723 23511
rect 13093 23477 13127 23511
rect 3893 23273 3927 23307
rect 5365 23273 5399 23307
rect 6745 23273 6779 23307
rect 7481 23273 7515 23307
rect 9045 23273 9079 23307
rect 12725 23273 12759 23307
rect 2605 23205 2639 23239
rect 3525 23205 3559 23239
rect 7205 23205 7239 23239
rect 10517 23205 10551 23239
rect 2789 23137 2823 23171
rect 4128 23137 4162 23171
rect 4905 23137 4939 23171
rect 5457 23137 5491 23171
rect 5733 23137 5767 23171
rect 6101 23137 6135 23171
rect 8033 23137 8067 23171
rect 8493 23137 8527 23171
rect 11897 23137 11931 23171
rect 12081 23137 12115 23171
rect 3157 23069 3191 23103
rect 8769 23069 8803 23103
rect 10241 23069 10275 23103
rect 10425 23069 10459 23103
rect 4215 23001 4249 23035
rect 10977 23001 11011 23035
rect 12173 22933 12207 22967
rect 2237 22729 2271 22763
rect 4353 22729 4387 22763
rect 4813 22729 4847 22763
rect 6469 22729 6503 22763
rect 8033 22729 8067 22763
rect 8953 22729 8987 22763
rect 11989 22729 12023 22763
rect 12909 22729 12943 22763
rect 6101 22661 6135 22695
rect 9965 22661 9999 22695
rect 12587 22661 12621 22695
rect 4905 22593 4939 22627
rect 7205 22593 7239 22627
rect 9045 22593 9079 22627
rect 11161 22593 11195 22627
rect 13599 22593 13633 22627
rect 2329 22525 2363 22559
rect 4077 22525 4111 22559
rect 12357 22525 12391 22559
rect 13496 22525 13530 22559
rect 13921 22525 13955 22559
rect 3433 22457 3467 22491
rect 3525 22457 3559 22491
rect 5226 22457 5260 22491
rect 6929 22457 6963 22491
rect 7021 22457 7055 22491
rect 10885 22457 10919 22491
rect 10977 22457 11011 22491
rect 2513 22389 2547 22423
rect 2881 22389 2915 22423
rect 3249 22389 3283 22423
rect 5825 22389 5859 22423
rect 8493 22389 8527 22423
rect 9413 22389 9447 22423
rect 10333 22389 10367 22423
rect 2697 22185 2731 22219
rect 3111 22185 3145 22219
rect 3433 22185 3467 22219
rect 4537 22185 4571 22219
rect 5365 22185 5399 22219
rect 6285 22185 6319 22219
rect 7021 22185 7055 22219
rect 9045 22185 9079 22219
rect 10977 22185 11011 22219
rect 4813 22117 4847 22151
rect 6653 22117 6687 22151
rect 8211 22117 8245 22151
rect 10010 22117 10044 22151
rect 11621 22117 11655 22151
rect 12449 22117 12483 22151
rect 13185 22117 13219 22151
rect 3040 22049 3074 22083
rect 4997 22049 5031 22083
rect 6837 22049 6871 22083
rect 8769 22049 8803 22083
rect 7389 21981 7423 22015
rect 7849 21981 7883 22015
rect 9689 21981 9723 22015
rect 11529 21981 11563 22015
rect 13093 21981 13127 22015
rect 13369 21981 13403 22015
rect 7665 21913 7699 21947
rect 12081 21913 12115 21947
rect 5917 21845 5951 21879
rect 10609 21845 10643 21879
rect 11345 21845 11379 21879
rect 4169 21641 4203 21675
rect 5641 21641 5675 21675
rect 7849 21641 7883 21675
rect 9137 21641 9171 21675
rect 9413 21641 9447 21675
rect 10517 21641 10551 21675
rect 11253 21641 11287 21675
rect 12173 21641 12207 21675
rect 13461 21641 13495 21675
rect 6561 21573 6595 21607
rect 11483 21573 11517 21607
rect 13829 21573 13863 21607
rect 3801 21505 3835 21539
rect 4721 21505 4755 21539
rect 4997 21505 5031 21539
rect 12817 21505 12851 21539
rect 6996 21437 7030 21471
rect 7389 21437 7423 21471
rect 7941 21437 7975 21471
rect 8401 21437 8435 21471
rect 9597 21437 9631 21471
rect 10793 21437 10827 21471
rect 11380 21437 11414 21471
rect 4813 21369 4847 21403
rect 8677 21369 8711 21403
rect 9918 21369 9952 21403
rect 12541 21369 12575 21403
rect 12633 21369 12667 21403
rect 3065 21301 3099 21335
rect 4537 21301 4571 21335
rect 7067 21301 7101 21335
rect 11805 21301 11839 21335
rect 7481 21097 7515 21131
rect 7941 21097 7975 21131
rect 8125 21097 8159 21131
rect 9045 21097 9079 21131
rect 10057 21097 10091 21131
rect 10609 21097 10643 21131
rect 12449 21097 12483 21131
rect 7205 21029 7239 21063
rect 11621 21029 11655 21063
rect 4905 20961 4939 20995
rect 6469 20961 6503 20995
rect 7021 20961 7055 20995
rect 8033 20961 8067 20995
rect 8493 20961 8527 20995
rect 13068 20961 13102 20995
rect 4445 20893 4479 20927
rect 9689 20893 9723 20927
rect 11529 20893 11563 20927
rect 12081 20825 12115 20859
rect 9505 20757 9539 20791
rect 10977 20757 11011 20791
rect 12817 20757 12851 20791
rect 13139 20757 13173 20791
rect 4261 20553 4295 20587
rect 5365 20553 5399 20587
rect 5733 20553 5767 20587
rect 6561 20553 6595 20587
rect 7205 20553 7239 20587
rect 8401 20553 8435 20587
rect 8861 20553 8895 20587
rect 10149 20553 10183 20587
rect 11713 20553 11747 20587
rect 12587 20553 12621 20587
rect 13277 20553 13311 20587
rect 13921 20553 13955 20587
rect 4997 20485 5031 20519
rect 11345 20485 11379 20519
rect 12081 20485 12115 20519
rect 8953 20417 8987 20451
rect 10793 20417 10827 20451
rect 13599 20417 13633 20451
rect 7389 20349 7423 20383
rect 7849 20349 7883 20383
rect 8125 20349 8159 20383
rect 9873 20349 9907 20383
rect 12357 20349 12391 20383
rect 13512 20349 13546 20383
rect 4445 20281 4479 20315
rect 4537 20281 4571 20315
rect 9315 20281 9349 20315
rect 10885 20281 10919 20315
rect 12909 20281 12943 20315
rect 3341 20213 3375 20247
rect 3801 20213 3835 20247
rect 6101 20213 6135 20247
rect 10609 20213 10643 20247
rect 8401 20009 8435 20043
rect 9505 20009 9539 20043
rect 11897 20009 11931 20043
rect 3111 19941 3145 19975
rect 10425 19941 10459 19975
rect 10517 19941 10551 19975
rect 11069 19941 11103 19975
rect 3024 19873 3058 19907
rect 4905 19873 4939 19907
rect 6469 19873 6503 19907
rect 7113 19873 7147 19907
rect 7389 19873 7423 19907
rect 7481 19873 7515 19907
rect 7665 19873 7699 19907
rect 9965 19873 9999 19907
rect 4997 19805 5031 19839
rect 7849 19805 7883 19839
rect 6837 19737 6871 19771
rect 7113 19737 7147 19771
rect 7205 19737 7239 19771
rect 5273 19669 5307 19703
rect 6101 19669 6135 19703
rect 8769 19669 8803 19703
rect 2973 19465 3007 19499
rect 4997 19465 5031 19499
rect 8217 19465 8251 19499
rect 10977 19465 11011 19499
rect 5273 19397 5307 19431
rect 6285 19397 6319 19431
rect 8493 19397 8527 19431
rect 4077 19329 4111 19363
rect 6929 19329 6963 19363
rect 3709 19261 3743 19295
rect 4169 19261 4203 19295
rect 5181 19261 5215 19295
rect 5457 19261 5491 19295
rect 6837 19261 6871 19295
rect 7113 19261 7147 19295
rect 7849 19261 7883 19295
rect 8401 19261 8435 19295
rect 8677 19261 8711 19295
rect 9965 19261 9999 19295
rect 10425 19261 10459 19295
rect 4721 19193 4755 19227
rect 6653 19193 6687 19227
rect 7573 19193 7607 19227
rect 4353 19125 4387 19159
rect 5641 19125 5675 19159
rect 8861 19125 8895 19159
rect 9781 19125 9815 19159
rect 10057 19125 10091 19159
rect 5181 18921 5215 18955
rect 5825 18921 5859 18955
rect 6101 18921 6135 18955
rect 7481 18921 7515 18955
rect 9873 18921 9907 18955
rect 10425 18921 10459 18955
rect 4629 18853 4663 18887
rect 7941 18853 7975 18887
rect 4721 18785 4755 18819
rect 4997 18785 5031 18819
rect 6285 18785 6319 18819
rect 6561 18785 6595 18819
rect 8033 18785 8067 18819
rect 8585 18785 8619 18819
rect 9689 18785 9723 18819
rect 10701 18785 10735 18819
rect 6377 18717 6411 18751
rect 7021 18717 7055 18751
rect 8769 18717 8803 18751
rect 11713 18717 11747 18751
rect 4813 18649 4847 18683
rect 10885 18581 10919 18615
rect 2881 18377 2915 18411
rect 9321 18377 9355 18411
rect 10701 18377 10735 18411
rect 3893 18309 3927 18343
rect 4813 18309 4847 18343
rect 6285 18309 6319 18343
rect 11345 18309 11379 18343
rect 8861 18241 8895 18275
rect 2973 18173 3007 18207
rect 3525 18173 3559 18207
rect 3985 18173 4019 18207
rect 5273 18173 5307 18207
rect 5457 18173 5491 18207
rect 6837 18173 6871 18207
rect 7573 18173 7607 18207
rect 7849 18173 7883 18207
rect 8401 18173 8435 18207
rect 8585 18173 8619 18207
rect 9413 18173 9447 18207
rect 11161 18173 11195 18207
rect 11621 18173 11655 18207
rect 7389 18105 7423 18139
rect 3157 18037 3191 18071
rect 4169 18037 4203 18071
rect 5089 18037 5123 18071
rect 7021 18037 7055 18071
rect 7573 18037 7607 18071
rect 7665 18037 7699 18071
rect 9781 18037 9815 18071
rect 10333 18037 10367 18071
rect 5273 17833 5307 17867
rect 6653 17833 6687 17867
rect 7021 17833 7055 17867
rect 9413 17833 9447 17867
rect 6377 17765 6411 17799
rect 8493 17765 8527 17799
rect 10010 17765 10044 17799
rect 11529 17765 11563 17799
rect 11621 17765 11655 17799
rect 2973 17697 3007 17731
rect 4905 17697 4939 17731
rect 7573 17697 7607 17731
rect 7941 17697 7975 17731
rect 9689 17697 9723 17731
rect 8033 17629 8067 17663
rect 12173 17629 12207 17663
rect 3157 17493 3191 17527
rect 4813 17493 4847 17527
rect 5825 17493 5859 17527
rect 10609 17493 10643 17527
rect 12541 17493 12575 17527
rect 3065 17289 3099 17323
rect 4629 17289 4663 17323
rect 7389 17289 7423 17323
rect 9045 17289 9079 17323
rect 10333 17289 10367 17323
rect 11713 17289 11747 17323
rect 12173 17289 12207 17323
rect 4261 17221 4295 17255
rect 6561 17153 6595 17187
rect 12817 17153 12851 17187
rect 3709 17085 3743 17119
rect 4721 17085 4755 17119
rect 5549 17085 5583 17119
rect 5733 17085 5767 17119
rect 6193 17085 6227 17119
rect 7573 17085 7607 17119
rect 8033 17085 8067 17119
rect 8309 17085 8343 17119
rect 9137 17085 9171 17119
rect 10057 17085 10091 17119
rect 10920 17085 10954 17119
rect 11345 17085 11379 17119
rect 9499 17017 9533 17051
rect 12541 17017 12575 17051
rect 12633 17017 12667 17051
rect 3893 16949 3927 16983
rect 4905 16949 4939 16983
rect 5273 16949 5307 16983
rect 5917 16949 5951 16983
rect 7113 16949 7147 16983
rect 11023 16949 11057 16983
rect 5825 16745 5859 16779
rect 9137 16745 9171 16779
rect 9873 16745 9907 16779
rect 11529 16745 11563 16779
rect 8211 16677 8245 16711
rect 10701 16677 10735 16711
rect 12265 16677 12299 16711
rect 12817 16677 12851 16711
rect 2973 16609 3007 16643
rect 4997 16609 5031 16643
rect 5273 16609 5307 16643
rect 6561 16609 6595 16643
rect 6837 16609 6871 16643
rect 7849 16609 7883 16643
rect 5457 16541 5491 16575
rect 7021 16541 7055 16575
rect 10609 16541 10643 16575
rect 11069 16541 11103 16575
rect 12173 16541 12207 16575
rect 3157 16405 3191 16439
rect 4629 16405 4663 16439
rect 7573 16405 7607 16439
rect 8769 16405 8803 16439
rect 4813 16201 4847 16235
rect 6377 16201 6411 16235
rect 7389 16201 7423 16235
rect 8585 16201 8619 16235
rect 8953 16201 8987 16235
rect 11023 16201 11057 16235
rect 11713 16201 11747 16235
rect 12173 16201 12207 16235
rect 12587 16201 12621 16235
rect 4261 16133 4295 16167
rect 7021 16133 7055 16167
rect 12909 16133 12943 16167
rect 9137 16065 9171 16099
rect 11345 16065 11379 16099
rect 4077 15997 4111 16031
rect 5089 15997 5123 16031
rect 5549 15997 5583 16031
rect 7849 15997 7883 16031
rect 8033 15997 8067 16031
rect 10920 15997 10954 16031
rect 12516 15997 12550 16031
rect 13277 15997 13311 16031
rect 5825 15929 5859 15963
rect 8309 15929 8343 15963
rect 9458 15929 9492 15963
rect 3065 15861 3099 15895
rect 3985 15861 4019 15895
rect 10057 15861 10091 15895
rect 10609 15861 10643 15895
rect 4813 15657 4847 15691
rect 6837 15657 6871 15691
rect 7021 15657 7055 15691
rect 7941 15657 7975 15691
rect 8309 15657 8343 15691
rect 9137 15657 9171 15691
rect 10057 15657 10091 15691
rect 5543 15589 5577 15623
rect 11529 15589 11563 15623
rect 11621 15589 11655 15623
rect 6929 15521 6963 15555
rect 7481 15521 7515 15555
rect 8493 15521 8527 15555
rect 9689 15521 9723 15555
rect 13001 15521 13035 15555
rect 5181 15453 5215 15487
rect 8677 15385 8711 15419
rect 12081 15385 12115 15419
rect 6101 15317 6135 15351
rect 10609 15317 10643 15351
rect 10977 15317 11011 15351
rect 13139 15317 13173 15351
rect 8033 15113 8067 15147
rect 8401 15113 8435 15147
rect 8861 15113 8895 15147
rect 10149 15113 10183 15147
rect 10609 15113 10643 15147
rect 11713 15113 11747 15147
rect 13001 15045 13035 15079
rect 4537 14977 4571 15011
rect 6837 14977 6871 15011
rect 8953 14977 8987 15011
rect 10793 14977 10827 15011
rect 13599 14977 13633 15011
rect 4905 14909 4939 14943
rect 5273 14909 5307 14943
rect 5549 14909 5583 14943
rect 12265 14909 12299 14943
rect 12516 14909 12550 14943
rect 13496 14909 13530 14943
rect 6101 14841 6135 14875
rect 6653 14841 6687 14875
rect 7199 14841 7233 14875
rect 9274 14841 9308 14875
rect 10885 14841 10919 14875
rect 11437 14841 11471 14875
rect 5273 14773 5307 14807
rect 7757 14773 7791 14807
rect 9873 14773 9907 14807
rect 12587 14773 12621 14807
rect 13921 14773 13955 14807
rect 5457 14569 5491 14603
rect 5825 14569 5859 14603
rect 7389 14569 7423 14603
rect 7849 14569 7883 14603
rect 8033 14569 8067 14603
rect 8953 14569 8987 14603
rect 9965 14569 9999 14603
rect 11437 14569 11471 14603
rect 6561 14501 6595 14535
rect 10517 14501 10551 14535
rect 12081 14501 12115 14535
rect 4905 14433 4939 14467
rect 7941 14433 7975 14467
rect 8401 14433 8435 14467
rect 11069 14433 11103 14467
rect 6469 14365 6503 14399
rect 6745 14365 6779 14399
rect 10425 14365 10459 14399
rect 11989 14365 12023 14399
rect 12541 14297 12575 14331
rect 5135 14229 5169 14263
rect 3019 14025 3053 14059
rect 6285 14025 6319 14059
rect 6653 14025 6687 14059
rect 7941 14025 7975 14059
rect 10057 14025 10091 14059
rect 11161 14025 11195 14059
rect 11621 14025 11655 14059
rect 12725 14025 12759 14059
rect 4031 13957 4065 13991
rect 11897 13957 11931 13991
rect 4445 13889 4479 13923
rect 4905 13889 4939 13923
rect 6929 13889 6963 13923
rect 7389 13889 7423 13923
rect 10885 13889 10919 13923
rect 2948 13821 2982 13855
rect 3960 13821 3994 13855
rect 8401 13821 8435 13855
rect 8861 13821 8895 13855
rect 9413 13821 9447 13855
rect 4813 13753 4847 13787
rect 7021 13753 7055 13787
rect 10241 13753 10275 13787
rect 10333 13753 10367 13787
rect 3433 13685 3467 13719
rect 5273 13685 5307 13719
rect 5825 13685 5859 13719
rect 8677 13685 8711 13719
rect 6745 13481 6779 13515
rect 7113 13481 7147 13515
rect 10701 13481 10735 13515
rect 11391 13481 11425 13515
rect 4353 13413 4387 13447
rect 5917 13413 5951 13447
rect 7941 13413 7975 13447
rect 9873 13413 9907 13447
rect 11320 13345 11354 13379
rect 4261 13277 4295 13311
rect 4905 13277 4939 13311
rect 5825 13277 5859 13311
rect 7665 13277 7699 13311
rect 9781 13277 9815 13311
rect 6377 13209 6411 13243
rect 8861 13209 8895 13243
rect 10333 13209 10367 13243
rect 5273 13141 5307 13175
rect 8585 13141 8619 13175
rect 3709 12937 3743 12971
rect 6193 12937 6227 12971
rect 7665 12937 7699 12971
rect 8953 12937 8987 12971
rect 10885 12937 10919 12971
rect 4077 12869 4111 12903
rect 6561 12869 6595 12903
rect 10517 12869 10551 12903
rect 7297 12801 7331 12835
rect 7757 12801 7791 12835
rect 9413 12801 9447 12835
rect 4220 12733 4254 12767
rect 11136 12733 11170 12767
rect 11529 12733 11563 12767
rect 4307 12665 4341 12699
rect 5273 12665 5307 12699
rect 5365 12665 5399 12699
rect 5917 12665 5951 12699
rect 8078 12665 8112 12699
rect 9597 12665 9631 12699
rect 9689 12665 9723 12699
rect 10241 12665 10275 12699
rect 4721 12597 4755 12631
rect 5089 12597 5123 12631
rect 8677 12597 8711 12631
rect 11207 12597 11241 12631
rect 11989 12597 12023 12631
rect 5043 12393 5077 12427
rect 5365 12393 5399 12427
rect 7849 12393 7883 12427
rect 6101 12325 6135 12359
rect 8217 12325 8251 12359
rect 9873 12325 9907 12359
rect 11345 12325 11379 12359
rect 11437 12325 11471 12359
rect 12868 12257 12902 12291
rect 6009 12189 6043 12223
rect 6285 12189 6319 12223
rect 8125 12189 8159 12223
rect 9781 12189 9815 12223
rect 12955 12189 12989 12223
rect 8677 12121 8711 12155
rect 10333 12121 10367 12155
rect 11897 12121 11931 12155
rect 4813 12053 4847 12087
rect 9505 12053 9539 12087
rect 4905 11849 4939 11883
rect 5641 11849 5675 11883
rect 6561 11849 6595 11883
rect 7297 11849 7331 11883
rect 7665 11849 7699 11883
rect 8677 11849 8711 11883
rect 11161 11849 11195 11883
rect 12081 11849 12115 11883
rect 13001 11849 13035 11883
rect 9597 11781 9631 11815
rect 13277 11781 13311 11815
rect 6285 11713 6319 11747
rect 9781 11713 9815 11747
rect 11391 11713 11425 11747
rect 4721 11645 4755 11679
rect 5800 11645 5834 11679
rect 7757 11645 7791 11679
rect 8953 11645 8987 11679
rect 11288 11645 11322 11679
rect 11713 11645 11747 11679
rect 12516 11645 12550 11679
rect 5273 11577 5307 11611
rect 8078 11577 8112 11611
rect 9873 11577 9907 11611
rect 10425 11577 10459 11611
rect 5871 11509 5905 11543
rect 10701 11509 10735 11543
rect 12587 11509 12621 11543
rect 5733 11305 5767 11339
rect 6101 11305 6135 11339
rect 7297 11305 7331 11339
rect 9137 11305 9171 11339
rect 9505 11305 9539 11339
rect 11391 11305 11425 11339
rect 7021 11237 7055 11271
rect 8170 11237 8204 11271
rect 9873 11237 9907 11271
rect 10425 11237 10459 11271
rect 4721 11169 4755 11203
rect 5273 11169 5307 11203
rect 6561 11169 6595 11203
rect 6837 11169 6871 11203
rect 11288 11169 11322 11203
rect 12332 11169 12366 11203
rect 5457 11101 5491 11135
rect 7849 11101 7883 11135
rect 9781 11101 9815 11135
rect 7757 11033 7791 11067
rect 12403 11033 12437 11067
rect 8769 10965 8803 10999
rect 4077 10761 4111 10795
rect 4813 10761 4847 10795
rect 7941 10761 7975 10795
rect 9505 10761 9539 10795
rect 11437 10761 11471 10795
rect 5549 10625 5583 10659
rect 7205 10625 7239 10659
rect 8585 10625 8619 10659
rect 8861 10625 8895 10659
rect 10425 10625 10459 10659
rect 11805 10625 11839 10659
rect 4169 10489 4203 10523
rect 5273 10489 5307 10523
rect 5365 10489 5399 10523
rect 6929 10489 6963 10523
rect 7021 10489 7055 10523
rect 8677 10489 8711 10523
rect 9965 10489 9999 10523
rect 10149 10489 10183 10523
rect 10241 10489 10275 10523
rect 6377 10421 6411 10455
rect 8401 10421 8435 10455
rect 11069 10421 11103 10455
rect 12633 10421 12667 10455
rect 5273 10217 5307 10251
rect 6837 10217 6871 10251
rect 8309 10217 8343 10251
rect 8677 10217 8711 10251
rect 10609 10217 10643 10251
rect 5911 10149 5945 10183
rect 7481 10149 7515 10183
rect 10010 10149 10044 10183
rect 11437 10149 11471 10183
rect 4537 10081 4571 10115
rect 6469 10081 6503 10115
rect 7113 10081 7147 10115
rect 5549 10013 5583 10047
rect 7389 10013 7423 10047
rect 7665 10013 7699 10047
rect 9689 10013 9723 10047
rect 9045 9945 9079 9979
rect 4721 9877 4755 9911
rect 4537 9673 4571 9707
rect 9781 9673 9815 9707
rect 5917 9605 5951 9639
rect 7849 9605 7883 9639
rect 10701 9537 10735 9571
rect 11345 9537 11379 9571
rect 4169 9469 4203 9503
rect 4997 9469 5031 9503
rect 7113 9469 7147 9503
rect 7297 9469 7331 9503
rect 8401 9469 8435 9503
rect 8861 9469 8895 9503
rect 10241 9469 10275 9503
rect 10425 9469 10459 9503
rect 4905 9401 4939 9435
rect 5359 9401 5393 9435
rect 6561 9401 6595 9435
rect 8309 9401 8343 9435
rect 9137 9401 9171 9435
rect 10977 9401 11011 9435
rect 6285 9333 6319 9367
rect 6929 9333 6963 9367
rect 5181 9129 5215 9163
rect 5457 9129 5491 9163
rect 6469 9129 6503 9163
rect 9827 9129 9861 9163
rect 7475 9061 7509 9095
rect 8401 9061 8435 9095
rect 4353 8993 4387 9027
rect 5549 8993 5583 9027
rect 5825 8993 5859 9027
rect 6929 8993 6963 9027
rect 9724 8993 9758 9027
rect 10701 8993 10735 9027
rect 7113 8925 7147 8959
rect 8769 8925 8803 8959
rect 10517 8925 10551 8959
rect 10241 8857 10275 8891
rect 10885 8857 10919 8891
rect 4491 8789 4525 8823
rect 8033 8789 8067 8823
rect 4353 8585 4387 8619
rect 4997 8585 5031 8619
rect 6193 8585 6227 8619
rect 9229 8585 9263 8619
rect 9505 8585 9539 8619
rect 9689 8585 9723 8619
rect 10793 8585 10827 8619
rect 4721 8517 4755 8551
rect 7757 8517 7791 8551
rect 5917 8449 5951 8483
rect 7021 8449 7055 8483
rect 8125 8449 8159 8483
rect 5181 8381 5215 8415
rect 5641 8381 5675 8415
rect 8217 8381 8251 8415
rect 8769 8381 8803 8415
rect 9505 8381 9539 8415
rect 9781 8381 9815 8415
rect 10241 8381 10275 8415
rect 8953 8313 8987 8347
rect 7205 8245 7239 8279
rect 9873 8245 9907 8279
rect 6561 7973 6595 8007
rect 8125 7973 8159 8007
rect 10010 7973 10044 8007
rect 5089 7905 5123 7939
rect 5273 7905 5307 7939
rect 9689 7905 9723 7939
rect 5549 7837 5583 7871
rect 6469 7837 6503 7871
rect 7113 7837 7147 7871
rect 8033 7837 8067 7871
rect 8677 7837 8711 7871
rect 11437 7837 11471 7871
rect 6193 7701 6227 7735
rect 10609 7701 10643 7735
rect 4537 7497 4571 7531
rect 4905 7497 4939 7531
rect 7757 7497 7791 7531
rect 8125 7497 8159 7531
rect 10793 7497 10827 7531
rect 9137 7429 9171 7463
rect 11115 7429 11149 7463
rect 6837 7361 6871 7395
rect 9229 7361 9263 7395
rect 5181 7293 5215 7327
rect 5641 7293 5675 7327
rect 11012 7293 11046 7327
rect 11437 7293 11471 7327
rect 5917 7225 5951 7259
rect 6285 7225 6319 7259
rect 7199 7225 7233 7259
rect 9591 7225 9625 7259
rect 10425 7225 10459 7259
rect 6653 7157 6687 7191
rect 8401 7157 8435 7191
rect 10149 7157 10183 7191
rect 4951 6953 4985 6987
rect 7573 6953 7607 6987
rect 8125 6953 8159 6987
rect 9229 6953 9263 6987
rect 10609 6953 10643 6987
rect 5273 6885 5307 6919
rect 6187 6885 6221 6919
rect 7021 6885 7055 6919
rect 10010 6885 10044 6919
rect 10885 6885 10919 6919
rect 11621 6885 11655 6919
rect 4848 6817 4882 6851
rect 5641 6817 5675 6851
rect 7757 6817 7791 6851
rect 9689 6817 9723 6851
rect 5825 6749 5859 6783
rect 11529 6749 11563 6783
rect 11989 6749 12023 6783
rect 6745 6613 6779 6647
rect 8677 6613 8711 6647
rect 4813 6409 4847 6443
rect 8401 6409 8435 6443
rect 9781 6409 9815 6443
rect 11437 6409 11471 6443
rect 6653 6341 6687 6375
rect 7941 6341 7975 6375
rect 8677 6273 8711 6307
rect 8953 6273 8987 6307
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 5784 6205 5818 6239
rect 5871 6137 5905 6171
rect 6929 6137 6963 6171
rect 7021 6137 7055 6171
rect 7573 6137 7607 6171
rect 8769 6137 8803 6171
rect 10425 6137 10459 6171
rect 10977 6137 11011 6171
rect 5641 6069 5675 6103
rect 6193 6069 6227 6103
rect 11805 6069 11839 6103
rect 6101 5865 6135 5899
rect 7389 5865 7423 5899
rect 8769 5865 8803 5899
rect 9873 5865 9907 5899
rect 7021 5797 7055 5831
rect 7757 5797 7791 5831
rect 7849 5797 7883 5831
rect 8401 5797 8435 5831
rect 10241 5797 10275 5831
rect 6009 5729 6043 5763
rect 6469 5729 6503 5763
rect 10793 5729 10827 5763
rect 11688 5729 11722 5763
rect 10149 5661 10183 5695
rect 11759 5525 11793 5559
rect 5641 5321 5675 5355
rect 6377 5321 6411 5355
rect 6561 5321 6595 5355
rect 7205 5321 7239 5355
rect 9137 5321 9171 5355
rect 10609 5321 10643 5355
rect 11713 5321 11747 5355
rect 12909 5321 12943 5355
rect 6285 5253 6319 5287
rect 5871 5185 5905 5219
rect 8493 5253 8527 5287
rect 5784 5117 5818 5151
rect 6377 5117 6411 5151
rect 7665 5117 7699 5151
rect 8217 5117 8251 5151
rect 10333 5185 10367 5219
rect 9413 5117 9447 5151
rect 9689 5117 9723 5151
rect 10860 5117 10894 5151
rect 12500 5117 12534 5151
rect 7573 5049 7607 5083
rect 8401 5049 8435 5083
rect 8493 5049 8527 5083
rect 12587 5049 12621 5083
rect 8677 4981 8711 5015
rect 9321 4981 9355 5015
rect 10931 4981 10965 5015
rect 11345 4981 11379 5015
rect 5273 4777 5307 4811
rect 7665 4777 7699 4811
rect 9321 4777 9355 4811
rect 6653 4709 6687 4743
rect 9873 4709 9907 4743
rect 5508 4641 5542 4675
rect 8033 4641 8067 4675
rect 8585 4641 8619 4675
rect 11253 4641 11287 4675
rect 12357 4641 12391 4675
rect 13461 4641 13495 4675
rect 5595 4573 5629 4607
rect 6009 4573 6043 4607
rect 6561 4573 6595 4607
rect 8769 4573 8803 4607
rect 9781 4573 9815 4607
rect 10149 4573 10183 4607
rect 7113 4505 7147 4539
rect 10701 4505 10735 4539
rect 12541 4505 12575 4539
rect 6285 4437 6319 4471
rect 11437 4437 11471 4471
rect 13645 4437 13679 4471
rect 5089 4233 5123 4267
rect 7941 4233 7975 4267
rect 11345 4233 11379 4267
rect 12265 4233 12299 4267
rect 13461 4233 13495 4267
rect 4629 4165 4663 4199
rect 9597 4165 9631 4199
rect 9965 4165 9999 4199
rect 10793 4165 10827 4199
rect 6285 4097 6319 4131
rect 7205 4097 7239 4131
rect 8217 4097 8251 4131
rect 10241 4097 10275 4131
rect 11621 4097 11655 4131
rect 4236 4029 4270 4063
rect 5181 4029 5215 4063
rect 5641 4029 5675 4063
rect 8401 4029 8435 4063
rect 12449 4029 12483 4063
rect 13001 4029 13035 4063
rect 13620 4029 13654 4063
rect 14013 4029 14047 4063
rect 5917 3961 5951 3995
rect 6929 3961 6963 3995
rect 7021 3961 7055 3995
rect 8722 3961 8756 3995
rect 10333 3961 10367 3995
rect 4307 3893 4341 3927
rect 6653 3893 6687 3927
rect 9321 3893 9355 3927
rect 12633 3893 12667 3927
rect 13691 3893 13725 3927
rect 9045 3689 9079 3723
rect 9413 3689 9447 3723
rect 11161 3689 11195 3723
rect 6279 3621 6313 3655
rect 8170 3621 8204 3655
rect 9873 3621 9907 3655
rect 11437 3621 11471 3655
rect 4629 3553 4663 3587
rect 4905 3553 4939 3587
rect 5089 3553 5123 3587
rect 7113 3553 7147 3587
rect 7849 3553 7883 3587
rect 10701 3553 10735 3587
rect 13461 3553 13495 3587
rect 5917 3485 5951 3519
rect 9781 3485 9815 3519
rect 10425 3485 10459 3519
rect 11345 3485 11379 3519
rect 5457 3417 5491 3451
rect 6837 3417 6871 3451
rect 11897 3417 11931 3451
rect 5733 3349 5767 3383
rect 7481 3349 7515 3383
rect 8769 3349 8803 3383
rect 13645 3349 13679 3383
rect 4077 3145 4111 3179
rect 4997 3145 5031 3179
rect 6285 3145 6319 3179
rect 6653 3145 6687 3179
rect 8125 3145 8159 3179
rect 8401 3145 8435 3179
rect 9505 3145 9539 3179
rect 9873 3145 9907 3179
rect 10149 3145 10183 3179
rect 11437 3145 11471 3179
rect 11805 3145 11839 3179
rect 13001 3145 13035 3179
rect 13369 3145 13403 3179
rect 4307 3077 4341 3111
rect 7757 3077 7791 3111
rect 11161 3077 11195 3111
rect 12633 3077 12667 3111
rect 5273 3009 5307 3043
rect 5917 3009 5951 3043
rect 6837 3009 6871 3043
rect 8585 3009 8619 3043
rect 10701 3009 10735 3043
rect 3224 2941 3258 2975
rect 4236 2941 4270 2975
rect 13691 3009 13725 3043
rect 12449 2941 12483 2975
rect 13604 2941 13638 2975
rect 14013 2941 14047 2975
rect 3709 2873 3743 2907
rect 5365 2873 5399 2907
rect 7199 2873 7233 2907
rect 8906 2873 8940 2907
rect 10425 2873 10459 2907
rect 10517 2873 10551 2907
rect 11161 2873 11195 2907
rect 3295 2805 3329 2839
rect 4721 2805 4755 2839
rect 4537 2601 4571 2635
rect 6285 2601 6319 2635
rect 6745 2601 6779 2635
rect 8033 2601 8067 2635
rect 9597 2601 9631 2635
rect 12817 2601 12851 2635
rect 7113 2533 7147 2567
rect 7205 2533 7239 2567
rect 7757 2533 7791 2567
rect 9965 2533 9999 2567
rect 10517 2533 10551 2567
rect 4328 2465 4362 2499
rect 4721 2465 4755 2499
rect 5917 2465 5951 2499
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 11161 2465 11195 2499
rect 11345 2465 11379 2499
rect 11897 2465 11931 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 5273 2397 5307 2431
rect 8401 2397 8435 2431
rect 9873 2397 9907 2431
rect 10793 2397 10827 2431
rect 5181 2329 5215 2363
rect 11529 2329 11563 2363
rect 8769 2261 8803 2295
<< metal1 >>
rect 290 39584 296 39636
rect 348 39584 354 39636
rect 1394 39584 1400 39636
rect 1452 39624 1458 39636
rect 2130 39624 2136 39636
rect 1452 39596 2136 39624
rect 1452 39584 1458 39596
rect 2130 39584 2136 39596
rect 2188 39584 2194 39636
rect 6914 39584 6920 39636
rect 6972 39624 6978 39636
rect 8846 39624 8852 39636
rect 6972 39596 8852 39624
rect 6972 39584 6978 39596
rect 8846 39584 8852 39596
rect 8904 39584 8910 39636
rect 308 39556 336 39584
rect 3418 39556 3424 39568
rect 308 39528 3424 39556
rect 3418 39516 3424 39528
rect 3476 39516 3482 39568
rect 8386 39244 8392 39296
rect 8444 39284 8450 39296
rect 9214 39284 9220 39296
rect 8444 39256 9220 39284
rect 8444 39244 8450 39256
rect 9214 39244 9220 39256
rect 9272 39244 9278 39296
rect 1486 38972 1492 39024
rect 1544 39012 1550 39024
rect 2406 39012 2412 39024
rect 1544 38984 2412 39012
rect 1544 38972 1550 38984
rect 2406 38972 2412 38984
rect 2464 38972 2470 39024
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 8113 37111 8171 37117
rect 8113 37077 8125 37111
rect 8159 37108 8171 37111
rect 8570 37108 8576 37120
rect 8159 37080 8576 37108
rect 8159 37077 8171 37080
rect 8113 37071 8171 37077
rect 8570 37068 8576 37080
rect 8628 37068 8634 37120
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 10965 36907 11023 36913
rect 10965 36873 10977 36907
rect 11011 36904 11023 36907
rect 11514 36904 11520 36916
rect 11011 36876 11520 36904
rect 11011 36873 11023 36876
rect 10965 36867 11023 36873
rect 11514 36864 11520 36876
rect 11572 36864 11578 36916
rect 5350 36728 5356 36780
rect 5408 36768 5414 36780
rect 5408 36740 7972 36768
rect 5408 36728 5414 36740
rect 3050 36660 3056 36712
rect 3108 36700 3114 36712
rect 6952 36703 7010 36709
rect 6952 36700 6964 36703
rect 3108 36672 6964 36700
rect 3108 36660 3114 36672
rect 6952 36669 6964 36672
rect 6998 36700 7010 36703
rect 6998 36672 7144 36700
rect 6998 36669 7010 36672
rect 6952 36663 7010 36669
rect 7116 36632 7144 36672
rect 7190 36660 7196 36712
rect 7248 36700 7254 36712
rect 7650 36700 7656 36712
rect 7248 36672 7656 36700
rect 7248 36660 7254 36672
rect 7650 36660 7656 36672
rect 7708 36660 7714 36712
rect 7944 36709 7972 36740
rect 7929 36703 7987 36709
rect 7929 36669 7941 36703
rect 7975 36700 7987 36703
rect 8021 36703 8079 36709
rect 8021 36700 8033 36703
rect 7975 36672 8033 36700
rect 7975 36669 7987 36672
rect 7929 36663 7987 36669
rect 8021 36669 8033 36672
rect 8067 36669 8079 36703
rect 8570 36700 8576 36712
rect 8531 36672 8576 36700
rect 8021 36663 8079 36669
rect 8570 36660 8576 36672
rect 8628 36660 8634 36712
rect 10781 36703 10839 36709
rect 10781 36669 10793 36703
rect 10827 36700 10839 36703
rect 10827 36672 11192 36700
rect 10827 36669 10839 36672
rect 10781 36663 10839 36669
rect 7377 36635 7435 36641
rect 7377 36632 7389 36635
rect 7116 36604 7389 36632
rect 7377 36601 7389 36604
rect 7423 36632 7435 36635
rect 10226 36632 10232 36644
rect 7423 36604 10232 36632
rect 7423 36601 7435 36604
rect 7377 36595 7435 36601
rect 10226 36592 10232 36604
rect 10284 36592 10290 36644
rect 11164 36576 11192 36672
rect 7055 36567 7113 36573
rect 7055 36533 7067 36567
rect 7101 36564 7113 36567
rect 7190 36564 7196 36576
rect 7101 36536 7196 36564
rect 7101 36533 7113 36536
rect 7055 36527 7113 36533
rect 7190 36524 7196 36536
rect 7248 36524 7254 36576
rect 8294 36564 8300 36576
rect 8255 36536 8300 36564
rect 8294 36524 8300 36536
rect 8352 36524 8358 36576
rect 11146 36524 11152 36576
rect 11204 36564 11210 36576
rect 11333 36567 11391 36573
rect 11333 36564 11345 36567
rect 11204 36536 11345 36564
rect 11204 36524 11210 36536
rect 11333 36533 11345 36536
rect 11379 36533 11391 36567
rect 11333 36527 11391 36533
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 9861 36363 9919 36369
rect 9861 36329 9873 36363
rect 9907 36360 9919 36363
rect 10410 36360 10416 36372
rect 9907 36332 10416 36360
rect 9907 36329 9919 36332
rect 9861 36323 9919 36329
rect 10410 36320 10416 36332
rect 10468 36320 10474 36372
rect 11425 36363 11483 36369
rect 11425 36329 11437 36363
rect 11471 36360 11483 36363
rect 12618 36360 12624 36372
rect 11471 36332 12624 36360
rect 11471 36329 11483 36332
rect 11425 36323 11483 36329
rect 12618 36320 12624 36332
rect 12676 36320 12682 36372
rect 6638 36252 6644 36304
rect 6696 36292 6702 36304
rect 7285 36295 7343 36301
rect 7285 36292 7297 36295
rect 6696 36264 7297 36292
rect 6696 36252 6702 36264
rect 7285 36261 7297 36264
rect 7331 36261 7343 36295
rect 7285 36255 7343 36261
rect 9674 36224 9680 36236
rect 9635 36196 9680 36224
rect 9674 36184 9680 36196
rect 9732 36184 9738 36236
rect 11238 36224 11244 36236
rect 11199 36196 11244 36224
rect 11238 36184 11244 36196
rect 11296 36184 11302 36236
rect 7190 36156 7196 36168
rect 7151 36128 7196 36156
rect 7190 36116 7196 36128
rect 7248 36116 7254 36168
rect 7742 36088 7748 36100
rect 7703 36060 7748 36088
rect 7742 36048 7748 36060
rect 7800 36048 7806 36100
rect 8570 35980 8576 36032
rect 8628 36020 8634 36032
rect 8757 36023 8815 36029
rect 8757 36020 8769 36023
rect 8628 35992 8769 36020
rect 8628 35980 8634 35992
rect 8757 35989 8769 35992
rect 8803 36020 8815 36023
rect 9490 36020 9496 36032
rect 8803 35992 9496 36020
rect 8803 35989 8815 35992
rect 8757 35983 8815 35989
rect 9490 35980 9496 35992
rect 9548 35980 9554 36032
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 7190 35776 7196 35828
rect 7248 35816 7254 35828
rect 8113 35819 8171 35825
rect 8113 35816 8125 35819
rect 7248 35788 8125 35816
rect 7248 35776 7254 35788
rect 8113 35785 8125 35788
rect 8159 35785 8171 35819
rect 8113 35779 8171 35785
rect 10413 35819 10471 35825
rect 10413 35785 10425 35819
rect 10459 35816 10471 35819
rect 11054 35816 11060 35828
rect 10459 35788 11060 35816
rect 10459 35785 10471 35788
rect 10413 35779 10471 35785
rect 11054 35776 11060 35788
rect 11112 35776 11118 35828
rect 11471 35819 11529 35825
rect 11471 35785 11483 35819
rect 11517 35816 11529 35819
rect 12066 35816 12072 35828
rect 11517 35788 12072 35816
rect 11517 35785 11529 35788
rect 11471 35779 11529 35785
rect 12066 35776 12072 35788
rect 12124 35776 12130 35828
rect 12621 35819 12679 35825
rect 12621 35785 12633 35819
rect 12667 35816 12679 35819
rect 13722 35816 13728 35828
rect 12667 35788 13728 35816
rect 12667 35785 12679 35788
rect 12621 35779 12679 35785
rect 13722 35776 13728 35788
rect 13780 35776 13786 35828
rect 7742 35748 7748 35760
rect 7703 35720 7748 35748
rect 7742 35708 7748 35720
rect 7800 35708 7806 35760
rect 7834 35572 7840 35624
rect 7892 35612 7898 35624
rect 8573 35615 8631 35621
rect 8573 35612 8585 35615
rect 7892 35584 8585 35612
rect 7892 35572 7898 35584
rect 8573 35581 8585 35584
rect 8619 35612 8631 35615
rect 8665 35615 8723 35621
rect 8665 35612 8677 35615
rect 8619 35584 8677 35612
rect 8619 35581 8631 35584
rect 8573 35575 8631 35581
rect 8665 35581 8677 35584
rect 8711 35581 8723 35615
rect 8665 35575 8723 35581
rect 9217 35615 9275 35621
rect 9217 35581 9229 35615
rect 9263 35612 9275 35615
rect 9490 35612 9496 35624
rect 9263 35584 9496 35612
rect 9263 35581 9275 35584
rect 9217 35575 9275 35581
rect 9490 35572 9496 35584
rect 9548 35572 9554 35624
rect 10226 35612 10232 35624
rect 10187 35584 10232 35612
rect 10226 35572 10232 35584
rect 10284 35612 10290 35624
rect 10781 35615 10839 35621
rect 10781 35612 10793 35615
rect 10284 35584 10793 35612
rect 10284 35572 10290 35584
rect 10781 35581 10793 35584
rect 10827 35581 10839 35615
rect 10781 35575 10839 35581
rect 11400 35615 11458 35621
rect 11400 35581 11412 35615
rect 11446 35612 11458 35615
rect 12434 35612 12440 35624
rect 11446 35584 12112 35612
rect 12395 35584 12440 35612
rect 11446 35581 11458 35584
rect 11400 35575 11458 35581
rect 6273 35547 6331 35553
rect 6273 35513 6285 35547
rect 6319 35544 6331 35547
rect 7006 35544 7012 35556
rect 6319 35516 7012 35544
rect 6319 35513 6331 35516
rect 6273 35507 6331 35513
rect 7006 35504 7012 35516
rect 7064 35504 7070 35556
rect 7190 35544 7196 35556
rect 7151 35516 7196 35544
rect 7190 35504 7196 35516
rect 7248 35504 7254 35556
rect 7285 35547 7343 35553
rect 7285 35513 7297 35547
rect 7331 35513 7343 35547
rect 7285 35507 7343 35513
rect 6638 35476 6644 35488
rect 6599 35448 6644 35476
rect 6638 35436 6644 35448
rect 6696 35436 6702 35488
rect 7024 35476 7052 35504
rect 7300 35476 7328 35507
rect 12084 35488 12112 35584
rect 12434 35572 12440 35584
rect 12492 35612 12498 35624
rect 12989 35615 13047 35621
rect 12989 35612 13001 35615
rect 12492 35584 13001 35612
rect 12492 35572 12498 35584
rect 12989 35581 13001 35584
rect 13035 35581 13047 35615
rect 12989 35575 13047 35581
rect 8754 35476 8760 35488
rect 7024 35448 7328 35476
rect 8715 35448 8760 35476
rect 8754 35436 8760 35448
rect 8812 35436 8818 35488
rect 9674 35436 9680 35488
rect 9732 35476 9738 35488
rect 9769 35479 9827 35485
rect 9769 35476 9781 35479
rect 9732 35448 9781 35476
rect 9732 35436 9738 35448
rect 9769 35445 9781 35448
rect 9815 35476 9827 35479
rect 10686 35476 10692 35488
rect 9815 35448 10692 35476
rect 9815 35445 9827 35448
rect 9769 35439 9827 35445
rect 10686 35436 10692 35448
rect 10744 35436 10750 35488
rect 11238 35436 11244 35488
rect 11296 35476 11302 35488
rect 11793 35479 11851 35485
rect 11793 35476 11805 35479
rect 11296 35448 11805 35476
rect 11296 35436 11302 35448
rect 11793 35445 11805 35448
rect 11839 35445 11851 35479
rect 11793 35439 11851 35445
rect 12066 35436 12072 35488
rect 12124 35476 12130 35488
rect 12161 35479 12219 35485
rect 12161 35476 12173 35479
rect 12124 35448 12173 35476
rect 12124 35436 12130 35448
rect 12161 35445 12173 35448
rect 12207 35445 12219 35479
rect 12161 35439 12219 35445
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 1762 35232 1768 35284
rect 1820 35272 1826 35284
rect 11701 35275 11759 35281
rect 1820 35244 8651 35272
rect 1820 35232 1826 35244
rect 7006 35204 7012 35216
rect 6967 35176 7012 35204
rect 7006 35164 7012 35176
rect 7064 35164 7070 35216
rect 8623 35148 8651 35244
rect 11701 35241 11713 35275
rect 11747 35272 11759 35275
rect 12802 35272 12808 35284
rect 11747 35244 12808 35272
rect 11747 35241 11759 35244
rect 11701 35235 11759 35241
rect 12802 35232 12808 35244
rect 12860 35232 12866 35284
rect 12897 35275 12955 35281
rect 12897 35241 12909 35275
rect 12943 35272 12955 35275
rect 14090 35272 14096 35284
rect 12943 35244 14096 35272
rect 12943 35241 12955 35244
rect 12897 35235 12955 35241
rect 14090 35232 14096 35244
rect 14148 35232 14154 35284
rect 9858 35164 9864 35216
rect 9916 35204 9922 35216
rect 9953 35207 10011 35213
rect 9953 35204 9965 35207
rect 9916 35176 9965 35204
rect 9916 35164 9922 35176
rect 9953 35173 9965 35176
rect 9999 35173 10011 35207
rect 9953 35167 10011 35173
rect 5880 35139 5938 35145
rect 5880 35105 5892 35139
rect 5926 35136 5938 35139
rect 6178 35136 6184 35148
rect 5926 35108 6184 35136
rect 5926 35105 5938 35108
rect 5880 35099 5938 35105
rect 6178 35096 6184 35108
rect 6236 35096 6242 35148
rect 8570 35136 8576 35148
rect 8628 35145 8651 35148
rect 8628 35139 8666 35145
rect 8518 35108 8576 35136
rect 8570 35096 8576 35108
rect 8654 35105 8666 35139
rect 11514 35136 11520 35148
rect 11475 35108 11520 35136
rect 8628 35099 8666 35105
rect 8628 35096 8634 35099
rect 11514 35096 11520 35108
rect 11572 35096 11578 35148
rect 12710 35136 12716 35148
rect 12671 35108 12716 35136
rect 12710 35096 12716 35108
rect 12768 35096 12774 35148
rect 6917 35071 6975 35077
rect 6917 35068 6929 35071
rect 6656 35040 6929 35068
rect 6656 35009 6684 35040
rect 6917 35037 6929 35040
rect 6963 35037 6975 35071
rect 6917 35031 6975 35037
rect 7561 35071 7619 35077
rect 7561 35037 7573 35071
rect 7607 35068 7619 35071
rect 7926 35068 7932 35080
rect 7607 35040 7932 35068
rect 7607 35037 7619 35040
rect 7561 35031 7619 35037
rect 7926 35028 7932 35040
rect 7984 35028 7990 35080
rect 8711 35071 8769 35077
rect 8711 35037 8723 35071
rect 8757 35068 8769 35071
rect 9398 35068 9404 35080
rect 8757 35040 9404 35068
rect 8757 35037 8769 35040
rect 8711 35031 8769 35037
rect 9398 35028 9404 35040
rect 9456 35068 9462 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9456 35040 9873 35068
rect 9456 35028 9462 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 10502 35068 10508 35080
rect 10463 35040 10508 35068
rect 9861 35031 9919 35037
rect 10502 35028 10508 35040
rect 10560 35028 10566 35080
rect 5951 35003 6009 35009
rect 5951 34969 5963 35003
rect 5997 35000 6009 35003
rect 6641 35003 6699 35009
rect 6641 35000 6653 35003
rect 5997 34972 6653 35000
rect 5997 34969 6009 34972
rect 5951 34963 6009 34969
rect 6641 34969 6653 34972
rect 6687 34969 6699 35003
rect 6641 34963 6699 34969
rect 5258 34932 5264 34944
rect 5219 34904 5264 34932
rect 5258 34892 5264 34904
rect 5316 34892 5322 34944
rect 7190 34892 7196 34944
rect 7248 34932 7254 34944
rect 7837 34935 7895 34941
rect 7837 34932 7849 34935
rect 7248 34904 7849 34932
rect 7248 34892 7254 34904
rect 7837 34901 7849 34904
rect 7883 34901 7895 34935
rect 10870 34932 10876 34944
rect 10831 34904 10876 34932
rect 7837 34895 7895 34901
rect 10870 34892 10876 34904
rect 10928 34892 10934 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 6178 34728 6184 34740
rect 6139 34700 6184 34728
rect 6178 34688 6184 34700
rect 6236 34688 6242 34740
rect 7006 34688 7012 34740
rect 7064 34728 7070 34740
rect 7745 34731 7803 34737
rect 7745 34728 7757 34731
rect 7064 34700 7757 34728
rect 7064 34688 7070 34700
rect 7745 34697 7757 34700
rect 7791 34697 7803 34731
rect 8570 34728 8576 34740
rect 8531 34700 8576 34728
rect 7745 34691 7803 34697
rect 8570 34688 8576 34700
rect 8628 34688 8634 34740
rect 13633 34731 13691 34737
rect 13633 34697 13645 34731
rect 13679 34728 13691 34731
rect 15746 34728 15752 34740
rect 13679 34700 15752 34728
rect 13679 34697 13691 34700
rect 13633 34691 13691 34697
rect 15746 34688 15752 34700
rect 15804 34688 15810 34740
rect 4295 34663 4353 34669
rect 4295 34629 4307 34663
rect 4341 34660 4353 34663
rect 7190 34660 7196 34672
rect 4341 34632 7196 34660
rect 4341 34629 4353 34632
rect 4295 34623 4353 34629
rect 7190 34620 7196 34632
rect 7248 34620 7254 34672
rect 10870 34660 10876 34672
rect 10520 34632 10876 34660
rect 5077 34595 5135 34601
rect 5077 34561 5089 34595
rect 5123 34592 5135 34595
rect 5534 34592 5540 34604
rect 5123 34564 5540 34592
rect 5123 34561 5135 34564
rect 5077 34555 5135 34561
rect 750 34484 756 34536
rect 808 34524 814 34536
rect 4224 34527 4282 34533
rect 4224 34524 4236 34527
rect 808 34496 4236 34524
rect 808 34484 814 34496
rect 4224 34493 4236 34496
rect 4270 34524 4282 34527
rect 4338 34524 4344 34536
rect 4270 34496 4344 34524
rect 4270 34493 4282 34496
rect 4224 34487 4282 34493
rect 4338 34484 4344 34496
rect 4396 34524 4402 34536
rect 5184 34533 5212 34564
rect 5534 34552 5540 34564
rect 5592 34592 5598 34604
rect 7834 34592 7840 34604
rect 5592 34564 7840 34592
rect 5592 34552 5598 34564
rect 7834 34552 7840 34564
rect 7892 34552 7898 34604
rect 8205 34595 8263 34601
rect 8205 34561 8217 34595
rect 8251 34592 8263 34595
rect 8665 34595 8723 34601
rect 8665 34592 8677 34595
rect 8251 34564 8677 34592
rect 8251 34561 8263 34564
rect 8205 34555 8263 34561
rect 8665 34561 8677 34564
rect 8711 34592 8723 34595
rect 8754 34592 8760 34604
rect 8711 34564 8760 34592
rect 8711 34561 8723 34564
rect 8665 34555 8723 34561
rect 8754 34552 8760 34564
rect 8812 34552 8818 34604
rect 10520 34601 10548 34632
rect 10870 34620 10876 34632
rect 10928 34660 10934 34672
rect 12158 34660 12164 34672
rect 10928 34632 12164 34660
rect 10928 34620 10934 34632
rect 12158 34620 12164 34632
rect 12216 34620 12222 34672
rect 10505 34595 10563 34601
rect 10505 34561 10517 34595
rect 10551 34561 10563 34595
rect 10962 34592 10968 34604
rect 10923 34564 10968 34592
rect 10505 34555 10563 34561
rect 10962 34552 10968 34564
rect 11020 34552 11026 34604
rect 12250 34552 12256 34604
rect 12308 34592 12314 34604
rect 12710 34592 12716 34604
rect 12308 34564 12716 34592
rect 12308 34552 12314 34564
rect 4617 34527 4675 34533
rect 4617 34524 4629 34527
rect 4396 34496 4629 34524
rect 4396 34484 4402 34496
rect 4617 34493 4629 34496
rect 4663 34493 4675 34527
rect 4617 34487 4675 34493
rect 5169 34527 5227 34533
rect 5169 34493 5181 34527
rect 5215 34493 5227 34527
rect 5169 34487 5227 34493
rect 5258 34484 5264 34536
rect 5316 34524 5322 34536
rect 5629 34527 5687 34533
rect 5629 34524 5641 34527
rect 5316 34496 5641 34524
rect 5316 34484 5322 34496
rect 5629 34493 5641 34496
rect 5675 34493 5687 34527
rect 5629 34487 5687 34493
rect 5905 34527 5963 34533
rect 5905 34493 5917 34527
rect 5951 34524 5963 34527
rect 6825 34527 6883 34533
rect 6825 34524 6837 34527
rect 5951 34496 6837 34524
rect 5951 34493 5963 34496
rect 5905 34487 5963 34493
rect 6825 34493 6837 34496
rect 6871 34524 6883 34527
rect 7374 34524 7380 34536
rect 6871 34496 7380 34524
rect 6871 34493 6883 34496
rect 6825 34487 6883 34493
rect 7374 34484 7380 34496
rect 7432 34484 7438 34536
rect 12487 34533 12515 34564
rect 12710 34552 12716 34564
rect 12768 34592 12774 34604
rect 12897 34595 12955 34601
rect 12897 34592 12909 34595
rect 12768 34564 12909 34592
rect 12768 34552 12774 34564
rect 12897 34561 12909 34564
rect 12943 34592 12955 34595
rect 13265 34595 13323 34601
rect 13265 34592 13277 34595
rect 12943 34564 13277 34592
rect 12943 34561 12955 34564
rect 12897 34555 12955 34561
rect 13265 34561 13277 34564
rect 13311 34561 13323 34595
rect 13265 34555 13323 34561
rect 12472 34527 12530 34533
rect 12472 34493 12484 34527
rect 12518 34493 12530 34527
rect 12472 34487 12530 34493
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13906 34524 13912 34536
rect 13495 34496 13912 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 13906 34484 13912 34496
rect 13964 34524 13970 34536
rect 14001 34527 14059 34533
rect 14001 34524 14013 34527
rect 13964 34496 14013 34524
rect 13964 34484 13970 34496
rect 14001 34493 14013 34496
rect 14047 34493 14059 34527
rect 14001 34487 14059 34493
rect 6641 34459 6699 34465
rect 6641 34425 6653 34459
rect 6687 34456 6699 34459
rect 6730 34456 6736 34468
rect 6687 34428 6736 34456
rect 6687 34425 6699 34428
rect 6641 34419 6699 34425
rect 6730 34416 6736 34428
rect 6788 34456 6794 34468
rect 7187 34459 7245 34465
rect 7187 34456 7199 34459
rect 6788 34428 7199 34456
rect 6788 34416 6794 34428
rect 7187 34425 7199 34428
rect 7233 34456 7245 34459
rect 9027 34459 9085 34465
rect 9027 34456 9039 34459
rect 7233 34428 9039 34456
rect 7233 34425 7245 34428
rect 7187 34419 7245 34425
rect 9027 34425 9039 34428
rect 9073 34456 9085 34459
rect 10042 34456 10048 34468
rect 9073 34428 10048 34456
rect 9073 34425 9085 34428
rect 9027 34419 9085 34425
rect 10042 34416 10048 34428
rect 10100 34416 10106 34468
rect 10597 34459 10655 34465
rect 10597 34425 10609 34459
rect 10643 34425 10655 34459
rect 10597 34419 10655 34425
rect 9585 34391 9643 34397
rect 9585 34357 9597 34391
rect 9631 34388 9643 34391
rect 9858 34388 9864 34400
rect 9631 34360 9864 34388
rect 9631 34357 9643 34360
rect 9585 34351 9643 34357
rect 9858 34348 9864 34360
rect 9916 34348 9922 34400
rect 10318 34388 10324 34400
rect 10279 34360 10324 34388
rect 10318 34348 10324 34360
rect 10376 34388 10382 34400
rect 10612 34388 10640 34419
rect 11514 34416 11520 34468
rect 11572 34456 11578 34468
rect 11609 34459 11667 34465
rect 11609 34456 11621 34459
rect 11572 34428 11621 34456
rect 11572 34416 11578 34428
rect 11609 34425 11621 34428
rect 11655 34456 11667 34459
rect 12342 34456 12348 34468
rect 11655 34428 12348 34456
rect 11655 34425 11667 34428
rect 11609 34419 11667 34425
rect 12342 34416 12348 34428
rect 12400 34416 12406 34468
rect 10376 34360 10640 34388
rect 10376 34348 10382 34360
rect 11974 34348 11980 34400
rect 12032 34388 12038 34400
rect 12575 34391 12633 34397
rect 12575 34388 12587 34391
rect 12032 34360 12587 34388
rect 12032 34348 12038 34360
rect 12575 34357 12587 34360
rect 12621 34357 12633 34391
rect 12575 34351 12633 34357
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 5350 34184 5356 34196
rect 5311 34156 5356 34184
rect 5350 34144 5356 34156
rect 5408 34144 5414 34196
rect 6178 34184 6184 34196
rect 6139 34156 6184 34184
rect 6178 34144 6184 34156
rect 6236 34144 6242 34196
rect 6638 34144 6644 34196
rect 6696 34184 6702 34196
rect 6733 34187 6791 34193
rect 6733 34184 6745 34187
rect 6696 34156 6745 34184
rect 6696 34144 6702 34156
rect 6733 34153 6745 34156
rect 6779 34153 6791 34187
rect 7006 34184 7012 34196
rect 6967 34156 7012 34184
rect 6733 34147 6791 34153
rect 6748 34116 6776 34147
rect 7006 34144 7012 34156
rect 7064 34144 7070 34196
rect 7374 34184 7380 34196
rect 7335 34156 7380 34184
rect 7374 34144 7380 34156
rect 7432 34144 7438 34196
rect 9398 34184 9404 34196
rect 9359 34156 9404 34184
rect 9398 34144 9404 34156
rect 9456 34144 9462 34196
rect 10042 34184 10048 34196
rect 10003 34156 10048 34184
rect 10042 34144 10048 34156
rect 10100 34144 10106 34196
rect 10597 34187 10655 34193
rect 10597 34153 10609 34187
rect 10643 34184 10655 34187
rect 13541 34187 13599 34193
rect 10643 34156 11652 34184
rect 10643 34153 10655 34156
rect 10597 34147 10655 34153
rect 7745 34119 7803 34125
rect 7745 34116 7757 34119
rect 6748 34088 7757 34116
rect 7745 34085 7757 34088
rect 7791 34116 7803 34119
rect 7834 34116 7840 34128
rect 7791 34088 7840 34116
rect 7791 34085 7803 34088
rect 7745 34079 7803 34085
rect 7834 34076 7840 34088
rect 7892 34076 7898 34128
rect 10502 34076 10508 34128
rect 10560 34116 10566 34128
rect 11514 34116 11520 34128
rect 10560 34088 11520 34116
rect 10560 34076 10566 34088
rect 11514 34076 11520 34088
rect 11572 34076 11578 34128
rect 11624 34125 11652 34156
rect 13541 34153 13553 34187
rect 13587 34184 13599 34187
rect 14734 34184 14740 34196
rect 13587 34156 14740 34184
rect 13587 34153 13599 34156
rect 13541 34147 13599 34153
rect 14734 34144 14740 34156
rect 14792 34144 14798 34196
rect 11609 34119 11667 34125
rect 11609 34085 11621 34119
rect 11655 34116 11667 34119
rect 11698 34116 11704 34128
rect 11655 34088 11704 34116
rect 11655 34085 11667 34088
rect 11609 34079 11667 34085
rect 11698 34076 11704 34088
rect 11756 34076 11762 34128
rect 3510 34008 3516 34060
rect 3568 34048 3574 34060
rect 4798 34048 4804 34060
rect 4856 34057 4862 34060
rect 4856 34051 4894 34057
rect 3568 34020 4804 34048
rect 3568 34008 3574 34020
rect 4798 34008 4804 34020
rect 4882 34017 4894 34051
rect 4856 34011 4894 34017
rect 13357 34051 13415 34057
rect 13357 34017 13369 34051
rect 13403 34048 13415 34051
rect 13538 34048 13544 34060
rect 13403 34020 13544 34048
rect 13403 34017 13415 34020
rect 13357 34011 13415 34017
rect 4856 34008 4862 34011
rect 13538 34008 13544 34020
rect 13596 34008 13602 34060
rect 5810 33980 5816 33992
rect 5771 33952 5816 33980
rect 5810 33940 5816 33952
rect 5868 33940 5874 33992
rect 7653 33983 7711 33989
rect 7653 33949 7665 33983
rect 7699 33949 7711 33983
rect 7926 33980 7932 33992
rect 7887 33952 7932 33980
rect 7653 33943 7711 33949
rect 4939 33915 4997 33921
rect 4939 33881 4951 33915
rect 4985 33912 4997 33915
rect 7668 33912 7696 33943
rect 7926 33940 7932 33952
rect 7984 33940 7990 33992
rect 9677 33983 9735 33989
rect 9677 33949 9689 33983
rect 9723 33980 9735 33983
rect 9766 33980 9772 33992
rect 9723 33952 9772 33980
rect 9723 33949 9735 33952
rect 9677 33943 9735 33949
rect 9766 33940 9772 33952
rect 9824 33940 9830 33992
rect 8846 33912 8852 33924
rect 4985 33884 8852 33912
rect 4985 33881 4997 33884
rect 4939 33875 4997 33881
rect 8846 33872 8852 33884
rect 8904 33872 8910 33924
rect 12066 33912 12072 33924
rect 12027 33884 12072 33912
rect 12066 33872 12072 33884
rect 12124 33872 12130 33924
rect 5626 33844 5632 33856
rect 5587 33816 5632 33844
rect 5626 33804 5632 33816
rect 5684 33804 5690 33856
rect 8662 33844 8668 33856
rect 8623 33816 8668 33844
rect 8662 33804 8668 33816
rect 8720 33804 8726 33856
rect 10686 33804 10692 33856
rect 10744 33844 10750 33856
rect 10873 33847 10931 33853
rect 10873 33844 10885 33847
rect 10744 33816 10885 33844
rect 10744 33804 10750 33816
rect 10873 33813 10885 33816
rect 10919 33813 10931 33847
rect 12526 33844 12532 33856
rect 12487 33816 12532 33844
rect 10873 33807 10931 33813
rect 12526 33804 12532 33816
rect 12584 33804 12590 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 6178 33600 6184 33652
rect 6236 33640 6242 33652
rect 6273 33643 6331 33649
rect 6273 33640 6285 33643
rect 6236 33612 6285 33640
rect 6236 33600 6242 33612
rect 6273 33609 6285 33612
rect 6319 33640 6331 33643
rect 6730 33640 6736 33652
rect 6319 33612 6736 33640
rect 6319 33609 6331 33612
rect 6273 33603 6331 33609
rect 6730 33600 6736 33612
rect 6788 33600 6794 33652
rect 7834 33640 7840 33652
rect 7795 33612 7840 33640
rect 7834 33600 7840 33612
rect 7892 33600 7898 33652
rect 8294 33640 8300 33652
rect 8255 33612 8300 33640
rect 8294 33600 8300 33612
rect 8352 33600 8358 33652
rect 10042 33640 10048 33652
rect 10003 33612 10048 33640
rect 10042 33600 10048 33612
rect 10100 33640 10106 33652
rect 10413 33643 10471 33649
rect 10413 33640 10425 33643
rect 10100 33612 10425 33640
rect 10100 33600 10106 33612
rect 10413 33609 10425 33612
rect 10459 33609 10471 33643
rect 11698 33640 11704 33652
rect 11659 33612 11704 33640
rect 10413 33603 10471 33609
rect 11698 33600 11704 33612
rect 11756 33600 11762 33652
rect 5736 33544 8248 33572
rect 4341 33507 4399 33513
rect 4341 33473 4353 33507
rect 4387 33504 4399 33507
rect 5736 33504 5764 33544
rect 4387 33476 5764 33504
rect 4387 33473 4399 33476
rect 4341 33467 4399 33473
rect 5810 33464 5816 33516
rect 5868 33504 5874 33516
rect 5905 33507 5963 33513
rect 5905 33504 5917 33507
rect 5868 33476 5917 33504
rect 5868 33464 5874 33476
rect 5905 33473 5917 33476
rect 5951 33504 5963 33507
rect 6549 33507 6607 33513
rect 6549 33504 6561 33507
rect 5951 33476 6561 33504
rect 5951 33473 5963 33476
rect 5905 33467 5963 33473
rect 6549 33473 6561 33476
rect 6595 33473 6607 33507
rect 6549 33467 6607 33473
rect 7561 33507 7619 33513
rect 7561 33473 7573 33507
rect 7607 33504 7619 33507
rect 7926 33504 7932 33516
rect 7607 33476 7932 33504
rect 7607 33473 7619 33476
rect 7561 33467 7619 33473
rect 7926 33464 7932 33476
rect 7984 33464 7990 33516
rect 3513 33439 3571 33445
rect 3513 33405 3525 33439
rect 3559 33436 3571 33439
rect 3605 33439 3663 33445
rect 3605 33436 3617 33439
rect 3559 33408 3617 33436
rect 3559 33405 3571 33408
rect 3513 33399 3571 33405
rect 3605 33405 3617 33408
rect 3651 33405 3663 33439
rect 4062 33436 4068 33448
rect 4023 33408 4068 33436
rect 3605 33399 3663 33405
rect 3620 33368 3648 33399
rect 4062 33396 4068 33408
rect 4120 33396 4126 33448
rect 5074 33436 5080 33448
rect 4172 33408 5080 33436
rect 4172 33368 4200 33408
rect 5074 33396 5080 33408
rect 5132 33396 5138 33448
rect 5169 33439 5227 33445
rect 5169 33405 5181 33439
rect 5215 33405 5227 33439
rect 5169 33399 5227 33405
rect 3620 33340 4200 33368
rect 5184 33368 5212 33399
rect 5258 33396 5264 33448
rect 5316 33436 5322 33448
rect 5629 33439 5687 33445
rect 5629 33436 5641 33439
rect 5316 33408 5641 33436
rect 5316 33396 5322 33408
rect 5629 33405 5641 33408
rect 5675 33405 5687 33439
rect 8220 33436 8248 33544
rect 8312 33504 8340 33600
rect 9677 33575 9735 33581
rect 9677 33541 9689 33575
rect 9723 33572 9735 33575
rect 10318 33572 10324 33584
rect 9723 33544 10324 33572
rect 9723 33541 9735 33544
rect 9677 33535 9735 33541
rect 10318 33532 10324 33544
rect 10376 33572 10382 33584
rect 10376 33544 12296 33572
rect 10376 33532 10382 33544
rect 8757 33507 8815 33513
rect 8757 33504 8769 33507
rect 8312 33476 8769 33504
rect 8757 33473 8769 33476
rect 8803 33473 8815 33507
rect 8757 33467 8815 33473
rect 10505 33439 10563 33445
rect 10505 33436 10517 33439
rect 8220 33408 10517 33436
rect 5629 33399 5687 33405
rect 10505 33405 10517 33408
rect 10551 33436 10563 33439
rect 10686 33436 10692 33448
rect 10551 33408 10692 33436
rect 10551 33405 10563 33408
rect 10505 33399 10563 33405
rect 5350 33368 5356 33380
rect 5184 33340 5356 33368
rect 5350 33328 5356 33340
rect 5408 33328 5414 33380
rect 4798 33300 4804 33312
rect 4759 33272 4804 33300
rect 4798 33260 4804 33272
rect 4856 33260 4862 33312
rect 5644 33300 5672 33399
rect 10686 33396 10692 33408
rect 10744 33396 10750 33448
rect 5718 33328 5724 33380
rect 5776 33368 5782 33380
rect 6917 33371 6975 33377
rect 6917 33368 6929 33371
rect 5776 33340 6929 33368
rect 5776 33328 5782 33340
rect 6917 33337 6929 33340
rect 6963 33337 6975 33371
rect 6917 33331 6975 33337
rect 7006 33328 7012 33380
rect 7064 33368 7070 33380
rect 8662 33368 8668 33380
rect 7064 33340 7109 33368
rect 8575 33340 8668 33368
rect 7064 33328 7070 33340
rect 8662 33328 8668 33340
rect 8720 33368 8726 33380
rect 9119 33371 9177 33377
rect 9119 33368 9131 33371
rect 8720 33340 9131 33368
rect 8720 33328 8726 33340
rect 9119 33337 9131 33340
rect 9165 33368 9177 33371
rect 10042 33368 10048 33380
rect 9165 33340 10048 33368
rect 9165 33337 9177 33340
rect 9119 33331 9177 33337
rect 10042 33328 10048 33340
rect 10100 33368 10106 33380
rect 12268 33377 12296 33544
rect 12526 33504 12532 33516
rect 12487 33476 12532 33504
rect 12526 33464 12532 33476
rect 12584 33464 12590 33516
rect 12802 33504 12808 33516
rect 12763 33476 12808 33504
rect 12802 33464 12808 33476
rect 12860 33464 12866 33516
rect 10826 33371 10884 33377
rect 10826 33368 10838 33371
rect 10100 33340 10838 33368
rect 10100 33328 10106 33340
rect 10826 33337 10838 33340
rect 10872 33337 10884 33371
rect 10826 33331 10884 33337
rect 12253 33371 12311 33377
rect 12253 33337 12265 33371
rect 12299 33368 12311 33371
rect 12621 33371 12679 33377
rect 12621 33368 12633 33371
rect 12299 33340 12633 33368
rect 12299 33337 12311 33340
rect 12253 33331 12311 33337
rect 12621 33337 12633 33340
rect 12667 33337 12679 33371
rect 12621 33331 12679 33337
rect 5810 33300 5816 33312
rect 5644 33272 5816 33300
rect 5810 33260 5816 33272
rect 5868 33260 5874 33312
rect 11422 33300 11428 33312
rect 11383 33272 11428 33300
rect 11422 33260 11428 33272
rect 11480 33260 11486 33312
rect 13538 33300 13544 33312
rect 13499 33272 13544 33300
rect 13538 33260 13544 33272
rect 13596 33260 13602 33312
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 3697 33099 3755 33105
rect 3697 33065 3709 33099
rect 3743 33096 3755 33099
rect 4062 33096 4068 33108
rect 3743 33068 4068 33096
rect 3743 33065 3755 33068
rect 3697 33059 3755 33065
rect 4062 33056 4068 33068
rect 4120 33056 4126 33108
rect 4847 33099 4905 33105
rect 4847 33065 4859 33099
rect 4893 33096 4905 33099
rect 5626 33096 5632 33108
rect 4893 33068 5632 33096
rect 4893 33065 4905 33068
rect 4847 33059 4905 33065
rect 5626 33056 5632 33068
rect 5684 33056 5690 33108
rect 8846 33096 8852 33108
rect 8807 33068 8852 33096
rect 8846 33056 8852 33068
rect 8904 33056 8910 33108
rect 11514 33096 11520 33108
rect 11427 33068 11520 33096
rect 11514 33056 11520 33068
rect 11572 33096 11578 33108
rect 11572 33068 12480 33096
rect 11572 33056 11578 33068
rect 6083 33031 6141 33037
rect 6083 32997 6095 33031
rect 6129 33028 6141 33031
rect 6178 33028 6184 33040
rect 6129 33000 6184 33028
rect 6129 32997 6141 33000
rect 6083 32991 6141 32997
rect 6178 32988 6184 33000
rect 6236 32988 6242 33040
rect 8018 33028 8024 33040
rect 7979 33000 8024 33028
rect 8018 32988 8024 33000
rect 8076 32988 8082 33040
rect 10318 33028 10324 33040
rect 10279 33000 10324 33028
rect 10318 32988 10324 33000
rect 10376 32988 10382 33040
rect 10873 33031 10931 33037
rect 10873 32997 10885 33031
rect 10919 33028 10931 33031
rect 10962 33028 10968 33040
rect 10919 33000 10968 33028
rect 10919 32997 10931 33000
rect 10873 32991 10931 32997
rect 10962 32988 10968 33000
rect 11020 32988 11026 33040
rect 11422 32988 11428 33040
rect 11480 33028 11486 33040
rect 11885 33031 11943 33037
rect 11885 33028 11897 33031
rect 11480 33000 11897 33028
rect 11480 32988 11486 33000
rect 11885 32997 11897 33000
rect 11931 32997 11943 33031
rect 11885 32991 11943 32997
rect 12066 32988 12072 33040
rect 12124 33028 12130 33040
rect 12250 33028 12256 33040
rect 12124 33000 12256 33028
rect 12124 32988 12130 33000
rect 12250 32988 12256 33000
rect 12308 32988 12314 33040
rect 12452 33037 12480 33068
rect 12437 33031 12495 33037
rect 12437 32997 12449 33031
rect 12483 33028 12495 33031
rect 12802 33028 12808 33040
rect 12483 33000 12808 33028
rect 12483 32997 12495 33000
rect 12437 32991 12495 32997
rect 12802 32988 12808 33000
rect 12860 32988 12866 33040
rect 4246 32920 4252 32972
rect 4304 32960 4310 32972
rect 4776 32963 4834 32969
rect 4776 32960 4788 32963
rect 4304 32932 4788 32960
rect 4304 32920 4310 32932
rect 4776 32929 4788 32932
rect 4822 32960 4834 32963
rect 5166 32960 5172 32972
rect 4822 32932 5172 32960
rect 4822 32929 4834 32932
rect 4776 32923 4834 32929
rect 5166 32920 5172 32932
rect 5224 32920 5230 32972
rect 13332 32963 13390 32969
rect 13332 32929 13344 32963
rect 13378 32960 13390 32963
rect 13538 32960 13544 32972
rect 13378 32932 13544 32960
rect 13378 32929 13390 32932
rect 13332 32923 13390 32929
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 5074 32852 5080 32904
rect 5132 32892 5138 32904
rect 5261 32895 5319 32901
rect 5261 32892 5273 32895
rect 5132 32864 5273 32892
rect 5132 32852 5138 32864
rect 5261 32861 5273 32864
rect 5307 32892 5319 32895
rect 5626 32892 5632 32904
rect 5307 32864 5632 32892
rect 5307 32861 5319 32864
rect 5261 32855 5319 32861
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32892 5779 32895
rect 5902 32892 5908 32904
rect 5767 32864 5908 32892
rect 5767 32861 5779 32864
rect 5721 32855 5779 32861
rect 5902 32852 5908 32864
rect 5960 32852 5966 32904
rect 7926 32892 7932 32904
rect 7887 32864 7932 32892
rect 7926 32852 7932 32864
rect 7984 32852 7990 32904
rect 8202 32892 8208 32904
rect 8163 32864 8208 32892
rect 8202 32852 8208 32864
rect 8260 32852 8266 32904
rect 9674 32852 9680 32904
rect 9732 32892 9738 32904
rect 10229 32895 10287 32901
rect 10229 32892 10241 32895
rect 9732 32864 10241 32892
rect 9732 32852 9738 32864
rect 10229 32861 10241 32864
rect 10275 32861 10287 32895
rect 10229 32855 10287 32861
rect 11793 32895 11851 32901
rect 11793 32861 11805 32895
rect 11839 32892 11851 32895
rect 12066 32892 12072 32904
rect 11839 32864 12072 32892
rect 11839 32861 11851 32864
rect 11793 32855 11851 32861
rect 12066 32852 12072 32864
rect 12124 32852 12130 32904
rect 4890 32784 4896 32836
rect 4948 32824 4954 32836
rect 8570 32824 8576 32836
rect 4948 32796 8576 32824
rect 4948 32784 4954 32796
rect 8570 32784 8576 32796
rect 8628 32784 8634 32836
rect 5629 32759 5687 32765
rect 5629 32725 5641 32759
rect 5675 32756 5687 32759
rect 5810 32756 5816 32768
rect 5675 32728 5816 32756
rect 5675 32725 5687 32728
rect 5629 32719 5687 32725
rect 5810 32716 5816 32728
rect 5868 32716 5874 32768
rect 6641 32759 6699 32765
rect 6641 32725 6653 32759
rect 6687 32756 6699 32759
rect 7006 32756 7012 32768
rect 6687 32728 7012 32756
rect 6687 32725 6699 32728
rect 6641 32719 6699 32725
rect 7006 32716 7012 32728
rect 7064 32716 7070 32768
rect 7374 32756 7380 32768
rect 7335 32728 7380 32756
rect 7374 32716 7380 32728
rect 7432 32716 7438 32768
rect 9766 32716 9772 32768
rect 9824 32756 9830 32768
rect 9950 32756 9956 32768
rect 9824 32728 9956 32756
rect 9824 32716 9830 32728
rect 9950 32716 9956 32728
rect 10008 32716 10014 32768
rect 10042 32716 10048 32768
rect 10100 32756 10106 32768
rect 13403 32759 13461 32765
rect 13403 32756 13415 32759
rect 10100 32728 13415 32756
rect 10100 32716 10106 32728
rect 13403 32725 13415 32728
rect 13449 32725 13461 32759
rect 13403 32719 13461 32725
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 8018 32512 8024 32564
rect 8076 32552 8082 32564
rect 8297 32555 8355 32561
rect 8297 32552 8309 32555
rect 8076 32524 8309 32552
rect 8076 32512 8082 32524
rect 8297 32521 8309 32524
rect 8343 32552 8355 32555
rect 8573 32555 8631 32561
rect 8573 32552 8585 32555
rect 8343 32524 8585 32552
rect 8343 32521 8355 32524
rect 8297 32515 8355 32521
rect 8573 32521 8585 32524
rect 8619 32521 8631 32555
rect 9858 32552 9864 32564
rect 9819 32524 9864 32552
rect 8573 32515 8631 32521
rect 9858 32512 9864 32524
rect 9916 32512 9922 32564
rect 10318 32512 10324 32564
rect 10376 32552 10382 32564
rect 10965 32555 11023 32561
rect 10965 32552 10977 32555
rect 10376 32524 10977 32552
rect 10376 32512 10382 32524
rect 10965 32521 10977 32524
rect 11011 32552 11023 32555
rect 11422 32552 11428 32564
rect 11011 32524 11428 32552
rect 11011 32521 11023 32524
rect 10965 32515 11023 32521
rect 11422 32512 11428 32524
rect 11480 32552 11486 32564
rect 11701 32555 11759 32561
rect 11701 32552 11713 32555
rect 11480 32524 11713 32552
rect 11480 32512 11486 32524
rect 11701 32521 11713 32524
rect 11747 32521 11759 32555
rect 12066 32552 12072 32564
rect 12027 32524 12072 32552
rect 11701 32515 11759 32521
rect 12066 32512 12072 32524
rect 12124 32512 12130 32564
rect 12158 32512 12164 32564
rect 12216 32552 12222 32564
rect 12575 32555 12633 32561
rect 12575 32552 12587 32555
rect 12216 32524 12587 32552
rect 12216 32512 12222 32524
rect 12575 32521 12587 32524
rect 12621 32521 12633 32555
rect 12575 32515 12633 32521
rect 5077 32487 5135 32493
rect 5077 32453 5089 32487
rect 5123 32484 5135 32487
rect 5166 32484 5172 32496
rect 5123 32456 5172 32484
rect 5123 32453 5135 32456
rect 5077 32447 5135 32453
rect 5166 32444 5172 32456
rect 5224 32484 5230 32496
rect 7558 32484 7564 32496
rect 5224 32456 7564 32484
rect 5224 32444 5230 32456
rect 7558 32444 7564 32456
rect 7616 32444 7622 32496
rect 9674 32444 9680 32496
rect 9732 32484 9738 32496
rect 11333 32487 11391 32493
rect 11333 32484 11345 32487
rect 9732 32456 11345 32484
rect 9732 32444 9738 32456
rect 11333 32453 11345 32456
rect 11379 32453 11391 32487
rect 11333 32447 11391 32453
rect 5810 32416 5816 32428
rect 5736 32388 5816 32416
rect 4246 32357 4252 32360
rect 4224 32351 4252 32357
rect 4224 32348 4236 32351
rect 4159 32320 4236 32348
rect 4224 32317 4236 32320
rect 4304 32348 4310 32360
rect 4617 32351 4675 32357
rect 4617 32348 4629 32351
rect 4304 32320 4629 32348
rect 4224 32311 4252 32317
rect 4246 32308 4252 32311
rect 4304 32308 4310 32320
rect 4617 32317 4629 32320
rect 4663 32317 4675 32351
rect 4617 32311 4675 32317
rect 5445 32351 5503 32357
rect 5445 32317 5457 32351
rect 5491 32348 5503 32351
rect 5626 32348 5632 32360
rect 5491 32320 5632 32348
rect 5491 32317 5503 32320
rect 5445 32311 5503 32317
rect 5626 32308 5632 32320
rect 5684 32308 5690 32360
rect 5736 32357 5764 32388
rect 5810 32376 5816 32388
rect 5868 32416 5874 32428
rect 6549 32419 6607 32425
rect 6549 32416 6561 32419
rect 5868 32388 6561 32416
rect 5868 32376 5874 32388
rect 6549 32385 6561 32388
rect 6595 32385 6607 32419
rect 6549 32379 6607 32385
rect 9493 32419 9551 32425
rect 9493 32385 9505 32419
rect 9539 32416 9551 32419
rect 10042 32416 10048 32428
rect 9539 32388 10048 32416
rect 9539 32385 9551 32388
rect 9493 32379 9551 32385
rect 10042 32376 10048 32388
rect 10100 32376 10106 32428
rect 10689 32419 10747 32425
rect 10689 32385 10701 32419
rect 10735 32416 10747 32419
rect 10962 32416 10968 32428
rect 10735 32388 10968 32416
rect 10735 32385 10747 32388
rect 10689 32379 10747 32385
rect 10962 32376 10968 32388
rect 11020 32376 11026 32428
rect 5721 32351 5779 32357
rect 5721 32317 5733 32351
rect 5767 32317 5779 32351
rect 5721 32311 5779 32317
rect 5994 32308 6000 32360
rect 6052 32348 6058 32360
rect 7374 32348 7380 32360
rect 6052 32320 7380 32348
rect 6052 32308 6058 32320
rect 7374 32308 7380 32320
rect 7432 32308 7438 32360
rect 12158 32308 12164 32360
rect 12216 32348 12222 32360
rect 12472 32351 12530 32357
rect 12472 32348 12484 32351
rect 12216 32320 12484 32348
rect 12216 32308 12222 32320
rect 12472 32317 12484 32320
rect 12518 32348 12530 32351
rect 12897 32351 12955 32357
rect 12897 32348 12909 32351
rect 12518 32320 12909 32348
rect 12518 32317 12530 32320
rect 12472 32311 12530 32317
rect 12897 32317 12909 32320
rect 12943 32317 12955 32351
rect 12897 32311 12955 32317
rect 5902 32280 5908 32292
rect 5863 32252 5908 32280
rect 5902 32240 5908 32252
rect 5960 32240 5966 32292
rect 7698 32283 7756 32289
rect 7698 32249 7710 32283
rect 7744 32249 7756 32283
rect 7698 32243 7756 32249
rect 10137 32283 10195 32289
rect 10137 32249 10149 32283
rect 10183 32249 10195 32283
rect 10137 32243 10195 32249
rect 4295 32215 4353 32221
rect 4295 32181 4307 32215
rect 4341 32212 4353 32215
rect 4522 32212 4528 32224
rect 4341 32184 4528 32212
rect 4341 32181 4353 32184
rect 4295 32175 4353 32181
rect 4522 32172 4528 32184
rect 4580 32172 4586 32224
rect 6178 32172 6184 32224
rect 6236 32212 6242 32224
rect 6273 32215 6331 32221
rect 6273 32212 6285 32215
rect 6236 32184 6285 32212
rect 6236 32172 6242 32184
rect 6273 32181 6285 32184
rect 6319 32212 6331 32215
rect 7098 32212 7104 32224
rect 6319 32184 7104 32212
rect 6319 32181 6331 32184
rect 6273 32175 6331 32181
rect 7098 32172 7104 32184
rect 7156 32212 7162 32224
rect 7193 32215 7251 32221
rect 7193 32212 7205 32215
rect 7156 32184 7205 32212
rect 7156 32172 7162 32184
rect 7193 32181 7205 32184
rect 7239 32212 7251 32215
rect 7713 32212 7741 32243
rect 7239 32184 7741 32212
rect 7239 32181 7251 32184
rect 7193 32175 7251 32181
rect 9858 32172 9864 32224
rect 9916 32212 9922 32224
rect 10152 32212 10180 32243
rect 9916 32184 10180 32212
rect 13357 32215 13415 32221
rect 9916 32172 9922 32184
rect 13357 32181 13369 32215
rect 13403 32212 13415 32215
rect 13538 32212 13544 32224
rect 13403 32184 13544 32212
rect 13403 32181 13415 32184
rect 13357 32175 13415 32181
rect 13538 32172 13544 32184
rect 13596 32172 13602 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 5902 31968 5908 32020
rect 5960 32008 5966 32020
rect 6273 32011 6331 32017
rect 6273 32008 6285 32011
rect 5960 31980 6285 32008
rect 5960 31968 5966 31980
rect 6273 31977 6285 31980
rect 6319 31977 6331 32011
rect 6273 31971 6331 31977
rect 8110 31968 8116 32020
rect 8168 32008 8174 32020
rect 8205 32011 8263 32017
rect 8205 32008 8217 32011
rect 8168 31980 8217 32008
rect 8168 31968 8174 31980
rect 8205 31977 8217 31980
rect 8251 31977 8263 32011
rect 8205 31971 8263 31977
rect 8711 32011 8769 32017
rect 8711 31977 8723 32011
rect 8757 32008 8769 32011
rect 9674 32008 9680 32020
rect 8757 31980 9680 32008
rect 8757 31977 8769 31980
rect 8711 31971 8769 31977
rect 9674 31968 9680 31980
rect 9732 31968 9738 32020
rect 9950 32008 9956 32020
rect 9911 31980 9956 32008
rect 9950 31968 9956 31980
rect 10008 31968 10014 32020
rect 11379 32011 11437 32017
rect 11379 31977 11391 32011
rect 11425 32008 11437 32011
rect 12526 32008 12532 32020
rect 11425 31980 12532 32008
rect 11425 31977 11437 31980
rect 11379 31971 11437 31977
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 566 31900 572 31952
rect 624 31940 630 31952
rect 4203 31943 4261 31949
rect 4203 31940 4215 31943
rect 624 31912 4215 31940
rect 624 31900 630 31912
rect 4203 31909 4215 31912
rect 4249 31909 4261 31943
rect 5994 31940 6000 31952
rect 5955 31912 6000 31940
rect 4203 31903 4261 31909
rect 5994 31900 6000 31912
rect 6052 31900 6058 31952
rect 7006 31940 7012 31952
rect 6967 31912 7012 31940
rect 7006 31900 7012 31912
rect 7064 31900 7070 31952
rect 7561 31943 7619 31949
rect 7561 31909 7573 31943
rect 7607 31940 7619 31943
rect 7837 31943 7895 31949
rect 7837 31940 7849 31943
rect 7607 31912 7849 31940
rect 7607 31909 7619 31912
rect 7561 31903 7619 31909
rect 7837 31909 7849 31912
rect 7883 31940 7895 31943
rect 7926 31940 7932 31952
rect 7883 31912 7932 31940
rect 7883 31909 7895 31912
rect 7837 31903 7895 31909
rect 7926 31900 7932 31912
rect 7984 31900 7990 31952
rect 3970 31872 3976 31884
rect 3931 31844 3976 31872
rect 3970 31832 3976 31844
rect 4028 31832 4034 31884
rect 5537 31875 5595 31881
rect 5537 31841 5549 31875
rect 5583 31872 5595 31875
rect 5626 31872 5632 31884
rect 5583 31844 5632 31872
rect 5583 31841 5595 31844
rect 5537 31835 5595 31841
rect 5626 31832 5632 31844
rect 5684 31832 5690 31884
rect 5810 31872 5816 31884
rect 5771 31844 5816 31872
rect 5810 31832 5816 31844
rect 5868 31832 5874 31884
rect 8481 31875 8539 31881
rect 8481 31841 8493 31875
rect 8527 31872 8539 31875
rect 8570 31872 8576 31884
rect 8527 31844 8576 31872
rect 8527 31841 8539 31844
rect 8481 31835 8539 31841
rect 8570 31832 8576 31844
rect 8628 31832 8634 31884
rect 9674 31872 9680 31884
rect 8817 31844 9680 31872
rect 4522 31764 4528 31816
rect 4580 31804 4586 31816
rect 6546 31804 6552 31816
rect 4580 31776 6552 31804
rect 4580 31764 4586 31776
rect 6546 31764 6552 31776
rect 6604 31804 6610 31816
rect 6917 31807 6975 31813
rect 6917 31804 6929 31807
rect 6604 31776 6929 31804
rect 6604 31764 6610 31776
rect 6917 31773 6929 31776
rect 6963 31773 6975 31807
rect 6917 31767 6975 31773
rect 6730 31696 6736 31748
rect 6788 31736 6794 31748
rect 8817 31736 8845 31844
rect 9674 31832 9680 31844
rect 9732 31832 9738 31884
rect 10137 31875 10195 31881
rect 10137 31841 10149 31875
rect 10183 31841 10195 31875
rect 10137 31835 10195 31841
rect 10152 31804 10180 31835
rect 11146 31832 11152 31884
rect 11204 31872 11210 31884
rect 11241 31875 11299 31881
rect 11241 31872 11253 31875
rect 11204 31844 11253 31872
rect 11204 31832 11210 31844
rect 11241 31841 11253 31844
rect 11287 31872 11299 31875
rect 11330 31872 11336 31884
rect 11287 31844 11336 31872
rect 11287 31841 11299 31844
rect 11241 31835 11299 31841
rect 11330 31832 11336 31844
rect 11388 31832 11394 31884
rect 6788 31708 8845 31736
rect 9508 31776 10180 31804
rect 6788 31696 6794 31708
rect 9508 31680 9536 31776
rect 4154 31628 4160 31680
rect 4212 31668 4218 31680
rect 8478 31668 8484 31680
rect 4212 31640 8484 31668
rect 4212 31628 4218 31640
rect 8478 31628 8484 31640
rect 8536 31668 8542 31680
rect 9033 31671 9091 31677
rect 9033 31668 9045 31671
rect 8536 31640 9045 31668
rect 8536 31628 8542 31640
rect 9033 31637 9045 31640
rect 9079 31668 9091 31671
rect 9490 31668 9496 31680
rect 9079 31640 9496 31668
rect 9079 31637 9091 31640
rect 9033 31631 9091 31637
rect 9490 31628 9496 31640
rect 9548 31628 9554 31680
rect 10781 31671 10839 31677
rect 10781 31637 10793 31671
rect 10827 31668 10839 31671
rect 10870 31668 10876 31680
rect 10827 31640 10876 31668
rect 10827 31637 10839 31640
rect 10781 31631 10839 31637
rect 10870 31628 10876 31640
rect 10928 31628 10934 31680
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 6546 31464 6552 31476
rect 6507 31436 6552 31464
rect 6546 31424 6552 31436
rect 6604 31424 6610 31476
rect 7006 31464 7012 31476
rect 6967 31436 7012 31464
rect 7006 31424 7012 31436
rect 7064 31424 7070 31476
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 10413 31467 10471 31473
rect 10413 31464 10425 31467
rect 9732 31436 10425 31464
rect 9732 31424 9738 31436
rect 10413 31433 10425 31436
rect 10459 31433 10471 31467
rect 10413 31427 10471 31433
rect 8110 31396 8116 31408
rect 7576 31368 8116 31396
rect 7576 31337 7604 31368
rect 8110 31356 8116 31368
rect 8168 31356 8174 31408
rect 7561 31331 7619 31337
rect 7561 31297 7573 31331
rect 7607 31297 7619 31331
rect 8202 31328 8208 31340
rect 8163 31300 8208 31328
rect 7561 31291 7619 31297
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 10781 31331 10839 31337
rect 10781 31297 10793 31331
rect 10827 31328 10839 31331
rect 10962 31328 10968 31340
rect 10827 31300 10968 31328
rect 10827 31297 10839 31300
rect 10781 31291 10839 31297
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 11425 31331 11483 31337
rect 11425 31297 11437 31331
rect 11471 31328 11483 31331
rect 12250 31328 12256 31340
rect 11471 31300 12256 31328
rect 11471 31297 11483 31300
rect 11425 31291 11483 31297
rect 12250 31288 12256 31300
rect 12308 31288 12314 31340
rect 4525 31263 4583 31269
rect 4525 31229 4537 31263
rect 4571 31260 4583 31263
rect 5261 31263 5319 31269
rect 5261 31260 5273 31263
rect 4571 31232 5273 31260
rect 4571 31229 4583 31232
rect 4525 31223 4583 31229
rect 5261 31229 5273 31232
rect 5307 31260 5319 31263
rect 5902 31260 5908 31272
rect 5307 31232 5908 31260
rect 5307 31229 5319 31232
rect 5261 31223 5319 31229
rect 5902 31220 5908 31232
rect 5960 31220 5966 31272
rect 9030 31260 9036 31272
rect 8991 31232 9036 31260
rect 9030 31220 9036 31232
rect 9088 31220 9094 31272
rect 9490 31260 9496 31272
rect 9451 31232 9496 31260
rect 9490 31220 9496 31232
rect 9548 31260 9554 31272
rect 10045 31263 10103 31269
rect 10045 31260 10057 31263
rect 9548 31232 10057 31260
rect 9548 31220 9554 31232
rect 10045 31229 10057 31232
rect 10091 31229 10103 31263
rect 10045 31223 10103 31229
rect 3970 31152 3976 31204
rect 4028 31192 4034 31204
rect 4157 31195 4215 31201
rect 4157 31192 4169 31195
rect 4028 31164 4169 31192
rect 4028 31152 4034 31164
rect 4157 31161 4169 31164
rect 4203 31192 4215 31195
rect 5350 31192 5356 31204
rect 4203 31164 5356 31192
rect 4203 31161 4215 31164
rect 4157 31155 4215 31161
rect 5350 31152 5356 31164
rect 5408 31152 5414 31204
rect 5721 31195 5779 31201
rect 5721 31161 5733 31195
rect 5767 31192 5779 31195
rect 5810 31192 5816 31204
rect 5767 31164 5816 31192
rect 5767 31161 5779 31164
rect 5721 31155 5779 31161
rect 5810 31152 5816 31164
rect 5868 31192 5874 31204
rect 7282 31192 7288 31204
rect 5868 31164 7288 31192
rect 5868 31152 5874 31164
rect 7282 31152 7288 31164
rect 7340 31152 7346 31204
rect 7653 31195 7711 31201
rect 7653 31161 7665 31195
rect 7699 31192 7711 31195
rect 7742 31192 7748 31204
rect 7699 31164 7748 31192
rect 7699 31161 7711 31164
rect 7653 31155 7711 31161
rect 7742 31152 7748 31164
rect 7800 31152 7806 31204
rect 9766 31192 9772 31204
rect 9727 31164 9772 31192
rect 9766 31152 9772 31164
rect 9824 31152 9830 31204
rect 10870 31152 10876 31204
rect 10928 31192 10934 31204
rect 10928 31164 10973 31192
rect 10928 31152 10934 31164
rect 4890 31124 4896 31136
rect 4851 31096 4896 31124
rect 4890 31084 4896 31096
rect 4948 31084 4954 31136
rect 5626 31084 5632 31136
rect 5684 31124 5690 31136
rect 6089 31127 6147 31133
rect 6089 31124 6101 31127
rect 5684 31096 6101 31124
rect 5684 31084 5690 31096
rect 6089 31093 6101 31096
rect 6135 31124 6147 31127
rect 6730 31124 6736 31136
rect 6135 31096 6736 31124
rect 6135 31093 6147 31096
rect 6089 31087 6147 31093
rect 6730 31084 6736 31096
rect 6788 31084 6794 31136
rect 8570 31084 8576 31136
rect 8628 31124 8634 31136
rect 8665 31127 8723 31133
rect 8665 31124 8677 31127
rect 8628 31096 8677 31124
rect 8628 31084 8634 31096
rect 8665 31093 8677 31096
rect 8711 31124 8723 31127
rect 9490 31124 9496 31136
rect 8711 31096 9496 31124
rect 8711 31093 8723 31096
rect 8665 31087 8723 31093
rect 9490 31084 9496 31096
rect 9548 31084 9554 31136
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 11701 31127 11759 31133
rect 11701 31124 11713 31127
rect 11388 31096 11713 31124
rect 11388 31084 11394 31096
rect 11701 31093 11713 31096
rect 11747 31093 11759 31127
rect 11701 31087 11759 31093
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 8294 30880 8300 30932
rect 8352 30920 8358 30932
rect 8754 30920 8760 30932
rect 8352 30892 8760 30920
rect 8352 30880 8358 30892
rect 8754 30880 8760 30892
rect 8812 30880 8818 30932
rect 10042 30920 10048 30932
rect 10003 30892 10048 30920
rect 10042 30880 10048 30892
rect 10100 30880 10106 30932
rect 10597 30923 10655 30929
rect 10597 30889 10609 30923
rect 10643 30920 10655 30923
rect 10870 30920 10876 30932
rect 10643 30892 10876 30920
rect 10643 30889 10655 30892
rect 10597 30883 10655 30889
rect 10870 30880 10876 30892
rect 10928 30880 10934 30932
rect 10962 30880 10968 30932
rect 11020 30920 11026 30932
rect 11020 30892 11065 30920
rect 11020 30880 11026 30892
rect 4801 30855 4859 30861
rect 4801 30821 4813 30855
rect 4847 30852 4859 30855
rect 4890 30852 4896 30864
rect 4847 30824 4896 30852
rect 4847 30821 4859 30824
rect 4801 30815 4859 30821
rect 4890 30812 4896 30824
rect 4948 30812 4954 30864
rect 7834 30852 7840 30864
rect 7795 30824 7840 30852
rect 7834 30812 7840 30824
rect 7892 30812 7898 30864
rect 11606 30852 11612 30864
rect 11567 30824 11612 30852
rect 11606 30812 11612 30824
rect 11664 30812 11670 30864
rect 12161 30855 12219 30861
rect 12161 30821 12173 30855
rect 12207 30852 12219 30855
rect 12250 30852 12256 30864
rect 12207 30824 12256 30852
rect 12207 30821 12219 30824
rect 12161 30815 12219 30821
rect 12250 30812 12256 30824
rect 12308 30812 12314 30864
rect 6086 30744 6092 30796
rect 6144 30784 6150 30796
rect 6273 30787 6331 30793
rect 6273 30784 6285 30787
rect 6144 30756 6285 30784
rect 6144 30744 6150 30756
rect 6273 30753 6285 30756
rect 6319 30753 6331 30787
rect 6454 30784 6460 30796
rect 6415 30756 6460 30784
rect 6273 30747 6331 30753
rect 6454 30744 6460 30756
rect 6512 30784 6518 30796
rect 6914 30784 6920 30796
rect 6512 30756 6920 30784
rect 6512 30744 6518 30756
rect 6914 30744 6920 30756
rect 6972 30744 6978 30796
rect 3970 30676 3976 30728
rect 4028 30716 4034 30728
rect 4709 30719 4767 30725
rect 4709 30716 4721 30719
rect 4028 30688 4721 30716
rect 4028 30676 4034 30688
rect 4709 30685 4721 30688
rect 4755 30685 4767 30719
rect 5350 30716 5356 30728
rect 5311 30688 5356 30716
rect 4709 30679 4767 30685
rect 5350 30676 5356 30688
rect 5408 30676 5414 30728
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30716 7803 30719
rect 8018 30716 8024 30728
rect 7791 30688 8024 30716
rect 7791 30685 7803 30688
rect 7745 30679 7803 30685
rect 8018 30676 8024 30688
rect 8076 30676 8082 30728
rect 8202 30716 8208 30728
rect 8163 30688 8208 30716
rect 8202 30676 8208 30688
rect 8260 30716 8266 30728
rect 8570 30716 8576 30728
rect 8260 30688 8576 30716
rect 8260 30676 8266 30688
rect 8570 30676 8576 30688
rect 8628 30716 8634 30728
rect 8665 30719 8723 30725
rect 8665 30716 8677 30719
rect 8628 30688 8677 30716
rect 8628 30676 8634 30688
rect 8665 30685 8677 30688
rect 8711 30685 8723 30719
rect 8665 30679 8723 30685
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9677 30719 9735 30725
rect 9677 30716 9689 30719
rect 8812 30688 9689 30716
rect 8812 30676 8818 30688
rect 9677 30685 9689 30688
rect 9723 30716 9735 30719
rect 10870 30716 10876 30728
rect 9723 30688 10876 30716
rect 9723 30685 9735 30688
rect 9677 30679 9735 30685
rect 10870 30676 10876 30688
rect 10928 30676 10934 30728
rect 11514 30716 11520 30728
rect 11475 30688 11520 30716
rect 11514 30676 11520 30688
rect 11572 30676 11578 30728
rect 6914 30608 6920 30660
rect 6972 30648 6978 30660
rect 9030 30648 9036 30660
rect 6972 30620 9036 30648
rect 6972 30608 6978 30620
rect 9030 30608 9036 30620
rect 9088 30608 9094 30660
rect 5721 30583 5779 30589
rect 5721 30549 5733 30583
rect 5767 30580 5779 30583
rect 5902 30580 5908 30592
rect 5767 30552 5908 30580
rect 5767 30549 5779 30552
rect 5721 30543 5779 30549
rect 5902 30540 5908 30552
rect 5960 30540 5966 30592
rect 6178 30540 6184 30592
rect 6236 30580 6242 30592
rect 6549 30583 6607 30589
rect 6549 30580 6561 30583
rect 6236 30552 6561 30580
rect 6236 30540 6242 30552
rect 6549 30549 6561 30552
rect 6595 30549 6607 30583
rect 7098 30580 7104 30592
rect 7059 30552 7104 30580
rect 6549 30543 6607 30549
rect 7098 30540 7104 30552
rect 7156 30540 7162 30592
rect 7561 30583 7619 30589
rect 7561 30549 7573 30583
rect 7607 30580 7619 30583
rect 7742 30580 7748 30592
rect 7607 30552 7748 30580
rect 7607 30549 7619 30552
rect 7561 30543 7619 30549
rect 7742 30540 7748 30552
rect 7800 30540 7806 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 3881 30379 3939 30385
rect 3881 30345 3893 30379
rect 3927 30376 3939 30379
rect 3970 30376 3976 30388
rect 3927 30348 3976 30376
rect 3927 30345 3939 30348
rect 3881 30339 3939 30345
rect 3970 30336 3976 30348
rect 4028 30336 4034 30388
rect 4709 30379 4767 30385
rect 4709 30345 4721 30379
rect 4755 30376 4767 30379
rect 4890 30376 4896 30388
rect 4755 30348 4896 30376
rect 4755 30345 4767 30348
rect 4709 30339 4767 30345
rect 4890 30336 4896 30348
rect 4948 30336 4954 30388
rect 7742 30376 7748 30388
rect 7703 30348 7748 30376
rect 7742 30336 7748 30348
rect 7800 30336 7806 30388
rect 8018 30376 8024 30388
rect 7979 30348 8024 30376
rect 8018 30336 8024 30348
rect 8076 30336 8082 30388
rect 8941 30379 8999 30385
rect 8941 30345 8953 30379
rect 8987 30376 8999 30379
rect 9306 30376 9312 30388
rect 8987 30348 9312 30376
rect 8987 30345 8999 30348
rect 8941 30339 8999 30345
rect 9306 30336 9312 30348
rect 9364 30336 9370 30388
rect 10870 30376 10876 30388
rect 10831 30348 10876 30376
rect 10870 30336 10876 30348
rect 10928 30336 10934 30388
rect 11514 30376 11520 30388
rect 11475 30348 11520 30376
rect 11514 30336 11520 30348
rect 11572 30336 11578 30388
rect 3988 30249 4016 30336
rect 10597 30311 10655 30317
rect 10597 30277 10609 30311
rect 10643 30308 10655 30311
rect 11606 30308 11612 30320
rect 10643 30280 11612 30308
rect 10643 30277 10655 30280
rect 10597 30271 10655 30277
rect 11606 30268 11612 30280
rect 11664 30308 11670 30320
rect 11793 30311 11851 30317
rect 11793 30308 11805 30311
rect 11664 30280 11805 30308
rect 11664 30268 11670 30280
rect 11793 30277 11805 30280
rect 11839 30277 11851 30311
rect 11793 30271 11851 30277
rect 3973 30243 4031 30249
rect 3973 30209 3985 30243
rect 4019 30209 4031 30243
rect 5350 30240 5356 30252
rect 5311 30212 5356 30240
rect 3973 30203 4031 30209
rect 5350 30200 5356 30212
rect 5408 30200 5414 30252
rect 9677 30243 9735 30249
rect 9677 30209 9689 30243
rect 9723 30240 9735 30243
rect 9766 30240 9772 30252
rect 9723 30212 9772 30240
rect 9723 30209 9735 30212
rect 9677 30203 9735 30209
rect 9766 30200 9772 30212
rect 9824 30200 9830 30252
rect 6825 30175 6883 30181
rect 6825 30141 6837 30175
rect 6871 30172 6883 30175
rect 7006 30172 7012 30184
rect 6871 30144 7012 30172
rect 6871 30141 6883 30144
rect 6825 30135 6883 30141
rect 7006 30132 7012 30144
rect 7064 30172 7070 30184
rect 8389 30175 8447 30181
rect 8389 30172 8401 30175
rect 7064 30144 8401 30172
rect 7064 30132 7070 30144
rect 8389 30141 8401 30144
rect 8435 30141 8447 30175
rect 8389 30135 8447 30141
rect 8570 30132 8576 30184
rect 8628 30172 8634 30184
rect 8700 30175 8758 30181
rect 8700 30172 8712 30175
rect 8628 30144 8712 30172
rect 8628 30132 8634 30144
rect 8700 30141 8712 30144
rect 8746 30141 8758 30175
rect 8700 30135 8758 30141
rect 5074 30104 5080 30116
rect 5035 30076 5080 30104
rect 5074 30064 5080 30076
rect 5132 30064 5138 30116
rect 5169 30107 5227 30113
rect 5169 30073 5181 30107
rect 5215 30104 5227 30107
rect 5902 30104 5908 30116
rect 5215 30076 5908 30104
rect 5215 30073 5227 30076
rect 5169 30067 5227 30073
rect 5902 30064 5908 30076
rect 5960 30064 5966 30116
rect 6454 30064 6460 30116
rect 6512 30064 6518 30116
rect 7098 30104 7104 30116
rect 7059 30076 7104 30104
rect 7098 30064 7104 30076
rect 7156 30064 7162 30116
rect 10042 30113 10048 30116
rect 9998 30107 10048 30113
rect 9998 30104 10010 30107
rect 9508 30076 10010 30104
rect 6365 30039 6423 30045
rect 6365 30005 6377 30039
rect 6411 30036 6423 30039
rect 6472 30036 6500 30064
rect 7466 30036 7472 30048
rect 6411 30008 7472 30036
rect 6411 30005 6423 30008
rect 6365 29999 6423 30005
rect 7466 29996 7472 30008
rect 7524 29996 7530 30048
rect 8294 29996 8300 30048
rect 8352 30036 8358 30048
rect 9508 30045 9536 30076
rect 9998 30073 10010 30076
rect 10044 30073 10048 30107
rect 9998 30067 10048 30073
rect 10042 30064 10048 30067
rect 10100 30064 10106 30116
rect 9125 30039 9183 30045
rect 9125 30036 9137 30039
rect 8352 30008 9137 30036
rect 8352 29996 8358 30008
rect 9125 30005 9137 30008
rect 9171 30036 9183 30039
rect 9493 30039 9551 30045
rect 9493 30036 9505 30039
rect 9171 30008 9505 30036
rect 9171 30005 9183 30008
rect 9125 29999 9183 30005
rect 9493 30005 9505 30008
rect 9539 30005 9551 30039
rect 9493 29999 9551 30005
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 4617 29835 4675 29841
rect 4617 29801 4629 29835
rect 4663 29832 4675 29835
rect 5074 29832 5080 29844
rect 4663 29804 5080 29832
rect 4663 29801 4675 29804
rect 4617 29795 4675 29801
rect 5074 29792 5080 29804
rect 5132 29832 5138 29844
rect 5350 29832 5356 29844
rect 5132 29804 5356 29832
rect 5132 29792 5138 29804
rect 5350 29792 5356 29804
rect 5408 29792 5414 29844
rect 7561 29835 7619 29841
rect 7561 29801 7573 29835
rect 7607 29832 7619 29835
rect 7834 29832 7840 29844
rect 7607 29804 7840 29832
rect 7607 29801 7619 29804
rect 7561 29795 7619 29801
rect 7834 29792 7840 29804
rect 7892 29792 7898 29844
rect 8018 29792 8024 29844
rect 8076 29832 8082 29844
rect 8389 29835 8447 29841
rect 8389 29832 8401 29835
rect 8076 29804 8401 29832
rect 8076 29792 8082 29804
rect 8389 29801 8401 29804
rect 8435 29801 8447 29835
rect 8389 29795 8447 29801
rect 9493 29835 9551 29841
rect 9493 29801 9505 29835
rect 9539 29832 9551 29835
rect 9766 29832 9772 29844
rect 9539 29804 9772 29832
rect 9539 29801 9551 29804
rect 9493 29795 9551 29801
rect 9766 29792 9772 29804
rect 9824 29792 9830 29844
rect 11241 29835 11299 29841
rect 11241 29801 11253 29835
rect 11287 29832 11299 29835
rect 11514 29832 11520 29844
rect 11287 29804 11520 29832
rect 11287 29801 11299 29804
rect 11241 29795 11299 29801
rect 11514 29792 11520 29804
rect 11572 29792 11578 29844
rect 4062 29724 4068 29776
rect 4120 29764 4126 29776
rect 4893 29767 4951 29773
rect 4893 29764 4905 29767
rect 4120 29736 4905 29764
rect 4120 29724 4126 29736
rect 4893 29733 4905 29736
rect 4939 29733 4951 29767
rect 4893 29727 4951 29733
rect 6546 29724 6552 29776
rect 6604 29764 6610 29776
rect 6962 29767 7020 29773
rect 6962 29764 6974 29767
rect 6604 29736 6974 29764
rect 6604 29724 6610 29736
rect 6962 29733 6974 29736
rect 7008 29764 7020 29767
rect 7098 29764 7104 29776
rect 7008 29736 7104 29764
rect 7008 29733 7020 29736
rect 6962 29727 7020 29733
rect 7098 29724 7104 29736
rect 7156 29724 7162 29776
rect 9861 29767 9919 29773
rect 9861 29733 9873 29767
rect 9907 29764 9919 29767
rect 10042 29764 10048 29776
rect 9907 29736 10048 29764
rect 9907 29733 9919 29736
rect 9861 29727 9919 29733
rect 10042 29724 10048 29736
rect 10100 29724 10106 29776
rect 12434 29724 12440 29776
rect 12492 29724 12498 29776
rect 12250 29696 12256 29708
rect 12211 29668 12256 29696
rect 12250 29656 12256 29668
rect 12308 29696 12314 29708
rect 12452 29696 12480 29724
rect 12308 29668 12480 29696
rect 12308 29656 12314 29668
rect 2869 29631 2927 29637
rect 2869 29597 2881 29631
rect 2915 29628 2927 29631
rect 3050 29628 3056 29640
rect 2915 29600 3056 29628
rect 2915 29597 2927 29600
rect 2869 29591 2927 29597
rect 3050 29588 3056 29600
rect 3108 29588 3114 29640
rect 4614 29588 4620 29640
rect 4672 29628 4678 29640
rect 4801 29631 4859 29637
rect 4801 29628 4813 29631
rect 4672 29600 4813 29628
rect 4672 29588 4678 29600
rect 4801 29597 4813 29600
rect 4847 29597 4859 29631
rect 6638 29628 6644 29640
rect 6599 29600 6644 29628
rect 4801 29591 4859 29597
rect 6638 29588 6644 29600
rect 6696 29588 6702 29640
rect 9766 29628 9772 29640
rect 9727 29600 9772 29628
rect 9766 29588 9772 29600
rect 9824 29588 9830 29640
rect 10413 29631 10471 29637
rect 10413 29597 10425 29631
rect 10459 29628 10471 29631
rect 12434 29628 12440 29640
rect 10459 29600 12440 29628
rect 10459 29597 10471 29600
rect 10413 29591 10471 29597
rect 12434 29588 12440 29600
rect 12492 29588 12498 29640
rect 5350 29560 5356 29572
rect 4126 29532 5028 29560
rect 5311 29532 5356 29560
rect 3099 29495 3157 29501
rect 3099 29461 3111 29495
rect 3145 29492 3157 29495
rect 4126 29492 4154 29532
rect 5000 29504 5028 29532
rect 5350 29520 5356 29532
rect 5408 29520 5414 29572
rect 3145 29464 4154 29492
rect 3145 29461 3157 29464
rect 3099 29455 3157 29461
rect 4982 29452 4988 29504
rect 5040 29492 5046 29504
rect 5721 29495 5779 29501
rect 5721 29492 5733 29495
rect 5040 29464 5733 29492
rect 5040 29452 5046 29464
rect 5721 29461 5733 29464
rect 5767 29461 5779 29495
rect 5721 29455 5779 29461
rect 6086 29452 6092 29504
rect 6144 29492 6150 29504
rect 6273 29495 6331 29501
rect 6273 29492 6285 29495
rect 6144 29464 6285 29492
rect 6144 29452 6150 29464
rect 6273 29461 6285 29464
rect 6319 29461 6331 29495
rect 6273 29455 6331 29461
rect 10410 29452 10416 29504
rect 10468 29492 10474 29504
rect 10689 29495 10747 29501
rect 10689 29492 10701 29495
rect 10468 29464 10701 29492
rect 10468 29452 10474 29464
rect 10689 29461 10701 29464
rect 10735 29461 10747 29495
rect 10689 29455 10747 29461
rect 10778 29452 10784 29504
rect 10836 29492 10842 29504
rect 12391 29495 12449 29501
rect 12391 29492 12403 29495
rect 10836 29464 12403 29492
rect 10836 29452 10842 29464
rect 12391 29461 12403 29464
rect 12437 29461 12449 29495
rect 12391 29455 12449 29461
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 4246 29248 4252 29300
rect 4304 29288 4310 29300
rect 12250 29288 12256 29300
rect 4304 29260 12256 29288
rect 4304 29248 4310 29260
rect 12250 29248 12256 29260
rect 12308 29288 12314 29300
rect 12897 29291 12955 29297
rect 12897 29288 12909 29291
rect 12308 29260 12909 29288
rect 12308 29248 12314 29260
rect 12897 29257 12909 29260
rect 12943 29257 12955 29291
rect 12897 29251 12955 29257
rect 4019 29223 4077 29229
rect 4019 29189 4031 29223
rect 4065 29220 4077 29223
rect 4614 29220 4620 29232
rect 4065 29192 4620 29220
rect 4065 29189 4077 29192
rect 4019 29183 4077 29189
rect 4614 29180 4620 29192
rect 4672 29180 4678 29232
rect 5074 29180 5080 29232
rect 5132 29220 5138 29232
rect 6546 29220 6552 29232
rect 5132 29192 6552 29220
rect 5132 29180 5138 29192
rect 6546 29180 6552 29192
rect 6604 29220 6610 29232
rect 8294 29220 8300 29232
rect 6604 29192 8300 29220
rect 6604 29180 6610 29192
rect 8294 29180 8300 29192
rect 8352 29220 8358 29232
rect 8389 29223 8447 29229
rect 8389 29220 8401 29223
rect 8352 29192 8401 29220
rect 8352 29180 8358 29192
rect 8389 29189 8401 29192
rect 8435 29189 8447 29223
rect 8389 29183 8447 29189
rect 4982 29152 4988 29164
rect 4943 29124 4988 29152
rect 4982 29112 4988 29124
rect 5040 29112 5046 29164
rect 5350 29152 5356 29164
rect 5311 29124 5356 29152
rect 5350 29112 5356 29124
rect 5408 29112 5414 29164
rect 10870 29152 10876 29164
rect 10831 29124 10876 29152
rect 10870 29112 10876 29124
rect 10928 29112 10934 29164
rect 3948 29087 4006 29093
rect 3948 29053 3960 29087
rect 3994 29084 4006 29087
rect 6825 29087 6883 29093
rect 6825 29084 6837 29087
rect 3994 29056 4154 29084
rect 3994 29053 4006 29056
rect 3948 29047 4006 29053
rect 3050 28948 3056 28960
rect 3011 28920 3056 28948
rect 3050 28908 3056 28920
rect 3108 28908 3114 28960
rect 4126 28948 4154 29056
rect 6196 29056 6837 29084
rect 4798 28976 4804 29028
rect 4856 29016 4862 29028
rect 5077 29019 5135 29025
rect 5077 29016 5089 29019
rect 4856 28988 5089 29016
rect 4856 28976 4862 28988
rect 5077 28985 5089 28988
rect 5123 28985 5135 29019
rect 5077 28979 5135 28985
rect 4338 28948 4344 28960
rect 4126 28920 4344 28948
rect 4338 28908 4344 28920
rect 4396 28948 4402 28960
rect 4433 28951 4491 28957
rect 4433 28948 4445 28951
rect 4396 28920 4445 28948
rect 4396 28908 4402 28920
rect 4433 28917 4445 28920
rect 4479 28948 4491 28951
rect 4522 28948 4528 28960
rect 4479 28920 4528 28948
rect 4479 28917 4491 28920
rect 4433 28911 4491 28917
rect 4522 28908 4528 28920
rect 4580 28908 4586 28960
rect 4706 28948 4712 28960
rect 4667 28920 4712 28948
rect 4706 28908 4712 28920
rect 4764 28908 4770 28960
rect 5626 28908 5632 28960
rect 5684 28948 5690 28960
rect 6196 28957 6224 29056
rect 6825 29053 6837 29056
rect 6871 29084 6883 29087
rect 6914 29084 6920 29096
rect 6871 29056 6920 29084
rect 6871 29053 6883 29056
rect 6825 29047 6883 29053
rect 6914 29044 6920 29056
rect 6972 29044 6978 29096
rect 7282 29084 7288 29096
rect 7243 29056 7288 29084
rect 7282 29044 7288 29056
rect 7340 29044 7346 29096
rect 8573 29087 8631 29093
rect 8573 29084 8585 29087
rect 8036 29056 8585 29084
rect 8036 28960 8064 29056
rect 8573 29053 8585 29056
rect 8619 29053 8631 29087
rect 8573 29047 8631 29053
rect 9493 29087 9551 29093
rect 9493 29053 9505 29087
rect 9539 29084 9551 29087
rect 9539 29056 10272 29084
rect 9539 29053 9551 29056
rect 9493 29047 9551 29053
rect 8294 28976 8300 29028
rect 8352 29016 8358 29028
rect 8894 29019 8952 29025
rect 8894 29016 8906 29019
rect 8352 28988 8906 29016
rect 8352 28976 8358 28988
rect 8894 28985 8906 28988
rect 8940 28985 8952 29019
rect 8894 28979 8952 28985
rect 6181 28951 6239 28957
rect 6181 28948 6193 28951
rect 5684 28920 6193 28948
rect 5684 28908 5690 28920
rect 6181 28917 6193 28920
rect 6227 28917 6239 28951
rect 6181 28911 6239 28917
rect 6638 28908 6644 28960
rect 6696 28948 6702 28960
rect 6917 28951 6975 28957
rect 6917 28948 6929 28951
rect 6696 28920 6929 28948
rect 6696 28908 6702 28920
rect 6917 28917 6929 28920
rect 6963 28917 6975 28951
rect 8018 28948 8024 28960
rect 7979 28920 8024 28948
rect 6917 28911 6975 28917
rect 8018 28908 8024 28920
rect 8076 28908 8082 28960
rect 9861 28951 9919 28957
rect 9861 28917 9873 28951
rect 9907 28948 9919 28951
rect 10042 28948 10048 28960
rect 9907 28920 10048 28948
rect 9907 28917 9919 28920
rect 9861 28911 9919 28917
rect 10042 28908 10048 28920
rect 10100 28908 10106 28960
rect 10244 28957 10272 29056
rect 12250 29044 12256 29096
rect 12308 29084 12314 29096
rect 12437 29087 12495 29093
rect 12437 29084 12449 29087
rect 12308 29056 12449 29084
rect 12308 29044 12314 29056
rect 12437 29053 12449 29056
rect 12483 29084 12495 29087
rect 13265 29087 13323 29093
rect 13265 29084 13277 29087
rect 12483 29056 13277 29084
rect 12483 29053 12495 29056
rect 12437 29047 12495 29053
rect 13265 29053 13277 29056
rect 13311 29053 13323 29087
rect 13265 29047 13323 29053
rect 13516 29087 13574 29093
rect 13516 29053 13528 29087
rect 13562 29084 13574 29087
rect 13722 29084 13728 29096
rect 13562 29056 13728 29084
rect 13562 29053 13574 29056
rect 13516 29047 13574 29053
rect 13722 29044 13728 29056
rect 13780 29084 13786 29096
rect 13909 29087 13967 29093
rect 13909 29084 13921 29087
rect 13780 29056 13921 29084
rect 13780 29044 13786 29056
rect 13909 29053 13921 29056
rect 13955 29053 13967 29087
rect 13909 29047 13967 29053
rect 10410 29016 10416 29028
rect 10371 28988 10416 29016
rect 10410 28976 10416 28988
rect 10468 28976 10474 29028
rect 10505 29019 10563 29025
rect 10505 28985 10517 29019
rect 10551 29016 10563 29019
rect 11514 29016 11520 29028
rect 10551 28988 11520 29016
rect 10551 28985 10563 28988
rect 10505 28979 10563 28985
rect 10229 28951 10287 28957
rect 10229 28917 10241 28951
rect 10275 28948 10287 28951
rect 10520 28948 10548 28979
rect 11514 28976 11520 28988
rect 11572 28976 11578 29028
rect 10275 28920 10548 28948
rect 10275 28917 10287 28920
rect 10229 28911 10287 28917
rect 10686 28908 10692 28960
rect 10744 28948 10750 28960
rect 12621 28951 12679 28957
rect 12621 28948 12633 28951
rect 10744 28920 12633 28948
rect 10744 28908 10750 28920
rect 12621 28917 12633 28920
rect 12667 28917 12679 28951
rect 12621 28911 12679 28917
rect 13354 28908 13360 28960
rect 13412 28948 13418 28960
rect 13587 28951 13645 28957
rect 13587 28948 13599 28951
rect 13412 28920 13599 28948
rect 13412 28908 13418 28920
rect 13587 28917 13599 28920
rect 13633 28917 13645 28951
rect 13587 28911 13645 28917
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 4614 28744 4620 28756
rect 4575 28716 4620 28744
rect 4614 28704 4620 28716
rect 4672 28704 4678 28756
rect 6181 28747 6239 28753
rect 6181 28713 6193 28747
rect 6227 28744 6239 28747
rect 6638 28744 6644 28756
rect 6227 28716 6644 28744
rect 6227 28713 6239 28716
rect 6181 28707 6239 28713
rect 6638 28704 6644 28716
rect 6696 28704 6702 28756
rect 9766 28704 9772 28756
rect 9824 28744 9830 28756
rect 9953 28747 10011 28753
rect 9953 28744 9965 28747
rect 9824 28716 9965 28744
rect 9824 28704 9830 28716
rect 9953 28713 9965 28716
rect 9999 28744 10011 28747
rect 13354 28744 13360 28756
rect 9999 28716 13360 28744
rect 9999 28713 10011 28716
rect 9953 28707 10011 28713
rect 13354 28704 13360 28716
rect 13412 28704 13418 28756
rect 4062 28636 4068 28688
rect 4120 28676 4126 28688
rect 4706 28676 4712 28688
rect 4120 28648 4712 28676
rect 4120 28636 4126 28648
rect 4706 28636 4712 28648
rect 4764 28636 4770 28688
rect 7006 28676 7012 28688
rect 6967 28648 7012 28676
rect 7006 28636 7012 28648
rect 7064 28636 7070 28688
rect 8754 28676 8760 28688
rect 8715 28648 8760 28676
rect 8754 28636 8760 28648
rect 8812 28636 8818 28688
rect 10321 28679 10379 28685
rect 10321 28645 10333 28679
rect 10367 28676 10379 28679
rect 11146 28676 11152 28688
rect 10367 28648 11152 28676
rect 10367 28645 10379 28648
rect 10321 28639 10379 28645
rect 11146 28636 11152 28648
rect 11204 28676 11210 28688
rect 11885 28679 11943 28685
rect 11885 28676 11897 28679
rect 11204 28648 11897 28676
rect 11204 28636 11210 28648
rect 11885 28645 11897 28648
rect 11931 28645 11943 28679
rect 12434 28676 12440 28688
rect 12395 28648 12440 28676
rect 11885 28639 11943 28645
rect 12434 28636 12440 28648
rect 12492 28636 12498 28688
rect 4798 28608 4804 28620
rect 4759 28580 4804 28608
rect 4798 28568 4804 28580
rect 4856 28608 4862 28620
rect 5721 28611 5779 28617
rect 5721 28608 5733 28611
rect 4856 28580 5733 28608
rect 4856 28568 4862 28580
rect 5721 28577 5733 28580
rect 5767 28577 5779 28611
rect 5721 28571 5779 28577
rect 6549 28611 6607 28617
rect 6549 28577 6561 28611
rect 6595 28577 6607 28611
rect 6549 28571 6607 28577
rect 6270 28500 6276 28552
rect 6328 28540 6334 28552
rect 6564 28540 6592 28571
rect 6638 28568 6644 28620
rect 6696 28608 6702 28620
rect 6733 28611 6791 28617
rect 6733 28608 6745 28611
rect 6696 28580 6745 28608
rect 6696 28568 6702 28580
rect 6733 28577 6745 28580
rect 6779 28608 6791 28611
rect 7282 28608 7288 28620
rect 6779 28580 7288 28608
rect 6779 28577 6791 28580
rect 6733 28571 6791 28577
rect 7282 28568 7288 28580
rect 7340 28568 7346 28620
rect 8110 28608 8116 28620
rect 8071 28580 8116 28608
rect 8110 28568 8116 28580
rect 8168 28568 8174 28620
rect 8478 28608 8484 28620
rect 8439 28580 8484 28608
rect 8478 28568 8484 28580
rect 8536 28568 8542 28620
rect 10870 28568 10876 28620
rect 10928 28608 10934 28620
rect 13262 28608 13268 28620
rect 10928 28580 10973 28608
rect 13223 28580 13268 28608
rect 10928 28568 10934 28580
rect 13262 28568 13268 28580
rect 13320 28568 13326 28620
rect 8128 28540 8156 28568
rect 6328 28512 8156 28540
rect 10229 28543 10287 28549
rect 6328 28500 6334 28512
rect 10229 28509 10241 28543
rect 10275 28540 10287 28543
rect 10318 28540 10324 28552
rect 10275 28512 10324 28540
rect 10275 28509 10287 28512
rect 10229 28503 10287 28509
rect 10318 28500 10324 28512
rect 10376 28500 10382 28552
rect 11793 28543 11851 28549
rect 11793 28509 11805 28543
rect 11839 28540 11851 28543
rect 11839 28512 12664 28540
rect 11839 28509 11851 28512
rect 11793 28503 11851 28509
rect 12636 28416 12664 28512
rect 12618 28364 12624 28416
rect 12676 28404 12682 28416
rect 13403 28407 13461 28413
rect 13403 28404 13415 28407
rect 12676 28376 13415 28404
rect 12676 28364 12682 28376
rect 13403 28373 13415 28376
rect 13449 28373 13461 28407
rect 13403 28367 13461 28373
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 4525 28203 4583 28209
rect 4525 28169 4537 28203
rect 4571 28200 4583 28203
rect 4798 28200 4804 28212
rect 4571 28172 4804 28200
rect 4571 28169 4583 28172
rect 4525 28163 4583 28169
rect 4798 28160 4804 28172
rect 4856 28200 4862 28212
rect 5905 28203 5963 28209
rect 5905 28200 5917 28203
rect 4856 28172 5917 28200
rect 4856 28160 4862 28172
rect 5905 28169 5917 28172
rect 5951 28169 5963 28203
rect 6270 28200 6276 28212
rect 6231 28172 6276 28200
rect 5905 28163 5963 28169
rect 6270 28160 6276 28172
rect 6328 28160 6334 28212
rect 8294 28200 8300 28212
rect 8255 28172 8300 28200
rect 8294 28160 8300 28172
rect 8352 28160 8358 28212
rect 8478 28160 8484 28212
rect 8536 28200 8542 28212
rect 9677 28203 9735 28209
rect 9677 28200 9689 28203
rect 8536 28172 9689 28200
rect 8536 28160 8542 28172
rect 9677 28169 9689 28172
rect 9723 28200 9735 28203
rect 10686 28200 10692 28212
rect 9723 28172 10692 28200
rect 9723 28169 9735 28172
rect 9677 28163 9735 28169
rect 10686 28160 10692 28172
rect 10744 28160 10750 28212
rect 11146 28200 11152 28212
rect 11107 28172 11152 28200
rect 11146 28160 11152 28172
rect 11204 28200 11210 28212
rect 11425 28203 11483 28209
rect 11425 28200 11437 28203
rect 11204 28172 11437 28200
rect 11204 28160 11210 28172
rect 11425 28169 11437 28172
rect 11471 28200 11483 28203
rect 11793 28203 11851 28209
rect 11793 28200 11805 28203
rect 11471 28172 11805 28200
rect 11471 28169 11483 28172
rect 11425 28163 11483 28169
rect 11793 28169 11805 28172
rect 11839 28169 11851 28203
rect 11793 28163 11851 28169
rect 12342 28160 12348 28212
rect 12400 28200 12406 28212
rect 13262 28200 13268 28212
rect 12400 28172 13268 28200
rect 12400 28160 12406 28172
rect 13262 28160 13268 28172
rect 13320 28200 13326 28212
rect 13633 28203 13691 28209
rect 13633 28200 13645 28203
rect 13320 28172 13645 28200
rect 13320 28160 13326 28172
rect 13633 28169 13645 28172
rect 13679 28169 13691 28203
rect 13633 28163 13691 28169
rect 4062 28092 4068 28144
rect 4120 28132 4126 28144
rect 6086 28132 6092 28144
rect 4120 28104 6092 28132
rect 4120 28092 4126 28104
rect 6086 28092 6092 28104
rect 6144 28092 6150 28144
rect 7466 28092 7472 28144
rect 7524 28132 7530 28144
rect 7524 28104 10364 28132
rect 7524 28092 7530 28104
rect 4080 28064 4108 28092
rect 3712 28036 4108 28064
rect 3712 28005 3740 28036
rect 5534 28024 5540 28076
rect 5592 28064 5598 28076
rect 6549 28067 6607 28073
rect 6549 28064 6561 28067
rect 5592 28036 6561 28064
rect 5592 28024 5598 28036
rect 6549 28033 6561 28036
rect 6595 28064 6607 28067
rect 8021 28067 8079 28073
rect 6595 28036 6960 28064
rect 6595 28033 6607 28036
rect 6549 28027 6607 28033
rect 3697 27999 3755 28005
rect 3697 27965 3709 27999
rect 3743 27965 3755 27999
rect 3697 27959 3755 27965
rect 3789 27999 3847 28005
rect 3789 27965 3801 27999
rect 3835 27996 3847 27999
rect 3970 27996 3976 28008
rect 3835 27968 3976 27996
rect 3835 27965 3847 27968
rect 3789 27959 3847 27965
rect 3970 27956 3976 27968
rect 4028 27956 4034 28008
rect 4157 27999 4215 28005
rect 4157 27965 4169 27999
rect 4203 27996 4215 27999
rect 4982 27996 4988 28008
rect 4203 27968 4237 27996
rect 4943 27968 4988 27996
rect 4203 27965 4215 27968
rect 4157 27959 4215 27965
rect 3329 27931 3387 27937
rect 3329 27897 3341 27931
rect 3375 27928 3387 27931
rect 4172 27928 4200 27959
rect 4982 27956 4988 27968
rect 5040 27956 5046 28008
rect 5074 27956 5080 28008
rect 5132 27996 5138 28008
rect 6932 28005 6960 28036
rect 8021 28033 8033 28067
rect 8067 28064 8079 28067
rect 8110 28064 8116 28076
rect 8067 28036 8116 28064
rect 8067 28033 8079 28036
rect 8021 28027 8079 28033
rect 8110 28024 8116 28036
rect 8168 28064 8174 28076
rect 9674 28064 9680 28076
rect 8168 28036 9680 28064
rect 8168 28024 8174 28036
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 6917 27999 6975 28005
rect 5132 27968 5349 27996
rect 5132 27956 5138 27968
rect 5321 27937 5349 27968
rect 6917 27965 6929 27999
rect 6963 27996 6975 27999
rect 7190 27996 7196 28008
rect 6963 27968 7196 27996
rect 6963 27965 6975 27968
rect 6917 27959 6975 27965
rect 7190 27956 7196 27968
rect 7248 27956 7254 28008
rect 7469 27999 7527 28005
rect 7469 27965 7481 27999
rect 7515 27965 7527 27999
rect 7469 27959 7527 27965
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27996 7711 27999
rect 8478 27996 8484 28008
rect 7699 27968 8484 27996
rect 7699 27965 7711 27968
rect 7653 27959 7711 27965
rect 5306 27931 5364 27937
rect 3375 27900 5212 27928
rect 3375 27897 3387 27900
rect 3329 27891 3387 27897
rect 4893 27863 4951 27869
rect 4893 27829 4905 27863
rect 4939 27860 4951 27863
rect 5074 27860 5080 27872
rect 4939 27832 5080 27860
rect 4939 27829 4951 27832
rect 4893 27823 4951 27829
rect 5074 27820 5080 27832
rect 5132 27820 5138 27872
rect 5184 27860 5212 27900
rect 5306 27897 5318 27931
rect 5352 27897 5364 27931
rect 5306 27891 5364 27897
rect 7006 27888 7012 27940
rect 7064 27928 7070 27940
rect 7484 27928 7512 27959
rect 8478 27956 8484 27968
rect 8536 27956 8542 28008
rect 9401 27999 9459 28005
rect 8680 27968 8846 27996
rect 8570 27928 8576 27940
rect 7064 27900 8576 27928
rect 7064 27888 7070 27900
rect 8570 27888 8576 27900
rect 8628 27888 8634 27940
rect 7466 27860 7472 27872
rect 5184 27832 7472 27860
rect 7466 27820 7472 27832
rect 7524 27820 7530 27872
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 8680 27860 8708 27968
rect 8818 27940 8846 27968
rect 9401 27965 9413 27999
rect 9447 27996 9459 27999
rect 10042 27996 10048 28008
rect 9447 27968 10048 27996
rect 9447 27965 9459 27968
rect 9401 27959 9459 27965
rect 10042 27956 10048 27968
rect 10100 27956 10106 28008
rect 10226 27996 10232 28008
rect 10187 27968 10232 27996
rect 10226 27956 10232 27968
rect 10284 27956 10290 28008
rect 10336 27996 10364 28104
rect 12621 27999 12679 28005
rect 12621 27996 12633 27999
rect 10336 27968 12633 27996
rect 12621 27965 12633 27968
rect 12667 27996 12679 27999
rect 13357 27999 13415 28005
rect 13357 27996 13369 27999
rect 12667 27968 13369 27996
rect 12667 27965 12679 27968
rect 12621 27959 12679 27965
rect 13357 27965 13369 27968
rect 13403 27965 13415 27999
rect 13357 27959 13415 27965
rect 8818 27937 8852 27940
rect 8803 27931 8852 27937
rect 8803 27897 8815 27931
rect 8849 27897 8852 27931
rect 8803 27891 8852 27897
rect 8846 27888 8852 27891
rect 8904 27928 8910 27940
rect 9858 27928 9864 27940
rect 8904 27900 9864 27928
rect 8904 27888 8910 27900
rect 9858 27888 9864 27900
rect 9916 27928 9922 27940
rect 10594 27937 10600 27940
rect 10591 27928 10600 27937
rect 9916 27900 10088 27928
rect 10555 27900 10600 27928
rect 9916 27888 9922 27900
rect 10060 27869 10088 27900
rect 10591 27891 10600 27900
rect 10594 27888 10600 27891
rect 10652 27888 10658 27940
rect 12437 27931 12495 27937
rect 12437 27897 12449 27931
rect 12483 27897 12495 27931
rect 12437 27891 12495 27897
rect 8352 27832 8708 27860
rect 10045 27863 10103 27869
rect 8352 27820 8358 27832
rect 10045 27829 10057 27863
rect 10091 27829 10103 27863
rect 10045 27823 10103 27829
rect 10502 27820 10508 27872
rect 10560 27860 10566 27872
rect 12161 27863 12219 27869
rect 12161 27860 12173 27863
rect 10560 27832 12173 27860
rect 10560 27820 10566 27832
rect 12161 27829 12173 27832
rect 12207 27860 12219 27863
rect 12452 27860 12480 27891
rect 12710 27860 12716 27872
rect 12207 27832 12480 27860
rect 12671 27832 12716 27860
rect 12207 27829 12219 27832
rect 12161 27823 12219 27829
rect 12710 27820 12716 27832
rect 12768 27820 12774 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 4709 27659 4767 27665
rect 4709 27625 4721 27659
rect 4755 27656 4767 27659
rect 4982 27656 4988 27668
rect 4755 27628 4988 27656
rect 4755 27625 4767 27628
rect 4709 27619 4767 27625
rect 4982 27616 4988 27628
rect 5040 27656 5046 27668
rect 5261 27659 5319 27665
rect 5261 27656 5273 27659
rect 5040 27628 5273 27656
rect 5040 27616 5046 27628
rect 5261 27625 5273 27628
rect 5307 27625 5319 27659
rect 7006 27656 7012 27668
rect 6967 27628 7012 27656
rect 5261 27619 5319 27625
rect 7006 27616 7012 27628
rect 7064 27616 7070 27668
rect 8018 27656 8024 27668
rect 7979 27628 8024 27656
rect 8018 27616 8024 27628
rect 8076 27616 8082 27668
rect 8478 27616 8484 27668
rect 8536 27656 8542 27668
rect 8941 27659 8999 27665
rect 8941 27656 8953 27659
rect 8536 27628 8953 27656
rect 8536 27616 8542 27628
rect 8941 27625 8953 27628
rect 8987 27625 8999 27659
rect 8941 27619 8999 27625
rect 10410 27616 10416 27668
rect 10468 27656 10474 27668
rect 12618 27656 12624 27668
rect 10468 27628 12480 27656
rect 12579 27628 12624 27656
rect 10468 27616 10474 27628
rect 6178 27588 6184 27600
rect 4172 27560 6184 27588
rect 4172 27532 4200 27560
rect 6178 27548 6184 27560
rect 6236 27548 6242 27600
rect 10042 27548 10048 27600
rect 10100 27588 10106 27600
rect 10137 27591 10195 27597
rect 10137 27588 10149 27591
rect 10100 27560 10149 27588
rect 10100 27548 10106 27560
rect 10137 27557 10149 27560
rect 10183 27557 10195 27591
rect 10137 27551 10195 27557
rect 10689 27591 10747 27597
rect 10689 27557 10701 27591
rect 10735 27588 10747 27591
rect 10870 27588 10876 27600
rect 10735 27560 10876 27588
rect 10735 27557 10747 27560
rect 10689 27551 10747 27557
rect 10870 27548 10876 27560
rect 10928 27588 10934 27600
rect 11333 27591 11391 27597
rect 11333 27588 11345 27591
rect 10928 27560 11345 27588
rect 10928 27548 10934 27560
rect 11333 27557 11345 27560
rect 11379 27557 11391 27591
rect 11698 27588 11704 27600
rect 11659 27560 11704 27588
rect 11333 27551 11391 27557
rect 11698 27548 11704 27560
rect 11756 27548 11762 27600
rect 12452 27588 12480 27628
rect 12618 27616 12624 27628
rect 12676 27616 12682 27668
rect 13219 27591 13277 27597
rect 13219 27588 13231 27591
rect 12452 27560 13231 27588
rect 13219 27557 13231 27560
rect 13265 27557 13277 27591
rect 13219 27551 13277 27557
rect 3513 27523 3571 27529
rect 3513 27489 3525 27523
rect 3559 27520 3571 27523
rect 4062 27520 4068 27532
rect 3559 27492 4068 27520
rect 3559 27489 3571 27492
rect 3513 27483 3571 27489
rect 4062 27480 4068 27492
rect 4120 27480 4126 27532
rect 4154 27480 4160 27532
rect 4212 27520 4218 27532
rect 5445 27523 5503 27529
rect 4212 27492 4305 27520
rect 4212 27480 4218 27492
rect 5445 27489 5457 27523
rect 5491 27520 5503 27523
rect 5534 27520 5540 27532
rect 5491 27492 5540 27520
rect 5491 27489 5503 27492
rect 5445 27483 5503 27489
rect 5534 27480 5540 27492
rect 5592 27480 5598 27532
rect 5629 27523 5687 27529
rect 5629 27489 5641 27523
rect 5675 27489 5687 27523
rect 5994 27520 6000 27532
rect 5955 27492 6000 27520
rect 5629 27483 5687 27489
rect 5644 27452 5672 27483
rect 5994 27480 6000 27492
rect 6052 27480 6058 27532
rect 7926 27520 7932 27532
rect 7887 27492 7932 27520
rect 7926 27480 7932 27492
rect 7984 27480 7990 27532
rect 8481 27523 8539 27529
rect 8481 27489 8493 27523
rect 8527 27520 8539 27523
rect 8570 27520 8576 27532
rect 8527 27492 8576 27520
rect 8527 27489 8539 27492
rect 8481 27483 8539 27489
rect 8570 27480 8576 27492
rect 8628 27480 8634 27532
rect 12253 27523 12311 27529
rect 12253 27489 12265 27523
rect 12299 27520 12311 27523
rect 12434 27520 12440 27532
rect 12299 27492 12440 27520
rect 12299 27489 12311 27492
rect 12253 27483 12311 27489
rect 12434 27480 12440 27492
rect 12492 27480 12498 27532
rect 13078 27520 13084 27532
rect 13039 27492 13084 27520
rect 13078 27480 13084 27492
rect 13136 27480 13142 27532
rect 6178 27452 6184 27464
rect 5552 27424 6184 27452
rect 4341 27387 4399 27393
rect 4341 27353 4353 27387
rect 4387 27384 4399 27387
rect 5552 27384 5580 27424
rect 6178 27412 6184 27424
rect 6236 27412 6242 27464
rect 10045 27455 10103 27461
rect 10045 27421 10057 27455
rect 10091 27452 10103 27455
rect 10134 27452 10140 27464
rect 10091 27424 10140 27452
rect 10091 27421 10103 27424
rect 10045 27415 10103 27421
rect 10134 27412 10140 27424
rect 10192 27452 10198 27464
rect 10778 27452 10784 27464
rect 10192 27424 10784 27452
rect 10192 27412 10198 27424
rect 10778 27412 10784 27424
rect 10836 27412 10842 27464
rect 11606 27452 11612 27464
rect 11567 27424 11612 27452
rect 11606 27412 11612 27424
rect 11664 27412 11670 27464
rect 4387 27356 5580 27384
rect 4387 27353 4399 27356
rect 4341 27347 4399 27353
rect 10226 27344 10232 27396
rect 10284 27384 10290 27396
rect 10965 27387 11023 27393
rect 10965 27384 10977 27387
rect 10284 27356 10977 27384
rect 10284 27344 10290 27356
rect 10965 27353 10977 27356
rect 11011 27353 11023 27387
rect 10965 27347 11023 27353
rect 5074 27316 5080 27328
rect 5035 27288 5080 27316
rect 5074 27276 5080 27288
rect 5132 27276 5138 27328
rect 6638 27316 6644 27328
rect 6599 27288 6644 27316
rect 6638 27276 6644 27288
rect 6696 27276 6702 27328
rect 9493 27319 9551 27325
rect 9493 27285 9505 27319
rect 9539 27316 9551 27319
rect 10318 27316 10324 27328
rect 9539 27288 10324 27316
rect 9539 27285 9551 27288
rect 9493 27279 9551 27285
rect 10318 27276 10324 27288
rect 10376 27316 10382 27328
rect 11790 27316 11796 27328
rect 10376 27288 11796 27316
rect 10376 27276 10382 27288
rect 11790 27276 11796 27288
rect 11848 27276 11854 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 4154 27072 4160 27124
rect 4212 27112 4218 27124
rect 5902 27112 5908 27124
rect 4212 27084 4257 27112
rect 5863 27084 5908 27112
rect 4212 27072 4218 27084
rect 5902 27072 5908 27084
rect 5960 27072 5966 27124
rect 6178 27112 6184 27124
rect 6139 27084 6184 27112
rect 6178 27072 6184 27084
rect 6236 27072 6242 27124
rect 6638 27072 6644 27124
rect 6696 27112 6702 27124
rect 7009 27115 7067 27121
rect 7009 27112 7021 27115
rect 6696 27084 7021 27112
rect 6696 27072 6702 27084
rect 7009 27081 7021 27084
rect 7055 27081 7067 27115
rect 10042 27112 10048 27124
rect 10003 27084 10048 27112
rect 7009 27075 7067 27081
rect 10042 27072 10048 27084
rect 10100 27072 10106 27124
rect 11609 27115 11667 27121
rect 11609 27081 11621 27115
rect 11655 27112 11667 27115
rect 11698 27112 11704 27124
rect 11655 27084 11704 27112
rect 11655 27081 11667 27084
rect 11609 27075 11667 27081
rect 11698 27072 11704 27084
rect 11756 27072 11762 27124
rect 11790 27072 11796 27124
rect 11848 27112 11854 27124
rect 12575 27115 12633 27121
rect 12575 27112 12587 27115
rect 11848 27084 12587 27112
rect 11848 27072 11854 27084
rect 12575 27081 12587 27084
rect 12621 27081 12633 27115
rect 13078 27112 13084 27124
rect 13039 27084 13084 27112
rect 12575 27075 12633 27081
rect 13078 27072 13084 27084
rect 13136 27072 13142 27124
rect 5442 27004 5448 27056
rect 5500 27044 5506 27056
rect 7377 27047 7435 27053
rect 7377 27044 7389 27047
rect 5500 27016 7389 27044
rect 5500 27004 5506 27016
rect 7377 27013 7389 27016
rect 7423 27044 7435 27047
rect 7926 27044 7932 27056
rect 7423 27016 7932 27044
rect 7423 27013 7435 27016
rect 7377 27007 7435 27013
rect 7926 27004 7932 27016
rect 7984 27004 7990 27056
rect 11238 27004 11244 27056
rect 11296 27044 11302 27056
rect 12802 27044 12808 27056
rect 11296 27016 12808 27044
rect 11296 27004 11302 27016
rect 12802 27004 12808 27016
rect 12860 27004 12866 27056
rect 4706 26936 4712 26988
rect 4764 26976 4770 26988
rect 4893 26979 4951 26985
rect 4893 26976 4905 26979
rect 4764 26948 4905 26976
rect 4764 26936 4770 26948
rect 4893 26945 4905 26948
rect 4939 26976 4951 26979
rect 5994 26976 6000 26988
rect 4939 26948 6000 26976
rect 4939 26945 4951 26948
rect 4893 26939 4951 26945
rect 5994 26936 6000 26948
rect 6052 26976 6058 26988
rect 7282 26976 7288 26988
rect 6052 26948 7288 26976
rect 6052 26936 6058 26948
rect 7282 26936 7288 26948
rect 7340 26936 7346 26988
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26976 8723 26979
rect 10226 26976 10232 26988
rect 8711 26948 10232 26976
rect 8711 26945 8723 26948
rect 8665 26939 8723 26945
rect 10226 26936 10232 26948
rect 10284 26936 10290 26988
rect 10505 26979 10563 26985
rect 10505 26945 10517 26979
rect 10551 26976 10563 26979
rect 10870 26976 10876 26988
rect 10551 26948 10876 26976
rect 10551 26945 10563 26948
rect 10505 26939 10563 26945
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 12066 26936 12072 26988
rect 12124 26976 12130 26988
rect 12161 26979 12219 26985
rect 12161 26976 12173 26979
rect 12124 26948 12173 26976
rect 12124 26936 12130 26948
rect 12161 26945 12173 26948
rect 12207 26976 12219 26979
rect 12207 26948 12515 26976
rect 12207 26945 12219 26948
rect 12161 26939 12219 26945
rect 4982 26908 4988 26920
rect 4943 26880 4988 26908
rect 4982 26868 4988 26880
rect 5040 26868 5046 26920
rect 12487 26917 12515 26948
rect 6825 26911 6883 26917
rect 6825 26877 6837 26911
rect 6871 26877 6883 26911
rect 7929 26911 7987 26917
rect 7929 26908 7941 26911
rect 6825 26871 6883 26877
rect 7852 26880 7941 26908
rect 5074 26800 5080 26852
rect 5132 26840 5138 26852
rect 5306 26843 5364 26849
rect 5306 26840 5318 26843
rect 5132 26812 5318 26840
rect 5132 26800 5138 26812
rect 5306 26809 5318 26812
rect 5352 26809 5364 26843
rect 5306 26803 5364 26809
rect 6086 26800 6092 26852
rect 6144 26840 6150 26852
rect 6549 26843 6607 26849
rect 6549 26840 6561 26843
rect 6144 26812 6561 26840
rect 6144 26800 6150 26812
rect 6549 26809 6561 26812
rect 6595 26840 6607 26843
rect 6840 26840 6868 26871
rect 6595 26812 6868 26840
rect 6595 26809 6607 26812
rect 6549 26803 6607 26809
rect 7852 26784 7880 26880
rect 7929 26877 7941 26880
rect 7975 26877 7987 26911
rect 7929 26871 7987 26877
rect 8481 26911 8539 26917
rect 8481 26877 8493 26911
rect 8527 26908 8539 26911
rect 12472 26911 12530 26917
rect 8527 26880 8616 26908
rect 8527 26877 8539 26880
rect 8481 26871 8539 26877
rect 8588 26784 8616 26880
rect 12472 26877 12484 26911
rect 12518 26877 12530 26911
rect 12472 26871 12530 26877
rect 10594 26800 10600 26852
rect 10652 26840 10658 26852
rect 11149 26843 11207 26849
rect 10652 26812 10697 26840
rect 10652 26800 10658 26812
rect 11149 26809 11161 26843
rect 11195 26840 11207 26843
rect 11238 26840 11244 26852
rect 11195 26812 11244 26840
rect 11195 26809 11207 26812
rect 11149 26803 11207 26809
rect 11238 26800 11244 26812
rect 11296 26800 11302 26852
rect 5718 26732 5724 26784
rect 5776 26772 5782 26784
rect 7834 26772 7840 26784
rect 5776 26744 7840 26772
rect 5776 26732 5782 26744
rect 7834 26732 7840 26744
rect 7892 26732 7898 26784
rect 8570 26732 8576 26784
rect 8628 26772 8634 26784
rect 8941 26775 8999 26781
rect 8941 26772 8953 26775
rect 8628 26744 8953 26772
rect 8628 26732 8634 26744
rect 8941 26741 8953 26744
rect 8987 26772 8999 26775
rect 9309 26775 9367 26781
rect 9309 26772 9321 26775
rect 8987 26744 9321 26772
rect 8987 26741 8999 26744
rect 8941 26735 8999 26741
rect 9309 26741 9321 26744
rect 9355 26741 9367 26775
rect 9309 26735 9367 26741
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 10045 26571 10103 26577
rect 10045 26537 10057 26571
rect 10091 26568 10103 26571
rect 10134 26568 10140 26580
rect 10091 26540 10140 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 10134 26528 10140 26540
rect 10192 26528 10198 26580
rect 10413 26571 10471 26577
rect 10413 26537 10425 26571
rect 10459 26568 10471 26571
rect 10594 26568 10600 26580
rect 10459 26540 10600 26568
rect 10459 26537 10471 26540
rect 10413 26531 10471 26537
rect 10594 26528 10600 26540
rect 10652 26528 10658 26580
rect 10962 26528 10968 26580
rect 11020 26568 11026 26580
rect 11514 26568 11520 26580
rect 11020 26540 11422 26568
rect 11475 26540 11520 26568
rect 11020 26528 11026 26540
rect 4062 26460 4068 26512
rect 4120 26500 4126 26512
rect 4801 26503 4859 26509
rect 4801 26500 4813 26503
rect 4120 26472 4813 26500
rect 4120 26460 4126 26472
rect 4801 26469 4813 26472
rect 4847 26469 4859 26503
rect 8386 26500 8392 26512
rect 4801 26463 4859 26469
rect 4908 26472 8392 26500
rect 4908 26444 4936 26472
rect 8386 26460 8392 26472
rect 8444 26500 8450 26512
rect 10318 26500 10324 26512
rect 8444 26472 10324 26500
rect 8444 26460 8450 26472
rect 10318 26460 10324 26472
rect 10376 26460 10382 26512
rect 10686 26500 10692 26512
rect 10647 26472 10692 26500
rect 10686 26460 10692 26472
rect 10744 26460 10750 26512
rect 11238 26500 11244 26512
rect 11199 26472 11244 26500
rect 11238 26460 11244 26472
rect 11296 26460 11302 26512
rect 11394 26500 11422 26540
rect 11514 26528 11520 26540
rect 11572 26568 11578 26580
rect 12207 26571 12265 26577
rect 12207 26568 12219 26571
rect 11572 26540 12219 26568
rect 11572 26528 11578 26540
rect 12207 26537 12219 26540
rect 12253 26537 12265 26571
rect 12207 26531 12265 26537
rect 11394 26472 11514 26500
rect 4890 26432 4896 26444
rect 4851 26404 4896 26432
rect 4890 26392 4896 26404
rect 4948 26392 4954 26444
rect 6454 26392 6460 26444
rect 6512 26432 6518 26444
rect 6914 26432 6920 26444
rect 6512 26404 6920 26432
rect 6512 26392 6518 26404
rect 6914 26392 6920 26404
rect 6972 26432 6978 26444
rect 7009 26435 7067 26441
rect 7009 26432 7021 26435
rect 6972 26404 7021 26432
rect 6972 26392 6978 26404
rect 7009 26401 7021 26404
rect 7055 26432 7067 26435
rect 7374 26432 7380 26444
rect 7055 26404 7380 26432
rect 7055 26401 7067 26404
rect 7009 26395 7067 26401
rect 7374 26392 7380 26404
rect 7432 26392 7438 26444
rect 8018 26432 8024 26444
rect 7979 26404 8024 26432
rect 8018 26392 8024 26404
rect 8076 26392 8082 26444
rect 8570 26432 8576 26444
rect 8531 26404 8576 26432
rect 8570 26392 8576 26404
rect 8628 26392 8634 26444
rect 11486 26432 11514 26472
rect 12066 26432 12072 26444
rect 12124 26441 12130 26444
rect 12124 26435 12162 26441
rect 11486 26404 12072 26432
rect 12066 26392 12072 26404
rect 12150 26401 12162 26435
rect 12124 26395 12162 26401
rect 12124 26392 12130 26395
rect 7098 26364 7104 26376
rect 7059 26336 7104 26364
rect 7098 26324 7104 26336
rect 7156 26324 7162 26376
rect 7837 26367 7895 26373
rect 7837 26333 7849 26367
rect 7883 26364 7895 26367
rect 8588 26364 8616 26392
rect 8754 26364 8760 26376
rect 7883 26336 8616 26364
rect 8715 26336 8760 26364
rect 7883 26333 7895 26336
rect 7837 26327 7895 26333
rect 8754 26324 8760 26336
rect 8812 26324 8818 26376
rect 10597 26367 10655 26373
rect 10597 26333 10609 26367
rect 10643 26364 10655 26367
rect 10778 26364 10784 26376
rect 10643 26336 10784 26364
rect 10643 26333 10655 26336
rect 10597 26327 10655 26333
rect 10778 26324 10784 26336
rect 10836 26324 10842 26376
rect 7558 26256 7564 26308
rect 7616 26296 7622 26308
rect 8386 26296 8392 26308
rect 7616 26268 8392 26296
rect 7616 26256 7622 26268
rect 8386 26256 8392 26268
rect 8444 26256 8450 26308
rect 4709 26231 4767 26237
rect 4709 26197 4721 26231
rect 4755 26228 4767 26231
rect 4982 26228 4988 26240
rect 4755 26200 4988 26228
rect 4755 26197 4767 26200
rect 4709 26191 4767 26197
rect 4982 26188 4988 26200
rect 5040 26228 5046 26240
rect 5350 26228 5356 26240
rect 5040 26200 5356 26228
rect 5040 26188 5046 26200
rect 5350 26188 5356 26200
rect 5408 26188 5414 26240
rect 5534 26188 5540 26240
rect 5592 26228 5598 26240
rect 5813 26231 5871 26237
rect 5813 26228 5825 26231
rect 5592 26200 5825 26228
rect 5592 26188 5598 26200
rect 5813 26197 5825 26200
rect 5859 26197 5871 26231
rect 9306 26228 9312 26240
rect 9267 26200 9312 26228
rect 5813 26191 5871 26197
rect 9306 26188 9312 26200
rect 9364 26188 9370 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 4890 26024 4896 26036
rect 4851 25996 4896 26024
rect 4890 25984 4896 25996
rect 4948 25984 4954 26036
rect 6454 26024 6460 26036
rect 6415 25996 6460 26024
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 8846 25984 8852 26036
rect 8904 26024 8910 26036
rect 9033 26027 9091 26033
rect 9033 26024 9045 26027
rect 8904 25996 9045 26024
rect 8904 25984 8910 25996
rect 9033 25993 9045 25996
rect 9079 26024 9091 26027
rect 9125 26027 9183 26033
rect 9125 26024 9137 26027
rect 9079 25996 9137 26024
rect 9079 25993 9091 25996
rect 9033 25987 9091 25993
rect 9125 25993 9137 25996
rect 9171 25993 9183 26027
rect 9125 25987 9183 25993
rect 10229 26027 10287 26033
rect 10229 25993 10241 26027
rect 10275 26024 10287 26027
rect 10594 26024 10600 26036
rect 10275 25996 10600 26024
rect 10275 25993 10287 25996
rect 10229 25987 10287 25993
rect 10594 25984 10600 25996
rect 10652 25984 10658 26036
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 10873 26027 10931 26033
rect 10873 26024 10885 26027
rect 10744 25996 10885 26024
rect 10744 25984 10750 25996
rect 10873 25993 10885 25996
rect 10919 25993 10931 26027
rect 10873 25987 10931 25993
rect 11471 26027 11529 26033
rect 11471 25993 11483 26027
rect 11517 26024 11529 26027
rect 11974 26024 11980 26036
rect 11517 25996 11980 26024
rect 11517 25993 11529 25996
rect 11471 25987 11529 25993
rect 11974 25984 11980 25996
rect 12032 25984 12038 26036
rect 12066 25984 12072 26036
rect 12124 26024 12130 26036
rect 12124 25996 12169 26024
rect 12124 25984 12130 25996
rect 5905 25891 5963 25897
rect 5905 25857 5917 25891
rect 5951 25888 5963 25891
rect 6086 25888 6092 25900
rect 5951 25860 6092 25888
rect 5951 25857 5963 25860
rect 5905 25851 5963 25857
rect 6086 25848 6092 25860
rect 6144 25848 6150 25900
rect 4525 25823 4583 25829
rect 4525 25789 4537 25823
rect 4571 25820 4583 25823
rect 5534 25820 5540 25832
rect 4571 25792 5540 25820
rect 4571 25789 4583 25792
rect 4525 25783 4583 25789
rect 5534 25780 5540 25792
rect 5592 25780 5598 25832
rect 7745 25823 7803 25829
rect 7745 25789 7757 25823
rect 7791 25789 7803 25823
rect 7745 25783 7803 25789
rect 8297 25823 8355 25829
rect 8297 25789 8309 25823
rect 8343 25820 8355 25823
rect 9306 25820 9312 25832
rect 8343 25792 8432 25820
rect 9219 25792 9312 25820
rect 8343 25789 8355 25792
rect 8297 25783 8355 25789
rect 5353 25755 5411 25761
rect 5353 25752 5365 25755
rect 5184 25724 5365 25752
rect 5074 25644 5080 25696
rect 5132 25684 5138 25696
rect 5184 25693 5212 25724
rect 5353 25721 5365 25724
rect 5399 25721 5411 25755
rect 5353 25715 5411 25721
rect 5626 25712 5632 25764
rect 5684 25752 5690 25764
rect 7561 25755 7619 25761
rect 7561 25752 7573 25755
rect 5684 25724 7573 25752
rect 5684 25712 5690 25724
rect 7561 25721 7573 25724
rect 7607 25752 7619 25755
rect 7760 25752 7788 25783
rect 7607 25724 7788 25752
rect 7607 25721 7619 25724
rect 7561 25715 7619 25721
rect 5169 25687 5227 25693
rect 5169 25684 5181 25687
rect 5132 25656 5181 25684
rect 5132 25644 5138 25656
rect 5169 25653 5181 25656
rect 5215 25653 5227 25687
rect 8404 25684 8432 25792
rect 9306 25780 9312 25792
rect 9364 25820 9370 25832
rect 9766 25820 9772 25832
rect 9364 25792 9772 25820
rect 9364 25780 9370 25792
rect 9766 25780 9772 25792
rect 9824 25780 9830 25832
rect 11238 25780 11244 25832
rect 11296 25820 11302 25832
rect 11368 25823 11426 25829
rect 11368 25820 11380 25823
rect 11296 25792 11380 25820
rect 11296 25780 11302 25792
rect 11368 25789 11380 25792
rect 11414 25789 11426 25823
rect 11368 25783 11426 25789
rect 8481 25755 8539 25761
rect 8481 25721 8493 25755
rect 8527 25752 8539 25755
rect 9398 25752 9404 25764
rect 8527 25724 9404 25752
rect 8527 25721 8539 25724
rect 8481 25715 8539 25721
rect 9398 25712 9404 25724
rect 9456 25712 9462 25764
rect 9631 25755 9689 25761
rect 9631 25721 9643 25755
rect 9677 25721 9689 25755
rect 9631 25715 9689 25721
rect 8570 25684 8576 25696
rect 8404 25656 8576 25684
rect 5169 25647 5227 25653
rect 8570 25644 8576 25656
rect 8628 25684 8634 25696
rect 8757 25687 8815 25693
rect 8757 25684 8769 25687
rect 8628 25656 8769 25684
rect 8628 25644 8634 25656
rect 8757 25653 8769 25656
rect 8803 25653 8815 25687
rect 8757 25647 8815 25653
rect 9033 25687 9091 25693
rect 9033 25653 9045 25687
rect 9079 25684 9091 25687
rect 9646 25684 9674 25715
rect 10042 25684 10048 25696
rect 9079 25656 10048 25684
rect 9079 25653 9091 25656
rect 9033 25647 9091 25653
rect 10042 25644 10048 25656
rect 10100 25644 10106 25696
rect 10597 25687 10655 25693
rect 10597 25653 10609 25687
rect 10643 25684 10655 25687
rect 10778 25684 10784 25696
rect 10643 25656 10784 25684
rect 10643 25653 10655 25656
rect 10597 25647 10655 25653
rect 10778 25644 10784 25656
rect 10836 25644 10842 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 5350 25480 5356 25492
rect 5311 25452 5356 25480
rect 5350 25440 5356 25452
rect 5408 25440 5414 25492
rect 5994 25440 6000 25492
rect 6052 25480 6058 25492
rect 6641 25483 6699 25489
rect 6641 25480 6653 25483
rect 6052 25452 6653 25480
rect 6052 25440 6058 25452
rect 6641 25449 6653 25452
rect 6687 25449 6699 25483
rect 7098 25480 7104 25492
rect 7059 25452 7104 25480
rect 6641 25443 6699 25449
rect 7098 25440 7104 25452
rect 7156 25440 7162 25492
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 9033 25483 9091 25489
rect 9033 25480 9045 25483
rect 8812 25452 9045 25480
rect 8812 25440 8818 25452
rect 9033 25449 9045 25452
rect 9079 25449 9091 25483
rect 9398 25480 9404 25492
rect 9359 25452 9404 25480
rect 9033 25443 9091 25449
rect 9398 25440 9404 25452
rect 9456 25440 9462 25492
rect 10042 25480 10048 25492
rect 10003 25452 10048 25480
rect 10042 25440 10048 25452
rect 10100 25440 10106 25492
rect 10597 25483 10655 25489
rect 10597 25449 10609 25483
rect 10643 25480 10655 25483
rect 10686 25480 10692 25492
rect 10643 25452 10692 25480
rect 10643 25449 10655 25452
rect 10597 25443 10655 25449
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 10778 25440 10784 25492
rect 10836 25480 10842 25492
rect 11425 25483 11483 25489
rect 11425 25480 11437 25483
rect 10836 25452 11437 25480
rect 10836 25440 10842 25452
rect 11425 25449 11437 25452
rect 11471 25449 11483 25483
rect 11425 25443 11483 25449
rect 5169 25415 5227 25421
rect 5169 25381 5181 25415
rect 5215 25412 5227 25415
rect 5215 25384 6132 25412
rect 5215 25381 5227 25384
rect 5169 25375 5227 25381
rect 6104 25356 6132 25384
rect 5534 25344 5540 25356
rect 5447 25316 5540 25344
rect 5534 25304 5540 25316
rect 5592 25344 5598 25356
rect 5902 25344 5908 25356
rect 5592 25316 5908 25344
rect 5592 25304 5598 25316
rect 5902 25304 5908 25316
rect 5960 25304 5966 25356
rect 6086 25344 6092 25356
rect 5999 25316 6092 25344
rect 6086 25304 6092 25316
rect 6144 25344 6150 25356
rect 7193 25347 7251 25353
rect 7193 25344 7205 25347
rect 6144 25316 7205 25344
rect 6144 25304 6150 25316
rect 7193 25313 7205 25316
rect 7239 25313 7251 25347
rect 7193 25307 7251 25313
rect 7282 25304 7288 25356
rect 7340 25344 7346 25356
rect 9416 25344 9444 25440
rect 11238 25372 11244 25424
rect 11296 25412 11302 25424
rect 11885 25415 11943 25421
rect 11885 25412 11897 25415
rect 11296 25384 11897 25412
rect 11296 25372 11302 25384
rect 11885 25381 11897 25384
rect 11931 25381 11943 25415
rect 11885 25375 11943 25381
rect 9677 25347 9735 25353
rect 9677 25344 9689 25347
rect 7340 25316 7385 25344
rect 9416 25316 9689 25344
rect 7340 25304 7346 25316
rect 9677 25313 9689 25316
rect 9723 25313 9735 25347
rect 9677 25307 9735 25313
rect 10870 25304 10876 25356
rect 10928 25344 10934 25356
rect 10965 25347 11023 25353
rect 10965 25344 10977 25347
rect 10928 25316 10977 25344
rect 10928 25304 10934 25316
rect 10965 25313 10977 25316
rect 11011 25344 11023 25347
rect 12434 25344 12440 25356
rect 11011 25316 12440 25344
rect 11011 25313 11023 25316
rect 10965 25307 11023 25313
rect 12434 25304 12440 25316
rect 12492 25304 12498 25356
rect 6178 25276 6184 25288
rect 6139 25248 6184 25276
rect 6178 25236 6184 25248
rect 6236 25236 6242 25288
rect 4430 25140 4436 25152
rect 4391 25112 4436 25140
rect 4430 25100 4436 25112
rect 4488 25100 4494 25152
rect 4801 25143 4859 25149
rect 4801 25109 4813 25143
rect 4847 25140 4859 25143
rect 5166 25140 5172 25152
rect 4847 25112 5172 25140
rect 4847 25109 4859 25112
rect 4801 25103 4859 25109
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 8018 25140 8024 25152
rect 6788 25112 8024 25140
rect 6788 25100 6794 25112
rect 8018 25100 8024 25112
rect 8076 25140 8082 25152
rect 8205 25143 8263 25149
rect 8205 25140 8217 25143
rect 8076 25112 8217 25140
rect 8076 25100 8082 25112
rect 8205 25109 8217 25112
rect 8251 25109 8263 25143
rect 8205 25103 8263 25109
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 4430 24896 4436 24948
rect 4488 24936 4494 24948
rect 5445 24939 5503 24945
rect 5445 24936 5457 24939
rect 4488 24908 5457 24936
rect 4488 24896 4494 24908
rect 5445 24905 5457 24908
rect 5491 24936 5503 24939
rect 7653 24939 7711 24945
rect 5491 24908 7328 24936
rect 5491 24905 5503 24908
rect 5445 24899 5503 24905
rect 7098 24828 7104 24880
rect 7156 24877 7162 24880
rect 7300 24877 7328 24908
rect 7653 24905 7665 24939
rect 7699 24936 7711 24939
rect 12250 24936 12256 24948
rect 7699 24908 12256 24936
rect 7699 24905 7711 24908
rect 7653 24899 7711 24905
rect 12250 24896 12256 24908
rect 12308 24896 12314 24948
rect 7156 24871 7205 24877
rect 7156 24837 7159 24871
rect 7193 24837 7205 24871
rect 7156 24831 7205 24837
rect 7285 24871 7343 24877
rect 7285 24837 7297 24871
rect 7331 24868 7343 24871
rect 8478 24868 8484 24880
rect 7331 24840 8484 24868
rect 7331 24837 7343 24840
rect 7285 24831 7343 24837
rect 7156 24828 7162 24831
rect 8478 24828 8484 24840
rect 8536 24828 8542 24880
rect 8846 24868 8852 24880
rect 8807 24840 8852 24868
rect 8846 24828 8852 24840
rect 8904 24868 8910 24880
rect 8904 24840 9536 24868
rect 8904 24828 8910 24840
rect 4798 24800 4804 24812
rect 3804 24772 4804 24800
rect 3804 24673 3832 24772
rect 4798 24760 4804 24772
rect 4856 24760 4862 24812
rect 5077 24803 5135 24809
rect 5077 24769 5089 24803
rect 5123 24800 5135 24803
rect 5537 24803 5595 24809
rect 5537 24800 5549 24803
rect 5123 24772 5549 24800
rect 5123 24769 5135 24772
rect 5077 24763 5135 24769
rect 5537 24769 5549 24772
rect 5583 24800 5595 24803
rect 6641 24803 6699 24809
rect 6641 24800 6653 24803
rect 5583 24772 6653 24800
rect 5583 24769 5595 24772
rect 5537 24763 5595 24769
rect 6641 24769 6653 24772
rect 6687 24800 6699 24803
rect 7006 24800 7012 24812
rect 6687 24772 7012 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 7006 24760 7012 24772
rect 7064 24800 7070 24812
rect 7377 24803 7435 24809
rect 7377 24800 7389 24803
rect 7064 24772 7389 24800
rect 7064 24760 7070 24772
rect 7377 24769 7389 24772
rect 7423 24769 7435 24803
rect 7377 24763 7435 24769
rect 8754 24760 8760 24812
rect 8812 24800 8818 24812
rect 9033 24803 9091 24809
rect 9033 24800 9045 24803
rect 8812 24772 9045 24800
rect 8812 24760 8818 24772
rect 9033 24769 9045 24772
rect 9079 24769 9091 24803
rect 9033 24763 9091 24769
rect 3970 24732 3976 24744
rect 3931 24704 3976 24732
rect 3970 24692 3976 24704
rect 4028 24692 4034 24744
rect 5350 24741 5356 24744
rect 5316 24735 5356 24741
rect 5316 24701 5328 24735
rect 5316 24695 5356 24701
rect 5350 24692 5356 24695
rect 5408 24692 5414 24744
rect 5442 24692 5448 24744
rect 5500 24732 5506 24744
rect 6730 24732 6736 24744
rect 5500 24704 6736 24732
rect 5500 24692 5506 24704
rect 6730 24692 6736 24704
rect 6788 24692 6794 24744
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7340 24704 8033 24732
rect 7340 24692 7346 24704
rect 8021 24701 8033 24704
rect 8067 24701 8079 24735
rect 8021 24695 8079 24701
rect 3789 24667 3847 24673
rect 3789 24633 3801 24667
rect 3835 24633 3847 24667
rect 3789 24627 3847 24633
rect 3142 24556 3148 24608
rect 3200 24596 3206 24608
rect 3605 24599 3663 24605
rect 3605 24596 3617 24599
rect 3200 24568 3617 24596
rect 3200 24556 3206 24568
rect 3605 24565 3617 24568
rect 3651 24596 3663 24599
rect 3804 24596 3832 24627
rect 3651 24568 3832 24596
rect 3988 24596 4016 24692
rect 4338 24664 4344 24676
rect 4299 24636 4344 24664
rect 4338 24624 4344 24636
rect 4396 24624 4402 24676
rect 5166 24664 5172 24676
rect 5127 24636 5172 24664
rect 5166 24624 5172 24636
rect 5224 24624 5230 24676
rect 5902 24664 5908 24676
rect 5863 24636 5908 24664
rect 5902 24624 5908 24636
rect 5960 24624 5966 24676
rect 6273 24667 6331 24673
rect 6273 24633 6285 24667
rect 6319 24664 6331 24667
rect 7009 24667 7067 24673
rect 7009 24664 7021 24667
rect 6319 24636 7021 24664
rect 6319 24633 6331 24636
rect 6273 24627 6331 24633
rect 7009 24633 7021 24636
rect 7055 24664 7067 24667
rect 8938 24664 8944 24676
rect 7055 24636 8944 24664
rect 7055 24633 7067 24636
rect 7009 24627 7067 24633
rect 4709 24599 4767 24605
rect 4709 24596 4721 24599
rect 3988 24568 4721 24596
rect 3651 24565 3663 24568
rect 3605 24559 3663 24565
rect 4709 24565 4721 24568
rect 4755 24596 4767 24599
rect 5074 24596 5080 24608
rect 4755 24568 5080 24596
rect 4755 24565 4767 24568
rect 4709 24559 4767 24565
rect 5074 24556 5080 24568
rect 5132 24596 5138 24608
rect 6288 24596 6316 24627
rect 8938 24624 8944 24636
rect 8996 24624 9002 24676
rect 9398 24673 9404 24676
rect 9395 24664 9404 24673
rect 9311 24636 9404 24664
rect 9395 24627 9404 24636
rect 9456 24664 9462 24676
rect 9508 24664 9536 24840
rect 10870 24800 10876 24812
rect 10831 24772 10876 24800
rect 10870 24760 10876 24772
rect 10928 24760 10934 24812
rect 11238 24800 11244 24812
rect 11199 24772 11244 24800
rect 11238 24760 11244 24772
rect 11296 24760 11302 24812
rect 9953 24735 10011 24741
rect 9953 24701 9965 24735
rect 9999 24732 10011 24735
rect 10597 24735 10655 24741
rect 10597 24732 10609 24735
rect 9999 24704 10609 24732
rect 9999 24701 10011 24704
rect 9953 24695 10011 24701
rect 10597 24701 10609 24704
rect 10643 24701 10655 24735
rect 10597 24695 10655 24701
rect 10229 24667 10287 24673
rect 10229 24664 10241 24667
rect 9456 24636 10241 24664
rect 9398 24624 9404 24627
rect 9456 24624 9462 24636
rect 10229 24633 10241 24636
rect 10275 24633 10287 24667
rect 10229 24627 10287 24633
rect 8478 24596 8484 24608
rect 5132 24568 6316 24596
rect 8439 24568 8484 24596
rect 5132 24556 5138 24568
rect 8478 24556 8484 24568
rect 8536 24556 8542 24608
rect 10612 24596 10640 24695
rect 10965 24667 11023 24673
rect 10965 24633 10977 24667
rect 11011 24633 11023 24667
rect 10965 24627 11023 24633
rect 10980 24596 11008 24627
rect 10612 24568 11008 24596
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 7193 24395 7251 24401
rect 7193 24392 7205 24395
rect 4126 24364 7205 24392
rect 2774 24216 2780 24268
rect 2832 24256 2838 24268
rect 2961 24259 3019 24265
rect 2961 24256 2973 24259
rect 2832 24228 2973 24256
rect 2832 24216 2838 24228
rect 2961 24225 2973 24228
rect 3007 24256 3019 24259
rect 4126 24256 4154 24364
rect 7193 24361 7205 24364
rect 7239 24361 7251 24395
rect 7193 24355 7251 24361
rect 7282 24352 7288 24404
rect 7340 24392 7346 24404
rect 7837 24395 7895 24401
rect 7837 24392 7849 24395
rect 7340 24364 7849 24392
rect 7340 24352 7346 24364
rect 7837 24361 7849 24364
rect 7883 24392 7895 24395
rect 8018 24392 8024 24404
rect 7883 24364 8024 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 8018 24352 8024 24364
rect 8076 24352 8082 24404
rect 9766 24392 9772 24404
rect 9727 24364 9772 24392
rect 9766 24352 9772 24364
rect 9824 24352 9830 24404
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10008 24364 11376 24392
rect 10008 24352 10014 24364
rect 5261 24327 5319 24333
rect 5261 24293 5273 24327
rect 5307 24324 5319 24327
rect 5350 24324 5356 24336
rect 5307 24296 5356 24324
rect 5307 24293 5319 24296
rect 5261 24287 5319 24293
rect 5350 24284 5356 24296
rect 5408 24324 5414 24336
rect 6641 24327 6699 24333
rect 6641 24324 6653 24327
rect 5408 24296 6653 24324
rect 5408 24284 5414 24296
rect 6641 24293 6653 24296
rect 6687 24324 6699 24327
rect 7098 24324 7104 24336
rect 6687 24296 7104 24324
rect 6687 24293 6699 24296
rect 6641 24287 6699 24293
rect 4246 24256 4252 24268
rect 3007 24228 4154 24256
rect 4207 24228 4252 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 4246 24216 4252 24228
rect 4304 24216 4310 24268
rect 5718 24256 5724 24268
rect 5679 24228 5724 24256
rect 5718 24216 5724 24228
rect 5776 24256 5782 24268
rect 6748 24265 6776 24296
rect 7098 24284 7104 24296
rect 7156 24284 7162 24336
rect 8478 24284 8484 24336
rect 8536 24324 8542 24336
rect 11241 24327 11299 24333
rect 11241 24324 11253 24327
rect 8536 24296 11253 24324
rect 8536 24284 8542 24296
rect 11241 24293 11253 24296
rect 11287 24293 11299 24327
rect 11241 24287 11299 24293
rect 6181 24259 6239 24265
rect 6181 24256 6193 24259
rect 5776 24228 6193 24256
rect 5776 24216 5782 24228
rect 6181 24225 6193 24228
rect 6227 24225 6239 24259
rect 6733 24259 6791 24265
rect 6733 24256 6745 24259
rect 6711 24228 6745 24256
rect 6181 24219 6239 24225
rect 6733 24225 6745 24228
rect 6779 24225 6791 24259
rect 7006 24256 7012 24268
rect 6967 24228 7012 24256
rect 6733 24219 6791 24225
rect 7006 24216 7012 24228
rect 7064 24216 7070 24268
rect 8297 24259 8355 24265
rect 8297 24225 8309 24259
rect 8343 24225 8355 24259
rect 8297 24219 8355 24225
rect 8757 24259 8815 24265
rect 8757 24225 8769 24259
rect 8803 24256 8815 24259
rect 9306 24256 9312 24268
rect 8803 24228 9312 24256
rect 8803 24225 8815 24228
rect 8757 24219 8815 24225
rect 3970 24148 3976 24200
rect 4028 24188 4034 24200
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 4028 24160 4169 24188
rect 4028 24148 4034 24160
rect 4157 24157 4169 24160
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 4338 24148 4344 24200
rect 4396 24188 4402 24200
rect 8312 24188 8340 24219
rect 9306 24216 9312 24228
rect 9364 24216 9370 24268
rect 9674 24256 9680 24268
rect 9635 24228 9680 24256
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10134 24256 10140 24268
rect 10095 24228 10140 24256
rect 10134 24216 10140 24228
rect 10192 24216 10198 24268
rect 11348 24265 11376 24364
rect 11333 24259 11391 24265
rect 11333 24225 11345 24259
rect 11379 24256 11391 24259
rect 11514 24256 11520 24268
rect 11379 24228 11520 24256
rect 11379 24225 11391 24228
rect 11333 24219 11391 24225
rect 11514 24216 11520 24228
rect 11572 24256 11578 24268
rect 12529 24259 12587 24265
rect 12529 24256 12541 24259
rect 11572 24228 12541 24256
rect 11572 24216 11578 24228
rect 12529 24225 12541 24228
rect 12575 24225 12587 24259
rect 12529 24219 12587 24225
rect 8846 24188 8852 24200
rect 4396 24160 8852 24188
rect 4396 24148 4402 24160
rect 8846 24148 8852 24160
rect 8904 24148 8910 24200
rect 8938 24148 8944 24200
rect 8996 24188 9002 24200
rect 12434 24188 12440 24200
rect 8996 24160 12440 24188
rect 8996 24148 9002 24160
rect 12434 24148 12440 24160
rect 12492 24148 12498 24200
rect 3326 24080 3332 24132
rect 3384 24120 3390 24132
rect 3513 24123 3571 24129
rect 3513 24120 3525 24123
rect 3384 24092 3525 24120
rect 3384 24080 3390 24092
rect 3513 24089 3525 24092
rect 3559 24120 3571 24123
rect 4430 24120 4436 24132
rect 3559 24092 4436 24120
rect 3559 24089 3571 24092
rect 3513 24083 3571 24089
rect 4430 24080 4436 24092
rect 4488 24080 4494 24132
rect 4614 24080 4620 24132
rect 4672 24120 4678 24132
rect 5629 24123 5687 24129
rect 5629 24120 5641 24123
rect 4672 24092 5641 24120
rect 4672 24080 4678 24092
rect 5629 24089 5641 24092
rect 5675 24120 5687 24123
rect 5810 24120 5816 24132
rect 5675 24092 5816 24120
rect 5675 24089 5687 24092
rect 5629 24083 5687 24089
rect 5810 24080 5816 24092
rect 5868 24120 5874 24132
rect 6178 24120 6184 24132
rect 5868 24092 6184 24120
rect 5868 24080 5874 24092
rect 6178 24080 6184 24092
rect 6236 24080 6242 24132
rect 6638 24080 6644 24132
rect 6696 24120 6702 24132
rect 6825 24123 6883 24129
rect 6825 24120 6837 24123
rect 6696 24092 6837 24120
rect 6696 24080 6702 24092
rect 6825 24089 6837 24092
rect 6871 24120 6883 24123
rect 7374 24120 7380 24132
rect 6871 24092 7380 24120
rect 6871 24089 6883 24092
rect 6825 24083 6883 24089
rect 7374 24080 7380 24092
rect 7432 24080 7438 24132
rect 8481 24123 8539 24129
rect 8481 24089 8493 24123
rect 8527 24120 8539 24123
rect 8570 24120 8576 24132
rect 8527 24092 8576 24120
rect 8527 24089 8539 24092
rect 8481 24083 8539 24089
rect 8570 24080 8576 24092
rect 8628 24120 8634 24132
rect 10134 24120 10140 24132
rect 8628 24092 10140 24120
rect 8628 24080 8634 24092
rect 10134 24080 10140 24092
rect 10192 24080 10198 24132
rect 3142 24052 3148 24064
rect 3103 24024 3148 24052
rect 3142 24012 3148 24024
rect 3200 24012 3206 24064
rect 4154 24012 4160 24064
rect 4212 24052 4218 24064
rect 4338 24052 4344 24064
rect 4212 24024 4344 24052
rect 4212 24012 4218 24024
rect 4338 24012 4344 24024
rect 4396 24012 4402 24064
rect 5905 24055 5963 24061
rect 5905 24021 5917 24055
rect 5951 24052 5963 24055
rect 5994 24052 6000 24064
rect 5951 24024 6000 24052
rect 5951 24021 5963 24024
rect 5905 24015 5963 24021
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 8754 24012 8760 24064
rect 8812 24052 8818 24064
rect 9125 24055 9183 24061
rect 9125 24052 9137 24055
rect 8812 24024 9137 24052
rect 8812 24012 8818 24024
rect 9125 24021 9137 24024
rect 9171 24021 9183 24055
rect 10686 24052 10692 24064
rect 10647 24024 10692 24052
rect 9125 24015 9183 24021
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 11149 24055 11207 24061
rect 11149 24021 11161 24055
rect 11195 24052 11207 24055
rect 11422 24052 11428 24064
rect 11195 24024 11428 24052
rect 11195 24021 11207 24024
rect 11149 24015 11207 24021
rect 11422 24012 11428 24024
rect 11480 24012 11486 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 2774 23848 2780 23860
rect 2735 23820 2780 23848
rect 2774 23808 2780 23820
rect 2832 23808 2838 23860
rect 4341 23851 4399 23857
rect 4341 23817 4353 23851
rect 4387 23848 4399 23851
rect 4614 23848 4620 23860
rect 4387 23820 4620 23848
rect 4387 23817 4399 23820
rect 4341 23811 4399 23817
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 6638 23848 6644 23860
rect 4764 23820 4809 23848
rect 6599 23820 6644 23848
rect 4764 23808 4770 23820
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 7098 23808 7104 23860
rect 7156 23848 7162 23860
rect 7561 23851 7619 23857
rect 7561 23848 7573 23851
rect 7156 23820 7573 23848
rect 7156 23808 7162 23820
rect 7561 23817 7573 23820
rect 7607 23817 7619 23851
rect 8202 23848 8208 23860
rect 8163 23820 8208 23848
rect 7561 23811 7619 23817
rect 8202 23808 8208 23820
rect 8260 23848 8266 23860
rect 8941 23851 8999 23857
rect 8941 23848 8953 23851
rect 8260 23820 8953 23848
rect 8260 23808 8266 23820
rect 8941 23817 8953 23820
rect 8987 23848 8999 23851
rect 9950 23848 9956 23860
rect 8987 23820 9956 23848
rect 8987 23817 8999 23820
rect 8941 23811 8999 23817
rect 9950 23808 9956 23820
rect 10008 23808 10014 23860
rect 10134 23848 10140 23860
rect 10095 23820 10140 23848
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 11514 23848 11520 23860
rect 11475 23820 11520 23848
rect 11514 23808 11520 23820
rect 11572 23848 11578 23860
rect 12713 23851 12771 23857
rect 12713 23848 12725 23851
rect 11572 23820 12725 23848
rect 11572 23808 11578 23820
rect 12713 23817 12725 23820
rect 12759 23817 12771 23851
rect 12713 23811 12771 23817
rect 3326 23780 3332 23792
rect 3287 23752 3332 23780
rect 3326 23740 3332 23752
rect 3384 23740 3390 23792
rect 6914 23740 6920 23792
rect 6972 23780 6978 23792
rect 7239 23783 7297 23789
rect 7239 23780 7251 23783
rect 6972 23752 7251 23780
rect 6972 23740 6978 23752
rect 7239 23749 7251 23752
rect 7285 23749 7297 23783
rect 7239 23743 7297 23749
rect 7374 23740 7380 23792
rect 7432 23780 7438 23792
rect 8220 23780 8248 23808
rect 7432 23752 8248 23780
rect 7432 23740 7438 23752
rect 8294 23740 8300 23792
rect 8352 23780 8358 23792
rect 8573 23783 8631 23789
rect 8573 23780 8585 23783
rect 8352 23752 8585 23780
rect 8352 23740 8358 23752
rect 8573 23749 8585 23752
rect 8619 23780 8631 23783
rect 8803 23783 8861 23789
rect 8803 23780 8815 23783
rect 8619 23752 8815 23780
rect 8619 23749 8631 23752
rect 8573 23743 8631 23749
rect 8803 23749 8815 23752
rect 8849 23749 8861 23783
rect 9306 23780 9312 23792
rect 8803 23743 8861 23749
rect 9048 23752 9312 23780
rect 3973 23715 4031 23721
rect 3973 23681 3985 23715
rect 4019 23712 4031 23715
rect 5718 23712 5724 23724
rect 4019 23684 5724 23712
rect 4019 23681 4031 23684
rect 3973 23675 4031 23681
rect 5718 23672 5724 23684
rect 5776 23672 5782 23724
rect 6273 23715 6331 23721
rect 6273 23681 6285 23715
rect 6319 23712 6331 23715
rect 7006 23712 7012 23724
rect 6319 23684 7012 23712
rect 6319 23681 6331 23684
rect 6273 23675 6331 23681
rect 7006 23672 7012 23684
rect 7064 23712 7070 23724
rect 7466 23712 7472 23724
rect 7064 23684 7472 23712
rect 7064 23672 7070 23684
rect 7466 23672 7472 23684
rect 7524 23712 7530 23724
rect 9048 23721 9076 23752
rect 9306 23740 9312 23752
rect 9364 23780 9370 23792
rect 9364 23752 11928 23780
rect 9364 23740 9370 23752
rect 9033 23715 9091 23721
rect 9033 23712 9045 23715
rect 7524 23684 9045 23712
rect 7524 23672 7530 23684
rect 9033 23681 9045 23684
rect 9079 23681 9091 23715
rect 9033 23675 9091 23681
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23712 10563 23715
rect 11422 23712 11428 23724
rect 10551 23684 11428 23712
rect 10551 23681 10563 23684
rect 10505 23675 10563 23681
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11900 23721 11928 23752
rect 12066 23740 12072 23792
rect 12124 23780 12130 23792
rect 12253 23783 12311 23789
rect 12253 23780 12265 23783
rect 12124 23752 12265 23780
rect 12124 23740 12130 23752
rect 12253 23749 12265 23752
rect 12299 23780 12311 23783
rect 12575 23783 12633 23789
rect 12575 23780 12587 23783
rect 12299 23752 12587 23780
rect 12299 23749 12311 23752
rect 12253 23743 12311 23749
rect 12575 23749 12587 23752
rect 12621 23749 12633 23783
rect 12575 23743 12633 23749
rect 11885 23715 11943 23721
rect 11885 23681 11897 23715
rect 11931 23712 11943 23715
rect 12805 23715 12863 23721
rect 12805 23712 12817 23715
rect 11931 23684 12817 23712
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 12805 23681 12817 23684
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 3145 23647 3203 23653
rect 3145 23613 3157 23647
rect 3191 23644 3203 23647
rect 3234 23644 3240 23656
rect 3191 23616 3240 23644
rect 3191 23613 3203 23616
rect 3145 23607 3203 23613
rect 3234 23604 3240 23616
rect 3292 23604 3298 23656
rect 3513 23647 3571 23653
rect 3513 23613 3525 23647
rect 3559 23644 3571 23647
rect 4062 23644 4068 23656
rect 3559 23616 4068 23644
rect 3559 23613 3571 23616
rect 3513 23607 3571 23613
rect 4062 23604 4068 23616
rect 4120 23604 4126 23656
rect 4798 23644 4804 23656
rect 4759 23616 4804 23644
rect 4798 23604 4804 23616
rect 4856 23644 4862 23656
rect 5074 23644 5080 23656
rect 4856 23616 5080 23644
rect 4856 23604 4862 23616
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 5629 23647 5687 23653
rect 5629 23644 5641 23647
rect 5321 23616 5641 23644
rect 4706 23536 4712 23588
rect 4764 23576 4770 23588
rect 5321 23576 5349 23616
rect 5629 23613 5641 23616
rect 5675 23613 5687 23647
rect 5810 23644 5816 23656
rect 5771 23616 5816 23644
rect 5629 23607 5687 23613
rect 5810 23604 5816 23616
rect 5868 23644 5874 23656
rect 5868 23616 7236 23644
rect 5868 23604 5874 23616
rect 4764 23548 5349 23576
rect 4764 23536 4770 23548
rect 5534 23536 5540 23588
rect 5592 23576 5598 23588
rect 5828 23576 5856 23604
rect 5592 23548 5856 23576
rect 7101 23579 7159 23585
rect 5592 23536 5598 23548
rect 7101 23545 7113 23579
rect 7147 23545 7159 23579
rect 7208 23576 7236 23616
rect 7558 23604 7564 23656
rect 7616 23644 7622 23656
rect 9401 23647 9459 23653
rect 9401 23644 9413 23647
rect 7616 23616 9413 23644
rect 7616 23604 7622 23616
rect 9401 23613 9413 23616
rect 9447 23613 9459 23647
rect 9401 23607 9459 23613
rect 8665 23579 8723 23585
rect 8665 23576 8677 23579
rect 7208 23548 8677 23576
rect 7101 23539 7159 23545
rect 8665 23545 8677 23548
rect 8711 23576 8723 23579
rect 8754 23576 8760 23588
rect 8711 23548 8760 23576
rect 8711 23545 8723 23548
rect 8665 23539 8723 23545
rect 4890 23508 4896 23520
rect 4851 23480 4896 23508
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 5166 23468 5172 23520
rect 5224 23508 5230 23520
rect 7116 23508 7144 23539
rect 8754 23536 8760 23548
rect 8812 23536 8818 23588
rect 10597 23579 10655 23585
rect 10597 23545 10609 23579
rect 10643 23576 10655 23579
rect 10686 23576 10692 23588
rect 10643 23548 10692 23576
rect 10643 23545 10655 23548
rect 10597 23539 10655 23545
rect 10686 23536 10692 23548
rect 10744 23536 10750 23588
rect 11149 23579 11207 23585
rect 11149 23545 11161 23579
rect 11195 23576 11207 23579
rect 11514 23576 11520 23588
rect 11195 23548 11520 23576
rect 11195 23545 11207 23548
rect 11149 23539 11207 23545
rect 11514 23536 11520 23548
rect 11572 23536 11578 23588
rect 12434 23576 12440 23588
rect 12395 23548 12440 23576
rect 12434 23536 12440 23548
rect 12492 23536 12498 23588
rect 7282 23508 7288 23520
rect 5224 23480 7288 23508
rect 5224 23468 5230 23480
rect 7282 23468 7288 23480
rect 7340 23468 7346 23520
rect 9306 23468 9312 23520
rect 9364 23508 9370 23520
rect 9674 23508 9680 23520
rect 9364 23480 9680 23508
rect 9364 23468 9370 23480
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 12250 23468 12256 23520
rect 12308 23508 12314 23520
rect 13081 23511 13139 23517
rect 13081 23508 13093 23511
rect 12308 23480 13093 23508
rect 12308 23468 12314 23480
rect 13081 23477 13093 23480
rect 13127 23477 13139 23511
rect 13081 23471 13139 23477
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 3881 23307 3939 23313
rect 3881 23273 3893 23307
rect 3927 23304 3939 23307
rect 4246 23304 4252 23316
rect 3927 23276 4252 23304
rect 3927 23273 3939 23276
rect 3881 23267 3939 23273
rect 4246 23264 4252 23276
rect 4304 23264 4310 23316
rect 4982 23264 4988 23316
rect 5040 23304 5046 23316
rect 5353 23307 5411 23313
rect 5353 23304 5365 23307
rect 5040 23276 5365 23304
rect 5040 23264 5046 23276
rect 5353 23273 5365 23276
rect 5399 23273 5411 23307
rect 5353 23267 5411 23273
rect 5442 23264 5448 23316
rect 5500 23304 5506 23316
rect 5718 23304 5724 23316
rect 5500 23276 5724 23304
rect 5500 23264 5506 23276
rect 5718 23264 5724 23276
rect 5776 23264 5782 23316
rect 6638 23264 6644 23316
rect 6696 23304 6702 23316
rect 6733 23307 6791 23313
rect 6733 23304 6745 23307
rect 6696 23276 6745 23304
rect 6696 23264 6702 23276
rect 6733 23273 6745 23276
rect 6779 23273 6791 23307
rect 7466 23304 7472 23316
rect 7427 23276 7472 23304
rect 6733 23267 6791 23273
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 8846 23264 8852 23316
rect 8904 23304 8910 23316
rect 9033 23307 9091 23313
rect 9033 23304 9045 23307
rect 8904 23276 9045 23304
rect 8904 23264 8910 23276
rect 9033 23273 9045 23276
rect 9079 23273 9091 23307
rect 12066 23304 12072 23316
rect 9033 23267 9091 23273
rect 9140 23276 12072 23304
rect 2222 23196 2228 23248
rect 2280 23236 2286 23248
rect 2593 23239 2651 23245
rect 2593 23236 2605 23239
rect 2280 23208 2605 23236
rect 2280 23196 2286 23208
rect 2593 23205 2605 23208
rect 2639 23236 2651 23239
rect 3142 23236 3148 23248
rect 2639 23208 3148 23236
rect 2639 23205 2651 23208
rect 2593 23199 2651 23205
rect 3142 23196 3148 23208
rect 3200 23196 3206 23248
rect 3513 23239 3571 23245
rect 3513 23205 3525 23239
rect 3559 23236 3571 23239
rect 3970 23236 3976 23248
rect 3559 23208 3976 23236
rect 3559 23205 3571 23208
rect 3513 23199 3571 23205
rect 3970 23196 3976 23208
rect 4028 23196 4034 23248
rect 6914 23196 6920 23248
rect 6972 23236 6978 23248
rect 7193 23239 7251 23245
rect 7193 23236 7205 23239
rect 6972 23208 7205 23236
rect 6972 23196 6978 23208
rect 7193 23205 7205 23208
rect 7239 23236 7251 23239
rect 8294 23236 8300 23248
rect 7239 23208 8300 23236
rect 7239 23205 7251 23208
rect 7193 23199 7251 23205
rect 8294 23196 8300 23208
rect 8352 23236 8358 23248
rect 9140 23236 9168 23276
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 12713 23307 12771 23313
rect 12713 23304 12725 23307
rect 12492 23276 12725 23304
rect 12492 23264 12498 23276
rect 12713 23273 12725 23276
rect 12759 23273 12771 23307
rect 12713 23267 12771 23273
rect 8352 23208 9168 23236
rect 8352 23196 8358 23208
rect 10410 23196 10416 23248
rect 10468 23236 10474 23248
rect 10505 23239 10563 23245
rect 10505 23236 10517 23239
rect 10468 23208 10517 23236
rect 10468 23196 10474 23208
rect 10505 23205 10517 23208
rect 10551 23236 10563 23239
rect 10686 23236 10692 23248
rect 10551 23208 10692 23236
rect 10551 23205 10563 23208
rect 10505 23199 10563 23205
rect 10686 23196 10692 23208
rect 10744 23196 10750 23248
rect 2682 23128 2688 23180
rect 2740 23168 2746 23180
rect 2777 23171 2835 23177
rect 2777 23168 2789 23171
rect 2740 23140 2789 23168
rect 2740 23128 2746 23140
rect 2777 23137 2789 23140
rect 2823 23168 2835 23171
rect 4116 23171 4174 23177
rect 2823 23140 3832 23168
rect 2823 23137 2835 23140
rect 2777 23131 2835 23137
rect 3145 23103 3203 23109
rect 3145 23069 3157 23103
rect 3191 23100 3203 23103
rect 3510 23100 3516 23112
rect 3191 23072 3516 23100
rect 3191 23069 3203 23072
rect 3145 23063 3203 23069
rect 3510 23060 3516 23072
rect 3568 23060 3574 23112
rect 3804 23100 3832 23140
rect 4116 23137 4128 23171
rect 4162 23168 4174 23171
rect 4522 23168 4528 23180
rect 4162 23140 4528 23168
rect 4162 23137 4174 23140
rect 4116 23131 4174 23137
rect 4522 23128 4528 23140
rect 4580 23128 4586 23180
rect 4893 23171 4951 23177
rect 4893 23137 4905 23171
rect 4939 23168 4951 23171
rect 5074 23168 5080 23180
rect 4939 23140 5080 23168
rect 4939 23137 4951 23140
rect 4893 23131 4951 23137
rect 5074 23128 5080 23140
rect 5132 23168 5138 23180
rect 5442 23168 5448 23180
rect 5132 23140 5448 23168
rect 5132 23128 5138 23140
rect 5442 23128 5448 23140
rect 5500 23128 5506 23180
rect 5534 23128 5540 23180
rect 5592 23168 5598 23180
rect 5721 23171 5779 23177
rect 5721 23168 5733 23171
rect 5592 23140 5733 23168
rect 5592 23128 5598 23140
rect 5721 23137 5733 23140
rect 5767 23137 5779 23171
rect 6086 23168 6092 23180
rect 6047 23140 6092 23168
rect 5721 23131 5779 23137
rect 6086 23128 6092 23140
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23168 7898 23180
rect 8021 23171 8079 23177
rect 8021 23168 8033 23171
rect 7892 23140 8033 23168
rect 7892 23128 7898 23140
rect 8021 23137 8033 23140
rect 8067 23137 8079 23171
rect 8478 23168 8484 23180
rect 8439 23140 8484 23168
rect 8021 23131 8079 23137
rect 8478 23128 8484 23140
rect 8536 23128 8542 23180
rect 11882 23168 11888 23180
rect 11440 23140 11888 23168
rect 5166 23100 5172 23112
rect 3804 23072 5172 23100
rect 5166 23060 5172 23072
rect 5224 23060 5230 23112
rect 5994 23060 6000 23112
rect 6052 23100 6058 23112
rect 8754 23100 8760 23112
rect 6052 23072 8432 23100
rect 8715 23072 8760 23100
rect 6052 23060 6058 23072
rect 4203 23035 4261 23041
rect 4203 23001 4215 23035
rect 4249 23032 4261 23035
rect 5626 23032 5632 23044
rect 4249 23004 5632 23032
rect 4249 23001 4261 23004
rect 4203 22995 4261 23001
rect 5626 22992 5632 23004
rect 5684 22992 5690 23044
rect 8404 22964 8432 23072
rect 8754 23060 8760 23072
rect 8812 23060 8818 23112
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23100 10287 23103
rect 10413 23103 10471 23109
rect 10413 23100 10425 23103
rect 10275 23072 10425 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 10413 23069 10425 23072
rect 10459 23100 10471 23103
rect 11330 23100 11336 23112
rect 10459 23072 11336 23100
rect 10459 23069 10471 23072
rect 10413 23063 10471 23069
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 10965 23035 11023 23041
rect 10965 23001 10977 23035
rect 11011 23032 11023 23035
rect 11146 23032 11152 23044
rect 11011 23004 11152 23032
rect 11011 23001 11023 23004
rect 10965 22995 11023 23001
rect 11146 22992 11152 23004
rect 11204 22992 11210 23044
rect 11440 22964 11468 23140
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 11974 23128 11980 23180
rect 12032 23168 12038 23180
rect 12069 23171 12127 23177
rect 12069 23168 12081 23171
rect 12032 23140 12081 23168
rect 12032 23128 12038 23140
rect 12069 23137 12081 23140
rect 12115 23168 12127 23171
rect 12710 23168 12716 23180
rect 12115 23140 12716 23168
rect 12115 23137 12127 23140
rect 12069 23131 12127 23137
rect 12710 23128 12716 23140
rect 12768 23128 12774 23180
rect 8404 22936 11468 22964
rect 12066 22924 12072 22976
rect 12124 22964 12130 22976
rect 12161 22967 12219 22973
rect 12161 22964 12173 22967
rect 12124 22936 12173 22964
rect 12124 22924 12130 22936
rect 12161 22933 12173 22936
rect 12207 22933 12219 22967
rect 12161 22927 12219 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2222 22760 2228 22772
rect 2183 22732 2228 22760
rect 2222 22720 2228 22732
rect 2280 22720 2286 22772
rect 4341 22763 4399 22769
rect 4341 22729 4353 22763
rect 4387 22760 4399 22763
rect 4522 22760 4528 22772
rect 4387 22732 4528 22760
rect 4387 22729 4399 22732
rect 4341 22723 4399 22729
rect 4522 22720 4528 22732
rect 4580 22720 4586 22772
rect 4798 22760 4804 22772
rect 4759 22732 4804 22760
rect 4798 22720 4804 22732
rect 4856 22720 4862 22772
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 6457 22763 6515 22769
rect 6457 22760 6469 22763
rect 5592 22732 6469 22760
rect 5592 22720 5598 22732
rect 6457 22729 6469 22732
rect 6503 22729 6515 22763
rect 6457 22723 6515 22729
rect 7282 22720 7288 22772
rect 7340 22760 7346 22772
rect 7834 22760 7840 22772
rect 7340 22732 7840 22760
rect 7340 22720 7346 22732
rect 7834 22720 7840 22732
rect 7892 22760 7898 22772
rect 8021 22763 8079 22769
rect 8021 22760 8033 22763
rect 7892 22732 8033 22760
rect 7892 22720 7898 22732
rect 8021 22729 8033 22732
rect 8067 22729 8079 22763
rect 8021 22723 8079 22729
rect 8941 22763 8999 22769
rect 8941 22729 8953 22763
rect 8987 22760 8999 22763
rect 9398 22760 9404 22772
rect 8987 22732 9404 22760
rect 8987 22729 8999 22732
rect 8941 22723 8999 22729
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 11974 22760 11980 22772
rect 11935 22732 11980 22760
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 12802 22720 12808 22772
rect 12860 22760 12866 22772
rect 12897 22763 12955 22769
rect 12897 22760 12909 22763
rect 12860 22732 12909 22760
rect 12860 22720 12866 22732
rect 12897 22729 12909 22732
rect 12943 22729 12955 22763
rect 12897 22723 12955 22729
rect 4154 22652 4160 22704
rect 4212 22692 4218 22704
rect 4430 22692 4436 22704
rect 4212 22664 4436 22692
rect 4212 22652 4218 22664
rect 4430 22652 4436 22664
rect 4488 22652 4494 22704
rect 5442 22652 5448 22704
rect 5500 22692 5506 22704
rect 6089 22695 6147 22701
rect 6089 22692 6101 22695
rect 5500 22664 6101 22692
rect 5500 22652 5506 22664
rect 6089 22661 6101 22664
rect 6135 22661 6147 22695
rect 6089 22655 6147 22661
rect 9953 22695 10011 22701
rect 9953 22661 9965 22695
rect 9999 22692 10011 22695
rect 10962 22692 10968 22704
rect 9999 22664 10968 22692
rect 9999 22661 10011 22664
rect 9953 22655 10011 22661
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 11422 22652 11428 22704
rect 11480 22692 11486 22704
rect 12575 22695 12633 22701
rect 12575 22692 12587 22695
rect 11480 22664 12587 22692
rect 11480 22652 11486 22664
rect 12575 22661 12587 22664
rect 12621 22661 12633 22695
rect 12575 22655 12633 22661
rect 4890 22624 4896 22636
rect 4851 22596 4896 22624
rect 4890 22584 4896 22596
rect 4948 22584 4954 22636
rect 7193 22627 7251 22633
rect 7193 22624 7205 22627
rect 5000 22596 7205 22624
rect 2317 22559 2375 22565
rect 2317 22525 2329 22559
rect 2363 22556 2375 22559
rect 2866 22556 2872 22568
rect 2363 22528 2872 22556
rect 2363 22525 2375 22528
rect 2317 22519 2375 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22556 4123 22559
rect 4154 22556 4160 22568
rect 4111 22528 4160 22556
rect 4111 22525 4123 22528
rect 4065 22519 4123 22525
rect 4154 22516 4160 22528
rect 4212 22556 4218 22568
rect 5000 22556 5028 22596
rect 7193 22593 7205 22596
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 9033 22627 9091 22633
rect 9033 22624 9045 22627
rect 8812 22596 9045 22624
rect 8812 22584 8818 22596
rect 9033 22593 9045 22596
rect 9079 22593 9091 22627
rect 11146 22624 11152 22636
rect 11107 22596 11152 22624
rect 9033 22587 9091 22593
rect 11146 22584 11152 22596
rect 11204 22584 11210 22636
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 13587 22627 13645 22633
rect 13587 22624 13599 22627
rect 11388 22596 13599 22624
rect 11388 22584 11394 22596
rect 13587 22593 13599 22596
rect 13633 22593 13645 22627
rect 13587 22587 13645 22593
rect 4212 22528 5028 22556
rect 12345 22559 12403 22565
rect 4212 22516 4218 22528
rect 12345 22525 12357 22559
rect 12391 22525 12403 22559
rect 12345 22519 12403 22525
rect 3418 22488 3424 22500
rect 3379 22460 3424 22488
rect 3418 22448 3424 22460
rect 3476 22448 3482 22500
rect 3513 22491 3571 22497
rect 3513 22457 3525 22491
rect 3559 22488 3571 22491
rect 3878 22488 3884 22500
rect 3559 22460 3884 22488
rect 3559 22457 3571 22460
rect 3513 22451 3571 22457
rect 2498 22420 2504 22432
rect 2459 22392 2504 22420
rect 2498 22380 2504 22392
rect 2556 22380 2562 22432
rect 2866 22420 2872 22432
rect 2827 22392 2872 22420
rect 2866 22380 2872 22392
rect 2924 22380 2930 22432
rect 3237 22423 3295 22429
rect 3237 22389 3249 22423
rect 3283 22420 3295 22423
rect 3528 22420 3556 22451
rect 3878 22448 3884 22460
rect 3936 22448 3942 22500
rect 4246 22448 4252 22500
rect 4304 22488 4310 22500
rect 4304 22460 4752 22488
rect 4304 22448 4310 22460
rect 3283 22392 3556 22420
rect 4724 22420 4752 22460
rect 4798 22448 4804 22500
rect 4856 22488 4862 22500
rect 5214 22491 5272 22497
rect 5214 22488 5226 22491
rect 4856 22460 5226 22488
rect 4856 22448 4862 22460
rect 5214 22457 5226 22460
rect 5260 22488 5272 22491
rect 5350 22488 5356 22500
rect 5260 22460 5356 22488
rect 5260 22457 5272 22460
rect 5214 22451 5272 22457
rect 5350 22448 5356 22460
rect 5408 22448 5414 22500
rect 6730 22448 6736 22500
rect 6788 22488 6794 22500
rect 6917 22491 6975 22497
rect 6917 22488 6929 22491
rect 6788 22460 6929 22488
rect 6788 22448 6794 22460
rect 6917 22457 6929 22460
rect 6963 22457 6975 22491
rect 6917 22451 6975 22457
rect 7009 22491 7067 22497
rect 7009 22457 7021 22491
rect 7055 22457 7067 22491
rect 7009 22451 7067 22457
rect 10873 22491 10931 22497
rect 10873 22457 10885 22491
rect 10919 22457 10931 22491
rect 10873 22451 10931 22457
rect 5813 22423 5871 22429
rect 5813 22420 5825 22423
rect 4724 22392 5825 22420
rect 3283 22389 3295 22392
rect 3237 22383 3295 22389
rect 5813 22389 5825 22392
rect 5859 22420 5871 22423
rect 6638 22420 6644 22432
rect 5859 22392 6644 22420
rect 5859 22389 5871 22392
rect 5813 22383 5871 22389
rect 6638 22380 6644 22392
rect 6696 22420 6702 22432
rect 7024 22420 7052 22451
rect 8478 22420 8484 22432
rect 6696 22392 7052 22420
rect 8439 22392 8484 22420
rect 6696 22380 6702 22392
rect 8478 22380 8484 22392
rect 8536 22380 8542 22432
rect 9398 22420 9404 22432
rect 9359 22392 9404 22420
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 10318 22420 10324 22432
rect 10279 22392 10324 22420
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 10888 22420 10916 22451
rect 10962 22448 10968 22500
rect 11020 22488 11026 22500
rect 11020 22460 11065 22488
rect 11020 22448 11026 22460
rect 12250 22448 12256 22500
rect 12308 22488 12314 22500
rect 12360 22488 12388 22519
rect 12894 22516 12900 22568
rect 12952 22556 12958 22568
rect 13484 22559 13542 22565
rect 13484 22556 13496 22559
rect 12952 22528 13496 22556
rect 12952 22516 12958 22528
rect 13484 22525 13496 22528
rect 13530 22556 13542 22559
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 13530 22528 13921 22556
rect 13530 22525 13542 22528
rect 13484 22519 13542 22525
rect 13909 22525 13921 22528
rect 13955 22525 13967 22559
rect 13909 22519 13967 22525
rect 12802 22488 12808 22500
rect 12308 22460 12808 22488
rect 12308 22448 12314 22460
rect 12802 22448 12808 22460
rect 12860 22448 12866 22500
rect 11330 22420 11336 22432
rect 10888 22392 11336 22420
rect 11330 22380 11336 22392
rect 11388 22380 11394 22432
rect 11422 22380 11428 22432
rect 11480 22420 11486 22432
rect 12066 22420 12072 22432
rect 11480 22392 12072 22420
rect 11480 22380 11486 22392
rect 12066 22380 12072 22392
rect 12124 22380 12130 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 2682 22216 2688 22228
rect 2643 22188 2688 22216
rect 2682 22176 2688 22188
rect 2740 22176 2746 22228
rect 3099 22219 3157 22225
rect 3099 22185 3111 22219
rect 3145 22216 3157 22219
rect 3418 22216 3424 22228
rect 3145 22188 3424 22216
rect 3145 22185 3157 22188
rect 3099 22179 3157 22185
rect 3418 22176 3424 22188
rect 3476 22176 3482 22228
rect 4525 22219 4583 22225
rect 4525 22185 4537 22219
rect 4571 22216 4583 22219
rect 4890 22216 4896 22228
rect 4571 22188 4896 22216
rect 4571 22185 4583 22188
rect 4525 22179 4583 22185
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 5350 22216 5356 22228
rect 5311 22188 5356 22216
rect 5350 22176 5356 22188
rect 5408 22176 5414 22228
rect 5626 22176 5632 22228
rect 5684 22216 5690 22228
rect 6273 22219 6331 22225
rect 6273 22216 6285 22219
rect 5684 22188 6285 22216
rect 5684 22176 5690 22188
rect 6273 22185 6285 22188
rect 6319 22216 6331 22219
rect 6730 22216 6736 22228
rect 6319 22188 6736 22216
rect 6319 22185 6331 22188
rect 6273 22179 6331 22185
rect 6730 22176 6736 22188
rect 6788 22176 6794 22228
rect 7006 22216 7012 22228
rect 6967 22188 7012 22216
rect 7006 22176 7012 22188
rect 7064 22176 7070 22228
rect 8754 22176 8760 22228
rect 8812 22216 8818 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8812 22188 9045 22216
rect 8812 22176 8818 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 10962 22216 10968 22228
rect 10875 22188 10968 22216
rect 9033 22179 9091 22185
rect 10962 22176 10968 22188
rect 11020 22216 11026 22228
rect 11020 22188 13216 22216
rect 11020 22176 11026 22188
rect 4801 22151 4859 22157
rect 4801 22117 4813 22151
rect 4847 22148 4859 22151
rect 6086 22148 6092 22160
rect 4847 22120 6092 22148
rect 4847 22117 4859 22120
rect 4801 22111 4859 22117
rect 6086 22108 6092 22120
rect 6144 22108 6150 22160
rect 6638 22148 6644 22160
rect 6599 22120 6644 22148
rect 6638 22108 6644 22120
rect 6696 22108 6702 22160
rect 8199 22151 8257 22157
rect 8199 22117 8211 22151
rect 8245 22148 8257 22151
rect 9398 22148 9404 22160
rect 8245 22120 9404 22148
rect 8245 22117 8257 22120
rect 8199 22111 8257 22117
rect 9398 22108 9404 22120
rect 9456 22148 9462 22160
rect 9998 22151 10056 22157
rect 9998 22148 10010 22151
rect 9456 22120 10010 22148
rect 9456 22108 9462 22120
rect 9998 22117 10010 22120
rect 10044 22117 10056 22151
rect 11606 22148 11612 22160
rect 11567 22120 11612 22148
rect 9998 22111 10056 22117
rect 11606 22108 11612 22120
rect 11664 22108 11670 22160
rect 11974 22108 11980 22160
rect 12032 22148 12038 22160
rect 13188 22157 13216 22188
rect 12437 22151 12495 22157
rect 12437 22148 12449 22151
rect 12032 22120 12449 22148
rect 12032 22108 12038 22120
rect 12437 22117 12449 22120
rect 12483 22117 12495 22151
rect 12437 22111 12495 22117
rect 13173 22151 13231 22157
rect 13173 22117 13185 22151
rect 13219 22148 13231 22151
rect 13446 22148 13452 22160
rect 13219 22120 13452 22148
rect 13219 22117 13231 22120
rect 13173 22111 13231 22117
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 3028 22083 3086 22089
rect 3028 22049 3040 22083
rect 3074 22080 3086 22083
rect 3326 22080 3332 22092
rect 3074 22052 3332 22080
rect 3074 22049 3086 22052
rect 3028 22043 3086 22049
rect 3326 22040 3332 22052
rect 3384 22040 3390 22092
rect 4982 22080 4988 22092
rect 4943 22052 4988 22080
rect 4982 22040 4988 22052
rect 5040 22040 5046 22092
rect 6822 22080 6828 22092
rect 6783 22052 6828 22080
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22080 8815 22083
rect 10318 22080 10324 22092
rect 8803 22052 10324 22080
rect 8803 22049 8815 22052
rect 8757 22043 8815 22049
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7837 22015 7895 22021
rect 7837 22012 7849 22015
rect 7423 21984 7849 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7837 21981 7849 21984
rect 7883 22012 7895 22015
rect 8110 22012 8116 22024
rect 7883 21984 8116 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 9674 22012 9680 22024
rect 9635 21984 9680 22012
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 11517 22015 11575 22021
rect 11517 21981 11529 22015
rect 11563 22012 11575 22015
rect 12158 22012 12164 22024
rect 11563 21984 12164 22012
rect 11563 21981 11575 21984
rect 11517 21975 11575 21981
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 13078 22012 13084 22024
rect 13039 21984 13084 22012
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 21981 13415 22015
rect 13357 21975 13415 21981
rect 2498 21904 2504 21956
rect 2556 21944 2562 21956
rect 7466 21944 7472 21956
rect 2556 21916 7472 21944
rect 2556 21904 2562 21916
rect 7466 21904 7472 21916
rect 7524 21944 7530 21956
rect 7653 21947 7711 21953
rect 7653 21944 7665 21947
rect 7524 21916 7665 21944
rect 7524 21904 7530 21916
rect 7653 21913 7665 21916
rect 7699 21913 7711 21947
rect 12066 21944 12072 21956
rect 12027 21916 12072 21944
rect 7653 21907 7711 21913
rect 12066 21904 12072 21916
rect 12124 21904 12130 21956
rect 12526 21904 12532 21956
rect 12584 21944 12590 21956
rect 13372 21944 13400 21975
rect 12584 21916 13400 21944
rect 12584 21904 12590 21916
rect 4890 21836 4896 21888
rect 4948 21876 4954 21888
rect 5905 21879 5963 21885
rect 5905 21876 5917 21879
rect 4948 21848 5917 21876
rect 4948 21836 4954 21848
rect 5905 21845 5917 21848
rect 5951 21845 5963 21879
rect 5905 21839 5963 21845
rect 10597 21879 10655 21885
rect 10597 21845 10609 21879
rect 10643 21876 10655 21879
rect 10778 21876 10784 21888
rect 10643 21848 10784 21876
rect 10643 21845 10655 21848
rect 10597 21839 10655 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 11330 21876 11336 21888
rect 11243 21848 11336 21876
rect 11330 21836 11336 21848
rect 11388 21876 11394 21888
rect 11974 21876 11980 21888
rect 11388 21848 11980 21876
rect 11388 21836 11394 21848
rect 11974 21836 11980 21848
rect 12032 21836 12038 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 4157 21675 4215 21681
rect 4157 21641 4169 21675
rect 4203 21672 4215 21675
rect 4982 21672 4988 21684
rect 4203 21644 4988 21672
rect 4203 21641 4215 21644
rect 4157 21635 4215 21641
rect 4982 21632 4988 21644
rect 5040 21632 5046 21684
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5408 21644 5641 21672
rect 5408 21632 5414 21644
rect 5629 21641 5641 21644
rect 5675 21641 5687 21675
rect 5629 21635 5687 21641
rect 7837 21675 7895 21681
rect 7837 21641 7849 21675
rect 7883 21672 7895 21675
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 7883 21644 9137 21672
rect 7883 21641 7895 21644
rect 7837 21635 7895 21641
rect 9125 21641 9137 21644
rect 9171 21672 9183 21675
rect 9398 21672 9404 21684
rect 9171 21644 9404 21672
rect 9171 21641 9183 21644
rect 9125 21635 9183 21641
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 10505 21675 10563 21681
rect 10505 21641 10517 21675
rect 10551 21672 10563 21675
rect 11241 21675 11299 21681
rect 11241 21672 11253 21675
rect 10551 21644 11253 21672
rect 10551 21641 10563 21644
rect 10505 21635 10563 21641
rect 11241 21641 11253 21644
rect 11287 21672 11299 21675
rect 11606 21672 11612 21684
rect 11287 21644 11612 21672
rect 11287 21641 11299 21644
rect 11241 21635 11299 21641
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 12158 21672 12164 21684
rect 12119 21644 12164 21672
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 13446 21672 13452 21684
rect 13407 21644 13452 21672
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 4430 21564 4436 21616
rect 4488 21604 4494 21616
rect 6549 21607 6607 21613
rect 6549 21604 6561 21607
rect 4488 21576 6561 21604
rect 4488 21564 4494 21576
rect 6549 21573 6561 21576
rect 6595 21604 6607 21607
rect 6822 21604 6828 21616
rect 6595 21576 6828 21604
rect 6595 21573 6607 21576
rect 6549 21567 6607 21573
rect 6822 21564 6828 21576
rect 6880 21564 6886 21616
rect 11471 21607 11529 21613
rect 11471 21573 11483 21607
rect 11517 21604 11529 21607
rect 13078 21604 13084 21616
rect 11517 21576 13084 21604
rect 11517 21573 11529 21576
rect 11471 21567 11529 21573
rect 13078 21564 13084 21576
rect 13136 21604 13142 21616
rect 13817 21607 13875 21613
rect 13817 21604 13829 21607
rect 13136 21576 13829 21604
rect 13136 21564 13142 21576
rect 13817 21573 13829 21576
rect 13863 21573 13875 21607
rect 13817 21567 13875 21573
rect 3789 21539 3847 21545
rect 3789 21505 3801 21539
rect 3835 21536 3847 21539
rect 4154 21536 4160 21548
rect 3835 21508 4160 21536
rect 3835 21505 3847 21508
rect 3789 21499 3847 21505
rect 4154 21496 4160 21508
rect 4212 21536 4218 21548
rect 4709 21539 4767 21545
rect 4709 21536 4721 21539
rect 4212 21508 4721 21536
rect 4212 21496 4218 21508
rect 4709 21505 4721 21508
rect 4755 21505 4767 21539
rect 4982 21536 4988 21548
rect 4943 21508 4988 21536
rect 4709 21499 4767 21505
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 6730 21496 6736 21548
rect 6788 21536 6794 21548
rect 7190 21536 7196 21548
rect 6788 21508 7196 21536
rect 6788 21496 6794 21508
rect 7190 21496 7196 21508
rect 7248 21536 7254 21548
rect 7248 21508 7972 21536
rect 7248 21496 7254 21508
rect 7944 21480 7972 21508
rect 12066 21496 12072 21548
rect 12124 21536 12130 21548
rect 12805 21539 12863 21545
rect 12805 21536 12817 21539
rect 12124 21508 12817 21536
rect 12124 21496 12130 21508
rect 12805 21505 12817 21508
rect 12851 21536 12863 21539
rect 13262 21536 13268 21548
rect 12851 21508 13268 21536
rect 12851 21505 12863 21508
rect 12805 21499 12863 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 6984 21471 7042 21477
rect 6984 21437 6996 21471
rect 7030 21468 7042 21471
rect 7374 21468 7380 21480
rect 7030 21440 7380 21468
rect 7030 21437 7042 21440
rect 6984 21431 7042 21437
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 7926 21468 7932 21480
rect 7839 21440 7932 21468
rect 7926 21428 7932 21440
rect 7984 21428 7990 21480
rect 8389 21471 8447 21477
rect 8389 21437 8401 21471
rect 8435 21437 8447 21471
rect 9582 21468 9588 21480
rect 9543 21440 9588 21468
rect 8389 21431 8447 21437
rect 4801 21403 4859 21409
rect 4801 21369 4813 21403
rect 4847 21400 4859 21403
rect 4890 21400 4896 21412
rect 4847 21372 4896 21400
rect 4847 21369 4859 21372
rect 4801 21363 4859 21369
rect 3053 21335 3111 21341
rect 3053 21301 3065 21335
rect 3099 21332 3111 21335
rect 3326 21332 3332 21344
rect 3099 21304 3332 21332
rect 3099 21301 3111 21304
rect 3053 21295 3111 21301
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 4525 21335 4583 21341
rect 4525 21301 4537 21335
rect 4571 21332 4583 21335
rect 4816 21332 4844 21363
rect 4890 21360 4896 21372
rect 4948 21360 4954 21412
rect 7466 21360 7472 21412
rect 7524 21400 7530 21412
rect 8404 21400 8432 21431
rect 9582 21428 9588 21440
rect 9640 21428 9646 21480
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10781 21471 10839 21477
rect 10781 21468 10793 21471
rect 9732 21440 10793 21468
rect 9732 21428 9738 21440
rect 10781 21437 10793 21440
rect 10827 21437 10839 21471
rect 10781 21431 10839 21437
rect 11368 21471 11426 21477
rect 11368 21437 11380 21471
rect 11414 21437 11426 21471
rect 11368 21431 11426 21437
rect 8478 21400 8484 21412
rect 7524 21372 8484 21400
rect 7524 21360 7530 21372
rect 8478 21360 8484 21372
rect 8536 21360 8542 21412
rect 8662 21400 8668 21412
rect 8623 21372 8668 21400
rect 8662 21360 8668 21372
rect 8720 21360 8726 21412
rect 9398 21360 9404 21412
rect 9456 21400 9462 21412
rect 9906 21403 9964 21409
rect 9906 21400 9918 21403
rect 9456 21372 9918 21400
rect 9456 21360 9462 21372
rect 9906 21369 9918 21372
rect 9952 21400 9964 21403
rect 10042 21400 10048 21412
rect 9952 21372 10048 21400
rect 9952 21369 9964 21372
rect 9906 21363 9964 21369
rect 10042 21360 10048 21372
rect 10100 21360 10106 21412
rect 11383 21344 11411 21431
rect 12526 21400 12532 21412
rect 12487 21372 12532 21400
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 12618 21360 12624 21412
rect 12676 21400 12682 21412
rect 12676 21372 12721 21400
rect 12676 21360 12682 21372
rect 4571 21304 4844 21332
rect 7055 21335 7113 21341
rect 4571 21301 4583 21304
rect 4525 21295 4583 21301
rect 7055 21301 7067 21335
rect 7101 21332 7113 21335
rect 7558 21332 7564 21344
rect 7101 21304 7564 21332
rect 7101 21301 7113 21304
rect 7055 21295 7113 21301
rect 7558 21292 7564 21304
rect 7616 21292 7622 21344
rect 11330 21292 11336 21344
rect 11388 21332 11411 21344
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11388 21304 11805 21332
rect 11388 21292 11394 21304
rect 11793 21301 11805 21304
rect 11839 21332 11851 21335
rect 12434 21332 12440 21344
rect 11839 21304 12440 21332
rect 11839 21301 11851 21304
rect 11793 21295 11851 21301
rect 12434 21292 12440 21304
rect 12492 21292 12498 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 1394 21088 1400 21140
rect 1452 21128 1458 21140
rect 3418 21128 3424 21140
rect 1452 21100 3424 21128
rect 1452 21088 1458 21100
rect 3418 21088 3424 21100
rect 3476 21128 3482 21140
rect 7374 21128 7380 21140
rect 3476 21100 7380 21128
rect 3476 21088 3482 21100
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 7466 21088 7472 21140
rect 7524 21128 7530 21140
rect 7926 21128 7932 21140
rect 7524 21100 7569 21128
rect 7887 21100 7932 21128
rect 7524 21088 7530 21100
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 8110 21128 8116 21140
rect 8071 21100 8116 21128
rect 8110 21088 8116 21100
rect 8168 21088 8174 21140
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 9033 21131 9091 21137
rect 9033 21128 9045 21131
rect 8720 21100 9045 21128
rect 8720 21088 8726 21100
rect 9033 21097 9045 21100
rect 9079 21097 9091 21131
rect 10042 21128 10048 21140
rect 10003 21100 10048 21128
rect 9033 21091 9091 21097
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 10597 21131 10655 21137
rect 10597 21097 10609 21131
rect 10643 21128 10655 21131
rect 12437 21131 12495 21137
rect 12437 21128 12449 21131
rect 10643 21100 12449 21128
rect 10643 21097 10655 21100
rect 10597 21091 10655 21097
rect 12437 21097 12449 21100
rect 12483 21128 12495 21131
rect 12618 21128 12624 21140
rect 12483 21100 12624 21128
rect 12483 21097 12495 21100
rect 12437 21091 12495 21097
rect 12618 21088 12624 21100
rect 12676 21088 12682 21140
rect 4246 21020 4252 21072
rect 4304 21060 4310 21072
rect 4430 21060 4436 21072
rect 4304 21032 4436 21060
rect 4304 21020 4310 21032
rect 4430 21020 4436 21032
rect 4488 21020 4494 21072
rect 7193 21063 7251 21069
rect 7193 21029 7205 21063
rect 7239 21060 7251 21063
rect 9674 21060 9680 21072
rect 7239 21032 9680 21060
rect 7239 21029 7251 21032
rect 7193 21023 7251 21029
rect 9674 21020 9680 21032
rect 9732 21020 9738 21072
rect 10778 21020 10784 21072
rect 10836 21060 10842 21072
rect 11609 21063 11667 21069
rect 11609 21060 11621 21063
rect 10836 21032 11621 21060
rect 10836 21020 10842 21032
rect 11609 21029 11621 21032
rect 11655 21060 11667 21063
rect 11698 21060 11704 21072
rect 11655 21032 11704 21060
rect 11655 21029 11667 21032
rect 11609 21023 11667 21029
rect 11698 21020 11704 21032
rect 11756 21020 11762 21072
rect 4890 20992 4896 21004
rect 4851 20964 4896 20992
rect 4890 20952 4896 20964
rect 4948 20952 4954 21004
rect 6178 20952 6184 21004
rect 6236 20992 6242 21004
rect 6457 20995 6515 21001
rect 6457 20992 6469 20995
rect 6236 20964 6469 20992
rect 6236 20952 6242 20964
rect 6457 20961 6469 20964
rect 6503 20961 6515 20995
rect 6457 20955 6515 20961
rect 4430 20924 4436 20936
rect 4391 20896 4436 20924
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 6472 20924 6500 20955
rect 6546 20952 6552 21004
rect 6604 20992 6610 21004
rect 7009 20995 7067 21001
rect 7009 20992 7021 20995
rect 6604 20964 7021 20992
rect 6604 20952 6610 20964
rect 7009 20961 7021 20964
rect 7055 20992 7067 20995
rect 7466 20992 7472 21004
rect 7055 20964 7472 20992
rect 7055 20961 7067 20964
rect 7009 20955 7067 20961
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 8018 20992 8024 21004
rect 7979 20964 8024 20992
rect 8018 20952 8024 20964
rect 8076 20952 8082 21004
rect 8478 20992 8484 21004
rect 8439 20964 8484 20992
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 13056 20995 13114 21001
rect 13056 20961 13068 20995
rect 13102 20992 13114 20995
rect 13262 20992 13268 21004
rect 13102 20964 13268 20992
rect 13102 20961 13114 20964
rect 13056 20955 13114 20961
rect 13262 20952 13268 20964
rect 13320 20952 13326 21004
rect 9306 20924 9312 20936
rect 6472 20896 9312 20924
rect 9306 20884 9312 20896
rect 9364 20884 9370 20936
rect 9674 20924 9680 20936
rect 9635 20896 9680 20924
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11204 20896 11529 20924
rect 11204 20884 11210 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 13170 20924 13176 20936
rect 11517 20887 11575 20893
rect 13142 20884 13176 20924
rect 13228 20884 13234 20936
rect 12066 20856 12072 20868
rect 12027 20828 12072 20856
rect 12066 20816 12072 20828
rect 12124 20816 12130 20868
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9582 20788 9588 20800
rect 9539 20760 9588 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9582 20748 9588 20760
rect 9640 20788 9646 20800
rect 10042 20788 10048 20800
rect 9640 20760 10048 20788
rect 9640 20748 9646 20760
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10962 20788 10968 20800
rect 10923 20760 10968 20788
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11514 20788 11520 20800
rect 11112 20760 11520 20788
rect 11112 20748 11118 20760
rect 11514 20748 11520 20760
rect 11572 20788 11578 20800
rect 12526 20788 12532 20800
rect 11572 20760 12532 20788
rect 11572 20748 11578 20760
rect 12526 20748 12532 20760
rect 12584 20788 12590 20800
rect 13142 20797 13170 20884
rect 12805 20791 12863 20797
rect 12805 20788 12817 20791
rect 12584 20760 12817 20788
rect 12584 20748 12590 20760
rect 12805 20757 12817 20760
rect 12851 20757 12863 20791
rect 12805 20751 12863 20757
rect 13127 20791 13185 20797
rect 13127 20757 13139 20791
rect 13173 20757 13185 20791
rect 13127 20751 13185 20757
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 4249 20587 4307 20593
rect 4249 20553 4261 20587
rect 4295 20584 4307 20587
rect 4430 20584 4436 20596
rect 4295 20556 4436 20584
rect 4295 20553 4307 20556
rect 4249 20547 4307 20553
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4890 20544 4896 20596
rect 4948 20584 4954 20596
rect 5353 20587 5411 20593
rect 5353 20584 5365 20587
rect 4948 20556 5365 20584
rect 4948 20544 4954 20556
rect 5353 20553 5365 20556
rect 5399 20553 5411 20587
rect 5718 20584 5724 20596
rect 5679 20556 5724 20584
rect 5353 20547 5411 20553
rect 5718 20544 5724 20556
rect 5776 20544 5782 20596
rect 6546 20584 6552 20596
rect 6507 20556 6552 20584
rect 6546 20544 6552 20556
rect 6604 20584 6610 20596
rect 7193 20587 7251 20593
rect 7193 20584 7205 20587
rect 6604 20556 7205 20584
rect 6604 20544 6610 20556
rect 7193 20553 7205 20556
rect 7239 20553 7251 20587
rect 7193 20547 7251 20553
rect 4982 20516 4988 20528
rect 4943 20488 4988 20516
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 7208 20448 7236 20547
rect 8018 20544 8024 20596
rect 8076 20584 8082 20596
rect 8389 20587 8447 20593
rect 8389 20584 8401 20587
rect 8076 20556 8401 20584
rect 8076 20544 8082 20556
rect 8389 20553 8401 20556
rect 8435 20553 8447 20587
rect 8389 20547 8447 20553
rect 8849 20587 8907 20593
rect 8849 20553 8861 20587
rect 8895 20584 8907 20587
rect 9398 20584 9404 20596
rect 8895 20556 9404 20584
rect 8895 20553 8907 20556
rect 8849 20547 8907 20553
rect 9398 20544 9404 20556
rect 9456 20584 9462 20596
rect 10137 20587 10195 20593
rect 10137 20584 10149 20587
rect 9456 20556 10149 20584
rect 9456 20544 9462 20556
rect 10137 20553 10149 20556
rect 10183 20553 10195 20587
rect 11698 20584 11704 20596
rect 11659 20556 11704 20584
rect 10137 20547 10195 20553
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 11974 20544 11980 20596
rect 12032 20584 12038 20596
rect 12575 20587 12633 20593
rect 12575 20584 12587 20587
rect 12032 20556 12587 20584
rect 12032 20544 12038 20556
rect 12575 20553 12587 20556
rect 12621 20553 12633 20587
rect 13262 20584 13268 20596
rect 13223 20556 13268 20584
rect 12575 20547 12633 20553
rect 13262 20544 13268 20556
rect 13320 20544 13326 20596
rect 13906 20584 13912 20596
rect 13867 20556 13912 20584
rect 13906 20544 13912 20556
rect 13964 20544 13970 20596
rect 11146 20476 11152 20528
rect 11204 20516 11210 20528
rect 11333 20519 11391 20525
rect 11333 20516 11345 20519
rect 11204 20488 11345 20516
rect 11204 20476 11210 20488
rect 11333 20485 11345 20488
rect 11379 20516 11391 20519
rect 12069 20519 12127 20525
rect 12069 20516 12081 20519
rect 11379 20488 12081 20516
rect 11379 20485 11391 20488
rect 11333 20479 11391 20485
rect 12069 20485 12081 20488
rect 12115 20485 12127 20519
rect 12069 20479 12127 20485
rect 7208 20420 7880 20448
rect 5718 20340 5724 20392
rect 5776 20380 5782 20392
rect 7374 20380 7380 20392
rect 5776 20352 7380 20380
rect 5776 20340 5782 20352
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 7852 20389 7880 20420
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 8941 20451 8999 20457
rect 8941 20448 8953 20451
rect 8720 20420 8953 20448
rect 8720 20408 8726 20420
rect 8941 20417 8953 20420
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 10962 20448 10968 20460
rect 10827 20420 10968 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 10962 20408 10968 20420
rect 11020 20448 11026 20460
rect 13587 20451 13645 20457
rect 13587 20448 13599 20451
rect 11020 20420 13599 20448
rect 11020 20408 11026 20420
rect 13587 20417 13599 20420
rect 13633 20417 13645 20451
rect 13587 20411 13645 20417
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 9674 20380 9680 20392
rect 8159 20352 9680 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 9674 20340 9680 20352
rect 9732 20340 9738 20392
rect 9861 20383 9919 20389
rect 9861 20349 9873 20383
rect 9907 20380 9919 20383
rect 12342 20380 12348 20392
rect 9907 20352 10640 20380
rect 12303 20352 12348 20380
rect 9907 20349 9919 20352
rect 9861 20343 9919 20349
rect 4433 20315 4491 20321
rect 4433 20312 4445 20315
rect 4126 20284 4445 20312
rect 3329 20247 3387 20253
rect 3329 20213 3341 20247
rect 3375 20244 3387 20247
rect 3789 20247 3847 20253
rect 3789 20244 3801 20247
rect 3375 20216 3801 20244
rect 3375 20213 3387 20216
rect 3329 20207 3387 20213
rect 3789 20213 3801 20216
rect 3835 20244 3847 20247
rect 4126 20244 4154 20284
rect 4433 20281 4445 20284
rect 4479 20281 4491 20315
rect 4433 20275 4491 20281
rect 4522 20272 4528 20324
rect 4580 20312 4586 20324
rect 9303 20315 9361 20321
rect 4580 20284 4625 20312
rect 4580 20272 4586 20284
rect 9303 20281 9315 20315
rect 9349 20312 9361 20315
rect 9398 20312 9404 20324
rect 9349 20284 9404 20312
rect 9349 20281 9361 20284
rect 9303 20275 9361 20281
rect 9398 20272 9404 20284
rect 9456 20272 9462 20324
rect 3835 20216 4154 20244
rect 3835 20213 3847 20216
rect 3789 20207 3847 20213
rect 5350 20204 5356 20256
rect 5408 20244 5414 20256
rect 6089 20247 6147 20253
rect 6089 20244 6101 20247
rect 5408 20216 6101 20244
rect 5408 20204 5414 20216
rect 6089 20213 6101 20216
rect 6135 20244 6147 20247
rect 6178 20244 6184 20256
rect 6135 20216 6184 20244
rect 6135 20213 6147 20216
rect 6089 20207 6147 20213
rect 6178 20204 6184 20216
rect 6236 20204 6242 20256
rect 10612 20253 10640 20352
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 12710 20340 12716 20392
rect 12768 20380 12774 20392
rect 13500 20383 13558 20389
rect 13500 20380 13512 20383
rect 12768 20352 13512 20380
rect 12768 20340 12774 20352
rect 13500 20349 13512 20352
rect 13546 20380 13558 20383
rect 13906 20380 13912 20392
rect 13546 20352 13912 20380
rect 13546 20349 13558 20352
rect 13500 20343 13558 20349
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 10873 20315 10931 20321
rect 10873 20281 10885 20315
rect 10919 20312 10931 20315
rect 10962 20312 10968 20324
rect 10919 20284 10968 20312
rect 10919 20281 10931 20284
rect 10873 20275 10931 20281
rect 10597 20247 10655 20253
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 10888 20244 10916 20275
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 12360 20312 12388 20340
rect 12897 20315 12955 20321
rect 12897 20312 12909 20315
rect 12360 20284 12909 20312
rect 12897 20281 12909 20284
rect 12943 20281 12955 20315
rect 12897 20275 12955 20281
rect 10643 20216 10916 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 7742 20040 7748 20052
rect 6472 20012 7748 20040
rect 106 19932 112 19984
rect 164 19972 170 19984
rect 3099 19975 3157 19981
rect 3099 19972 3111 19975
rect 164 19944 3111 19972
rect 164 19932 170 19944
rect 3099 19941 3111 19944
rect 3145 19941 3157 19975
rect 4982 19972 4988 19984
rect 3099 19935 3157 19941
rect 4126 19944 4988 19972
rect 2958 19904 2964 19916
rect 2922 19876 2964 19904
rect 2958 19864 2964 19876
rect 3016 19913 3022 19916
rect 3016 19907 3070 19913
rect 3016 19873 3024 19907
rect 3058 19904 3070 19907
rect 4126 19904 4154 19944
rect 4982 19932 4988 19944
rect 5040 19932 5046 19984
rect 4890 19904 4896 19916
rect 3058 19876 4154 19904
rect 4851 19876 4896 19904
rect 3058 19873 3070 19876
rect 3016 19867 3070 19873
rect 3016 19864 3022 19867
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 6270 19864 6276 19916
rect 6328 19904 6334 19916
rect 6472 19913 6500 20012
rect 7484 19913 7512 20012
rect 7742 20000 7748 20012
rect 7800 20040 7806 20052
rect 8294 20040 8300 20052
rect 7800 20012 8300 20040
rect 7800 20000 7806 20012
rect 8294 20000 8300 20012
rect 8352 20040 8358 20052
rect 8389 20043 8447 20049
rect 8389 20040 8401 20043
rect 8352 20012 8401 20040
rect 8352 20000 8358 20012
rect 8389 20009 8401 20012
rect 8435 20009 8447 20043
rect 8389 20003 8447 20009
rect 9493 20043 9551 20049
rect 9493 20009 9505 20043
rect 9539 20040 9551 20043
rect 9674 20040 9680 20052
rect 9539 20012 9680 20040
rect 9539 20009 9551 20012
rect 9493 20003 9551 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 12158 20040 12164 20052
rect 11931 20012 12164 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 10410 19972 10416 19984
rect 7616 19944 10416 19972
rect 7616 19932 7622 19944
rect 10410 19932 10416 19944
rect 10468 19932 10474 19984
rect 10505 19975 10563 19981
rect 10505 19941 10517 19975
rect 10551 19972 10563 19975
rect 10870 19972 10876 19984
rect 10551 19944 10876 19972
rect 10551 19941 10563 19944
rect 10505 19935 10563 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 11054 19972 11060 19984
rect 11015 19944 11060 19972
rect 11054 19932 11060 19944
rect 11112 19932 11118 19984
rect 6457 19907 6515 19913
rect 6457 19904 6469 19907
rect 6328 19876 6469 19904
rect 6328 19864 6334 19876
rect 6457 19873 6469 19876
rect 6503 19873 6515 19907
rect 6457 19867 6515 19873
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19904 7159 19907
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 7147 19876 7389 19904
rect 7147 19873 7159 19876
rect 7101 19867 7159 19873
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 7469 19907 7527 19913
rect 7469 19873 7481 19907
rect 7515 19873 7527 19907
rect 7469 19867 7527 19873
rect 7653 19907 7711 19913
rect 7653 19873 7665 19907
rect 7699 19904 7711 19907
rect 7742 19904 7748 19916
rect 7699 19876 7748 19904
rect 7699 19873 7711 19876
rect 7653 19867 7711 19873
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 8478 19864 8484 19916
rect 8536 19904 8542 19916
rect 9953 19907 10011 19913
rect 9953 19904 9965 19907
rect 8536 19876 9965 19904
rect 8536 19864 8542 19876
rect 9953 19873 9965 19876
rect 9999 19904 10011 19907
rect 10226 19904 10232 19916
rect 9999 19876 10232 19904
rect 9999 19873 10011 19876
rect 9953 19867 10011 19873
rect 10226 19864 10232 19876
rect 10284 19864 10290 19916
rect 4982 19836 4988 19848
rect 4895 19808 4988 19836
rect 4982 19796 4988 19808
rect 5040 19836 5046 19848
rect 7834 19836 7840 19848
rect 5040 19808 7604 19836
rect 7795 19808 7840 19836
rect 5040 19796 5046 19808
rect 5994 19728 6000 19780
rect 6052 19768 6058 19780
rect 6822 19768 6828 19780
rect 6052 19740 6828 19768
rect 6052 19728 6058 19740
rect 6822 19728 6828 19740
rect 6880 19768 6886 19780
rect 7101 19771 7159 19777
rect 7101 19768 7113 19771
rect 6880 19740 7113 19768
rect 6880 19728 6886 19740
rect 7101 19737 7113 19740
rect 7147 19768 7159 19771
rect 7193 19771 7251 19777
rect 7193 19768 7205 19771
rect 7147 19740 7205 19768
rect 7147 19737 7159 19740
rect 7101 19731 7159 19737
rect 7193 19737 7205 19740
rect 7239 19737 7251 19771
rect 7576 19768 7604 19808
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 7576 19740 8708 19768
rect 7193 19731 7251 19737
rect 8680 19712 8708 19740
rect 5258 19700 5264 19712
rect 5219 19672 5264 19700
rect 5258 19660 5264 19672
rect 5316 19700 5322 19712
rect 6086 19700 6092 19712
rect 5316 19672 6092 19700
rect 5316 19660 5322 19672
rect 6086 19660 6092 19672
rect 6144 19660 6150 19712
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 8757 19703 8815 19709
rect 8757 19700 8769 19703
rect 8720 19672 8769 19700
rect 8720 19660 8726 19672
rect 8757 19669 8769 19672
rect 8803 19669 8815 19703
rect 8757 19663 8815 19669
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 2958 19496 2964 19508
rect 2919 19468 2964 19496
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 4706 19456 4712 19508
rect 4764 19496 4770 19508
rect 4985 19499 5043 19505
rect 4985 19496 4997 19499
rect 4764 19468 4997 19496
rect 4764 19456 4770 19468
rect 4985 19465 4997 19468
rect 5031 19496 5043 19499
rect 8205 19499 8263 19505
rect 8205 19496 8217 19499
rect 5031 19468 8217 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 8205 19465 8217 19468
rect 8251 19465 8263 19499
rect 10962 19496 10968 19508
rect 10923 19468 10968 19496
rect 8205 19459 8263 19465
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19360 4123 19363
rect 4111 19332 4752 19360
rect 4111 19329 4123 19332
rect 4065 19323 4123 19329
rect 3697 19295 3755 19301
rect 3697 19261 3709 19295
rect 3743 19292 3755 19295
rect 4154 19292 4160 19304
rect 3743 19264 4160 19292
rect 3743 19261 3755 19264
rect 3697 19255 3755 19261
rect 4154 19252 4160 19264
rect 4212 19292 4218 19304
rect 4212 19264 4257 19292
rect 4212 19252 4218 19264
rect 4724 19233 4752 19332
rect 5000 19292 5028 19459
rect 5258 19428 5264 19440
rect 5219 19400 5264 19428
rect 5258 19388 5264 19400
rect 5316 19388 5322 19440
rect 6270 19428 6276 19440
rect 6231 19400 6276 19428
rect 6270 19388 6276 19400
rect 6328 19388 6334 19440
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 6917 19363 6975 19369
rect 6917 19360 6929 19363
rect 6144 19332 6929 19360
rect 6144 19320 6150 19332
rect 6917 19329 6929 19332
rect 6963 19329 6975 19363
rect 6917 19323 6975 19329
rect 5166 19292 5172 19304
rect 5000 19264 5172 19292
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19261 5503 19295
rect 6822 19292 6828 19304
rect 6783 19264 6828 19292
rect 5445 19255 5503 19261
rect 4709 19227 4767 19233
rect 4709 19193 4721 19227
rect 4755 19224 4767 19227
rect 4890 19224 4896 19236
rect 4755 19196 4896 19224
rect 4755 19193 4767 19196
rect 4709 19187 4767 19193
rect 4890 19184 4896 19196
rect 4948 19224 4954 19236
rect 5460 19224 5488 19255
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 7101 19295 7159 19301
rect 7101 19292 7113 19295
rect 6932 19264 7113 19292
rect 6932 19236 6960 19264
rect 7101 19261 7113 19264
rect 7147 19292 7159 19295
rect 7742 19292 7748 19304
rect 7147 19264 7748 19292
rect 7147 19261 7159 19264
rect 7101 19255 7159 19261
rect 7742 19252 7748 19264
rect 7800 19292 7806 19304
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 7800 19264 7849 19292
rect 7800 19252 7806 19264
rect 7837 19261 7849 19264
rect 7883 19261 7895 19295
rect 8220 19292 8248 19459
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 8294 19388 8300 19440
rect 8352 19428 8358 19440
rect 8481 19431 8539 19437
rect 8481 19428 8493 19431
rect 8352 19400 8493 19428
rect 8352 19388 8358 19400
rect 8481 19397 8493 19400
rect 8527 19397 8539 19431
rect 8481 19391 8539 19397
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8220 19264 8401 19292
rect 7837 19255 7895 19261
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8662 19292 8668 19304
rect 8623 19264 8668 19292
rect 8389 19255 8447 19261
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 9916 19264 9965 19292
rect 9916 19252 9922 19264
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 10226 19252 10232 19304
rect 10284 19292 10290 19304
rect 10413 19295 10471 19301
rect 10413 19292 10425 19295
rect 10284 19264 10425 19292
rect 10284 19252 10290 19264
rect 10413 19261 10425 19264
rect 10459 19261 10471 19295
rect 10413 19255 10471 19261
rect 6641 19227 6699 19233
rect 6641 19224 6653 19227
rect 4948 19196 6653 19224
rect 4948 19184 4954 19196
rect 6641 19193 6653 19196
rect 6687 19224 6699 19227
rect 6914 19224 6920 19236
rect 6687 19196 6920 19224
rect 6687 19193 6699 19196
rect 6641 19187 6699 19193
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 7561 19227 7619 19233
rect 7561 19193 7573 19227
rect 7607 19224 7619 19227
rect 10686 19224 10692 19236
rect 7607 19196 10692 19224
rect 7607 19193 7619 19196
rect 7561 19187 7619 19193
rect 10686 19184 10692 19196
rect 10744 19184 10750 19236
rect 4341 19159 4399 19165
rect 4341 19125 4353 19159
rect 4387 19156 4399 19159
rect 5442 19156 5448 19168
rect 4387 19128 5448 19156
rect 4387 19125 4399 19128
rect 4341 19119 4399 19125
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 5626 19156 5632 19168
rect 5587 19128 5632 19156
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 9364 19128 9781 19156
rect 9364 19116 9370 19128
rect 9769 19125 9781 19128
rect 9815 19156 9827 19159
rect 9858 19156 9864 19168
rect 9815 19128 9864 19156
rect 9815 19125 9827 19128
rect 9769 19119 9827 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 4154 18912 4160 18964
rect 4212 18952 4218 18964
rect 5169 18955 5227 18961
rect 5169 18952 5181 18955
rect 4212 18924 5181 18952
rect 4212 18912 4218 18924
rect 5169 18921 5181 18924
rect 5215 18921 5227 18955
rect 5810 18952 5816 18964
rect 5771 18924 5816 18952
rect 5169 18915 5227 18921
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 6086 18952 6092 18964
rect 6047 18924 6092 18952
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 7469 18955 7527 18961
rect 7469 18921 7481 18955
rect 7515 18952 7527 18955
rect 8294 18952 8300 18964
rect 7515 18924 8300 18952
rect 7515 18921 7527 18924
rect 7469 18915 7527 18921
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 9861 18955 9919 18961
rect 9861 18952 9873 18955
rect 8588 18924 9873 18952
rect 4617 18887 4675 18893
rect 4617 18853 4629 18887
rect 4663 18884 4675 18887
rect 6822 18884 6828 18896
rect 4663 18856 6828 18884
rect 4663 18853 4675 18856
rect 4617 18847 4675 18853
rect 4724 18825 4752 18856
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 7929 18887 7987 18893
rect 7929 18853 7941 18887
rect 7975 18884 7987 18887
rect 8588 18884 8616 18924
rect 9861 18921 9873 18924
rect 9907 18921 9919 18955
rect 10410 18952 10416 18964
rect 10371 18924 10416 18952
rect 9861 18915 9919 18921
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 7975 18856 8616 18884
rect 7975 18853 7987 18856
rect 7929 18847 7987 18853
rect 4709 18819 4767 18825
rect 4709 18816 4721 18819
rect 4687 18788 4721 18816
rect 4709 18785 4721 18788
rect 4755 18785 4767 18819
rect 4982 18816 4988 18828
rect 4943 18788 4988 18816
rect 4709 18779 4767 18785
rect 4982 18776 4988 18788
rect 5040 18776 5046 18828
rect 5166 18776 5172 18828
rect 5224 18816 5230 18828
rect 6270 18816 6276 18828
rect 5224 18788 6276 18816
rect 5224 18776 5230 18788
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18816 6607 18819
rect 6914 18816 6920 18828
rect 6595 18788 6920 18816
rect 6595 18785 6607 18788
rect 6549 18779 6607 18785
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 7558 18816 7564 18828
rect 7432 18788 7564 18816
rect 7432 18776 7438 18788
rect 7558 18776 7564 18788
rect 7616 18816 7622 18828
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7616 18788 8033 18816
rect 7616 18776 7622 18788
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8478 18776 8484 18828
rect 8536 18816 8542 18828
rect 8588 18825 8616 18856
rect 8573 18819 8631 18825
rect 8573 18816 8585 18819
rect 8536 18788 8585 18816
rect 8536 18776 8542 18788
rect 8573 18785 8585 18788
rect 8619 18785 8631 18819
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 8573 18779 8631 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10686 18816 10692 18828
rect 10647 18788 10692 18816
rect 10686 18776 10692 18788
rect 10744 18776 10750 18828
rect 4062 18708 4068 18760
rect 4120 18748 4126 18760
rect 5000 18748 5028 18776
rect 4120 18720 5028 18748
rect 4120 18708 4126 18720
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 6236 18720 6377 18748
rect 6236 18708 6242 18720
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18748 7067 18751
rect 8202 18748 8208 18760
rect 7055 18720 8208 18748
rect 7055 18717 7067 18720
rect 7009 18711 7067 18717
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 9582 18748 9588 18760
rect 8803 18720 9588 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 11514 18708 11520 18760
rect 11572 18748 11578 18760
rect 11701 18751 11759 18757
rect 11701 18748 11713 18751
rect 11572 18720 11713 18748
rect 11572 18708 11578 18720
rect 11701 18717 11713 18720
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 4798 18680 4804 18692
rect 4711 18652 4804 18680
rect 4798 18640 4804 18652
rect 4856 18680 4862 18692
rect 6196 18680 6224 18708
rect 4856 18652 6224 18680
rect 4856 18640 4862 18652
rect 5442 18572 5448 18624
rect 5500 18612 5506 18624
rect 7374 18612 7380 18624
rect 5500 18584 7380 18612
rect 5500 18572 5506 18584
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 7466 18572 7472 18624
rect 7524 18612 7530 18624
rect 10873 18615 10931 18621
rect 10873 18612 10885 18615
rect 7524 18584 10885 18612
rect 7524 18572 7530 18584
rect 10873 18581 10885 18584
rect 10919 18581 10931 18615
rect 10873 18575 10931 18581
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 2869 18411 2927 18417
rect 2869 18377 2881 18411
rect 2915 18408 2927 18411
rect 8846 18408 8852 18420
rect 2915 18380 8852 18408
rect 2915 18377 2927 18380
rect 2869 18371 2927 18377
rect 2976 18213 3004 18380
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 9309 18411 9367 18417
rect 9309 18377 9321 18411
rect 9355 18408 9367 18411
rect 9398 18408 9404 18420
rect 9355 18380 9404 18408
rect 9355 18377 9367 18380
rect 9309 18371 9367 18377
rect 9398 18368 9404 18380
rect 9456 18408 9462 18420
rect 9766 18408 9772 18420
rect 9456 18380 9772 18408
rect 9456 18368 9462 18380
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 10686 18408 10692 18420
rect 10647 18380 10692 18408
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 3881 18343 3939 18349
rect 3881 18309 3893 18343
rect 3927 18340 3939 18343
rect 4062 18340 4068 18352
rect 3927 18312 4068 18340
rect 3927 18309 3939 18312
rect 3881 18303 3939 18309
rect 4062 18300 4068 18312
rect 4120 18300 4126 18352
rect 4798 18340 4804 18352
rect 4759 18312 4804 18340
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 6270 18340 6276 18352
rect 6231 18312 6276 18340
rect 6270 18300 6276 18312
rect 6328 18300 6334 18352
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 7742 18340 7748 18352
rect 7432 18312 7748 18340
rect 7432 18300 7438 18312
rect 7742 18300 7748 18312
rect 7800 18340 7806 18352
rect 7800 18312 9806 18340
rect 7800 18300 7806 18312
rect 5810 18272 5816 18284
rect 5276 18244 5816 18272
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18173 3019 18207
rect 2961 18167 3019 18173
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3970 18204 3976 18216
rect 3559 18176 3976 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 5276 18213 5304 18244
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 5902 18232 5908 18284
rect 5960 18272 5966 18284
rect 8849 18275 8907 18281
rect 8849 18272 8861 18275
rect 5960 18244 8861 18272
rect 5960 18232 5966 18244
rect 8849 18241 8861 18244
rect 8895 18272 8907 18275
rect 9674 18272 9680 18284
rect 8895 18244 9680 18272
rect 8895 18241 8907 18244
rect 8849 18235 8907 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 5261 18207 5319 18213
rect 5261 18173 5273 18207
rect 5307 18173 5319 18207
rect 5261 18167 5319 18173
rect 5445 18207 5503 18213
rect 5445 18173 5457 18207
rect 5491 18173 5503 18207
rect 5445 18167 5503 18173
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 7006 18204 7012 18216
rect 6871 18176 7012 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 4798 18096 4804 18148
rect 4856 18136 4862 18148
rect 5460 18136 5488 18167
rect 7006 18164 7012 18176
rect 7064 18204 7070 18216
rect 7466 18204 7472 18216
rect 7064 18176 7472 18204
rect 7064 18164 7070 18176
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7607 18176 7849 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 8478 18204 8484 18216
rect 8435 18176 8484 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 7374 18136 7380 18148
rect 4856 18108 5488 18136
rect 7287 18108 7380 18136
rect 4856 18096 4862 18108
rect 7374 18096 7380 18108
rect 7432 18136 7438 18148
rect 8404 18136 8432 18167
rect 8478 18164 8484 18176
rect 8536 18164 8542 18216
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 9398 18204 9404 18216
rect 8619 18176 9404 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9778 18204 9806 18312
rect 9858 18300 9864 18352
rect 9916 18340 9922 18352
rect 11333 18343 11391 18349
rect 11333 18340 11345 18343
rect 9916 18312 11345 18340
rect 9916 18300 9922 18312
rect 11333 18309 11345 18312
rect 11379 18309 11391 18343
rect 11333 18303 11391 18309
rect 11149 18207 11207 18213
rect 11149 18204 11161 18207
rect 9778 18176 11161 18204
rect 11149 18173 11161 18176
rect 11195 18204 11207 18207
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 11195 18176 11621 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 11609 18173 11621 18176
rect 11655 18173 11667 18207
rect 11609 18167 11667 18173
rect 9306 18136 9312 18148
rect 7432 18108 8432 18136
rect 9140 18108 9312 18136
rect 7432 18096 7438 18108
rect 3145 18071 3203 18077
rect 3145 18037 3157 18071
rect 3191 18068 3203 18071
rect 4062 18068 4068 18080
rect 3191 18040 4068 18068
rect 3191 18037 3203 18040
rect 3145 18031 3203 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4157 18071 4215 18077
rect 4157 18037 4169 18071
rect 4203 18068 4215 18071
rect 4522 18068 4528 18080
rect 4203 18040 4528 18068
rect 4203 18037 4215 18040
rect 4157 18031 4215 18037
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 5074 18068 5080 18080
rect 5035 18040 5080 18068
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 7009 18071 7067 18077
rect 7009 18068 7021 18071
rect 5868 18040 7021 18068
rect 5868 18028 5874 18040
rect 7009 18037 7021 18040
rect 7055 18068 7067 18071
rect 7561 18071 7619 18077
rect 7561 18068 7573 18071
rect 7055 18040 7573 18068
rect 7055 18037 7067 18040
rect 7009 18031 7067 18037
rect 7561 18037 7573 18040
rect 7607 18068 7619 18071
rect 7653 18071 7711 18077
rect 7653 18068 7665 18071
rect 7607 18040 7665 18068
rect 7607 18037 7619 18040
rect 7561 18031 7619 18037
rect 7653 18037 7665 18040
rect 7699 18068 7711 18071
rect 9140 18068 9168 18108
rect 9306 18096 9312 18108
rect 9364 18096 9370 18148
rect 9766 18068 9772 18080
rect 7699 18040 9168 18068
rect 9727 18040 9772 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 5258 17864 5264 17876
rect 5219 17836 5264 17864
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 6641 17867 6699 17873
rect 6641 17864 6653 17867
rect 6236 17836 6653 17864
rect 6236 17824 6242 17836
rect 6641 17833 6653 17836
rect 6687 17833 6699 17867
rect 7006 17864 7012 17876
rect 6967 17836 7012 17864
rect 6641 17827 6699 17833
rect 7006 17824 7012 17836
rect 7064 17864 7070 17876
rect 7190 17864 7196 17876
rect 7064 17836 7196 17864
rect 7064 17824 7070 17836
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 9398 17864 9404 17876
rect 9359 17836 9404 17864
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 9824 17836 10041 17864
rect 9824 17824 9830 17836
rect 6365 17799 6423 17805
rect 6365 17765 6377 17799
rect 6411 17796 6423 17799
rect 6914 17796 6920 17808
rect 6411 17768 6920 17796
rect 6411 17765 6423 17768
rect 6365 17759 6423 17765
rect 6914 17756 6920 17768
rect 6972 17756 6978 17808
rect 8481 17799 8539 17805
rect 8481 17796 8493 17799
rect 7576 17768 8493 17796
rect 7576 17740 7604 17768
rect 8481 17765 8493 17768
rect 8527 17796 8539 17799
rect 9858 17796 9864 17808
rect 8527 17768 9864 17796
rect 8527 17765 8539 17768
rect 8481 17759 8539 17765
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 10013 17805 10041 17836
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 11422 17864 11428 17876
rect 10376 17836 11428 17864
rect 10376 17824 10382 17836
rect 11422 17824 11428 17836
rect 11480 17864 11486 17876
rect 11480 17836 11652 17864
rect 11480 17824 11486 17836
rect 9998 17799 10056 17805
rect 9998 17765 10010 17799
rect 10044 17765 10056 17799
rect 11514 17796 11520 17808
rect 11475 17768 11520 17796
rect 9998 17759 10056 17765
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 11624 17805 11652 17836
rect 11609 17799 11667 17805
rect 11609 17765 11621 17799
rect 11655 17765 11667 17799
rect 11609 17759 11667 17765
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17697 3019 17731
rect 2961 17691 3019 17697
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 5074 17728 5080 17740
rect 4939 17700 5080 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 2976 17660 3004 17691
rect 5074 17688 5080 17700
rect 5132 17688 5138 17740
rect 7558 17728 7564 17740
rect 7519 17700 7564 17728
rect 7558 17688 7564 17700
rect 7616 17688 7622 17740
rect 7926 17728 7932 17740
rect 7887 17700 7932 17728
rect 7926 17688 7932 17700
rect 7984 17688 7990 17740
rect 9582 17688 9588 17740
rect 9640 17728 9646 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9640 17700 9689 17728
rect 9640 17688 9646 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 3050 17660 3056 17672
rect 2963 17632 3056 17660
rect 3050 17620 3056 17632
rect 3108 17660 3114 17672
rect 7650 17660 7656 17672
rect 3108 17632 7656 17660
rect 3108 17620 3114 17632
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 8018 17660 8024 17672
rect 7979 17632 8024 17660
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17660 12219 17663
rect 12802 17660 12808 17672
rect 12207 17632 12808 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 4430 17552 4436 17604
rect 4488 17592 4494 17604
rect 12710 17592 12716 17604
rect 4488 17564 12716 17592
rect 4488 17552 4494 17564
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 3145 17527 3203 17533
rect 3145 17493 3157 17527
rect 3191 17524 3203 17527
rect 4798 17524 4804 17536
rect 3191 17496 4804 17524
rect 3191 17493 3203 17496
rect 3145 17487 3203 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 5718 17484 5724 17536
rect 5776 17524 5782 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5776 17496 5825 17524
rect 5776 17484 5782 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 5813 17487 5871 17493
rect 10597 17527 10655 17533
rect 10597 17493 10609 17527
rect 10643 17524 10655 17527
rect 12158 17524 12164 17536
rect 10643 17496 12164 17524
rect 10643 17493 10655 17496
rect 10597 17487 10655 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 4617 17323 4675 17329
rect 4617 17289 4629 17323
rect 4663 17320 4675 17323
rect 5074 17320 5080 17332
rect 4663 17292 5080 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8352 17292 9045 17320
rect 8352 17280 8358 17292
rect 9033 17289 9045 17292
rect 9079 17320 9091 17323
rect 9766 17320 9772 17332
rect 9079 17292 9772 17320
rect 9079 17289 9091 17292
rect 9033 17283 9091 17289
rect 4249 17255 4307 17261
rect 4249 17252 4261 17255
rect 4126 17224 4261 17252
rect 4126 17184 4154 17224
rect 4249 17221 4261 17224
rect 4295 17252 4307 17255
rect 7834 17252 7840 17264
rect 4295 17224 7840 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 3712 17156 4154 17184
rect 3712 17125 3740 17156
rect 4522 17144 4528 17196
rect 4580 17184 4586 17196
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 4580 17156 6561 17184
rect 4580 17144 4586 17156
rect 6549 17153 6561 17156
rect 6595 17184 6607 17187
rect 7926 17184 7932 17196
rect 6595 17156 7932 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17085 3755 17119
rect 3697 17079 3755 17085
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4709 17119 4767 17125
rect 4709 17116 4721 17119
rect 4120 17088 4721 17116
rect 4120 17076 4126 17088
rect 4709 17085 4721 17088
rect 4755 17116 4767 17119
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 4755 17088 5549 17116
rect 4755 17085 4767 17088
rect 4709 17079 4767 17085
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 5552 17048 5580 17079
rect 5626 17076 5632 17128
rect 5684 17116 5690 17128
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 5684 17088 5733 17116
rect 5684 17076 5690 17088
rect 5721 17085 5733 17088
rect 5767 17116 5779 17119
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 5767 17088 6193 17116
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 6181 17085 6193 17088
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 7374 17076 7380 17128
rect 7432 17116 7438 17128
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 7432 17088 7573 17116
rect 7432 17076 7438 17088
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 7650 17076 7656 17128
rect 7708 17116 7714 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7708 17088 8033 17116
rect 7708 17076 7714 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 9122 17116 9128 17128
rect 8343 17088 9128 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 6914 17048 6920 17060
rect 5552 17020 6920 17048
rect 6914 17008 6920 17020
rect 6972 17008 6978 17060
rect 9502 17057 9530 17292
rect 9766 17280 9772 17292
rect 9824 17320 9830 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 9824 17292 10333 17320
rect 9824 17280 9830 17292
rect 10321 17289 10333 17292
rect 10367 17289 10379 17323
rect 10321 17283 10379 17289
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 11572 17292 11713 17320
rect 11572 17280 11578 17292
rect 11701 17289 11713 17292
rect 11747 17289 11759 17323
rect 12158 17320 12164 17332
rect 12119 17292 12164 17320
rect 11701 17283 11759 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12802 17184 12808 17196
rect 12763 17156 12808 17184
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 10045 17119 10103 17125
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 10778 17116 10784 17128
rect 10091 17088 10784 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 10870 17076 10876 17128
rect 10928 17125 10934 17128
rect 10928 17119 10966 17125
rect 10954 17116 10966 17119
rect 11333 17119 11391 17125
rect 11333 17116 11345 17119
rect 10954 17088 11345 17116
rect 10954 17085 10966 17088
rect 10928 17079 10966 17085
rect 11333 17085 11345 17088
rect 11379 17116 11391 17119
rect 12250 17116 12256 17128
rect 11379 17088 12256 17116
rect 11379 17085 11391 17088
rect 11333 17079 11391 17085
rect 10928 17076 10934 17079
rect 12250 17076 12256 17088
rect 12308 17076 12314 17128
rect 9487 17051 9545 17057
rect 9487 17017 9499 17051
rect 9533 17017 9545 17051
rect 9487 17011 9545 17017
rect 12066 17008 12072 17060
rect 12124 17048 12130 17060
rect 12526 17048 12532 17060
rect 12124 17020 12532 17048
rect 12124 17008 12130 17020
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17017 12679 17051
rect 12621 17011 12679 17017
rect 3881 16983 3939 16989
rect 3881 16949 3893 16983
rect 3927 16980 3939 16983
rect 3970 16980 3976 16992
rect 3927 16952 3976 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4890 16980 4896 16992
rect 4851 16952 4896 16980
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5902 16980 5908 16992
rect 5863 16952 5908 16980
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 7101 16983 7159 16989
rect 7101 16949 7113 16983
rect 7147 16980 7159 16983
rect 7558 16980 7564 16992
rect 7147 16952 7564 16980
rect 7147 16949 7159 16952
rect 7101 16943 7159 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 11011 16983 11069 16989
rect 11011 16949 11023 16983
rect 11057 16980 11069 16983
rect 11238 16980 11244 16992
rect 11057 16952 11244 16980
rect 11057 16949 11069 16952
rect 11011 16943 11069 16949
rect 11238 16940 11244 16952
rect 11296 16940 11302 16992
rect 12158 16940 12164 16992
rect 12216 16980 12222 16992
rect 12636 16980 12664 17011
rect 12216 16952 12664 16980
rect 12216 16940 12222 16952
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 5813 16779 5871 16785
rect 5813 16776 5825 16779
rect 4948 16748 5825 16776
rect 4948 16736 4954 16748
rect 2961 16643 3019 16649
rect 2961 16609 2973 16643
rect 3007 16640 3019 16643
rect 3050 16640 3056 16652
rect 3007 16612 3056 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 5000 16649 5028 16748
rect 5813 16745 5825 16748
rect 5859 16776 5871 16779
rect 7282 16776 7288 16788
rect 5859 16748 7288 16776
rect 5859 16745 5871 16748
rect 5813 16739 5871 16745
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 9122 16776 9128 16788
rect 9083 16748 9128 16776
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9582 16736 9588 16788
rect 9640 16776 9646 16788
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9640 16748 9873 16776
rect 9640 16736 9646 16748
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11480 16748 11529 16776
rect 11480 16736 11486 16748
rect 11517 16745 11529 16748
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 8199 16711 8257 16717
rect 5276 16680 6868 16708
rect 5276 16649 5304 16680
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 4985 16603 5043 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 6730 16640 6736 16652
rect 6595 16612 6736 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 6840 16649 6868 16680
rect 8199 16677 8211 16711
rect 8245 16708 8257 16711
rect 8294 16708 8300 16720
rect 8245 16680 8300 16708
rect 8245 16677 8257 16680
rect 8199 16671 8257 16677
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 10686 16708 10692 16720
rect 10647 16680 10692 16708
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 10778 16668 10784 16720
rect 10836 16708 10842 16720
rect 12158 16708 12164 16720
rect 10836 16680 12164 16708
rect 10836 16668 10842 16680
rect 12158 16668 12164 16680
rect 12216 16708 12222 16720
rect 12253 16711 12311 16717
rect 12253 16708 12265 16711
rect 12216 16680 12265 16708
rect 12216 16668 12222 16680
rect 12253 16677 12265 16680
rect 12299 16677 12311 16711
rect 12802 16708 12808 16720
rect 12763 16680 12808 16708
rect 12253 16671 12311 16677
rect 12802 16668 12808 16680
rect 12860 16668 12866 16720
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16640 6883 16643
rect 7374 16640 7380 16652
rect 6871 16612 7380 16640
rect 6871 16609 6883 16612
rect 6825 16603 6883 16609
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8018 16640 8024 16652
rect 7883 16612 8024 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 5442 16572 5448 16584
rect 5403 16544 5448 16572
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16572 7067 16575
rect 9674 16572 9680 16584
rect 7055 16544 9680 16572
rect 7055 16541 7067 16544
rect 7009 16535 7067 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 10594 16572 10600 16584
rect 10555 16544 10600 16572
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 11054 16572 11060 16584
rect 11015 16544 11060 16572
rect 11054 16532 11060 16544
rect 11112 16572 11118 16584
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 11112 16544 12173 16572
rect 11112 16532 11118 16544
rect 12161 16541 12173 16544
rect 12207 16572 12219 16575
rect 12894 16572 12900 16584
rect 12207 16544 12900 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 12894 16532 12900 16544
rect 12952 16532 12958 16584
rect 3142 16436 3148 16448
rect 3103 16408 3148 16436
rect 3142 16396 3148 16408
rect 3200 16396 3206 16448
rect 4617 16439 4675 16445
rect 4617 16405 4629 16439
rect 4663 16436 4675 16439
rect 4798 16436 4804 16448
rect 4663 16408 4804 16436
rect 4663 16405 4675 16408
rect 4617 16399 4675 16405
rect 4798 16396 4804 16408
rect 4856 16436 4862 16448
rect 5534 16436 5540 16448
rect 4856 16408 5540 16436
rect 4856 16396 4862 16408
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 5902 16396 5908 16448
rect 5960 16436 5966 16448
rect 7561 16439 7619 16445
rect 7561 16436 7573 16439
rect 5960 16408 7573 16436
rect 5960 16396 5966 16408
rect 7561 16405 7573 16408
rect 7607 16436 7619 16439
rect 7650 16436 7656 16448
rect 7607 16408 7656 16436
rect 7607 16405 7619 16408
rect 7561 16399 7619 16405
rect 7650 16396 7656 16408
rect 7708 16396 7714 16448
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16436 8815 16439
rect 9306 16436 9312 16448
rect 8803 16408 9312 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 4801 16235 4859 16241
rect 4801 16201 4813 16235
rect 4847 16232 4859 16235
rect 6365 16235 6423 16241
rect 6365 16232 6377 16235
rect 4847 16204 6377 16232
rect 4847 16201 4859 16204
rect 4801 16195 4859 16201
rect 6365 16201 6377 16204
rect 6411 16232 6423 16235
rect 7374 16232 7380 16244
rect 6411 16204 7380 16232
rect 6411 16201 6423 16204
rect 6365 16195 6423 16201
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8573 16235 8631 16241
rect 8573 16232 8585 16235
rect 8352 16204 8585 16232
rect 8352 16192 8358 16204
rect 8573 16201 8585 16204
rect 8619 16232 8631 16235
rect 8846 16232 8852 16244
rect 8619 16204 8852 16232
rect 8619 16201 8631 16204
rect 8573 16195 8631 16201
rect 8846 16192 8852 16204
rect 8904 16232 8910 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 8904 16204 8953 16232
rect 8904 16192 8910 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 6730 16164 6736 16176
rect 4295 16136 6736 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 6730 16124 6736 16136
rect 6788 16164 6794 16176
rect 7009 16167 7067 16173
rect 7009 16164 7021 16167
rect 6788 16136 7021 16164
rect 6788 16124 6794 16136
rect 7009 16133 7021 16136
rect 7055 16133 7067 16167
rect 7009 16127 7067 16133
rect 7834 16124 7840 16176
rect 7892 16164 7898 16176
rect 8110 16164 8116 16176
rect 7892 16136 8116 16164
rect 7892 16124 7898 16136
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 8956 16164 8984 16195
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 11011 16235 11069 16241
rect 11011 16232 11023 16235
rect 10652 16204 11023 16232
rect 10652 16192 10658 16204
rect 11011 16201 11023 16204
rect 11057 16232 11069 16235
rect 11701 16235 11759 16241
rect 11701 16232 11713 16235
rect 11057 16204 11713 16232
rect 11057 16201 11069 16204
rect 11011 16195 11069 16201
rect 11701 16201 11713 16204
rect 11747 16201 11759 16235
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 11701 16195 11759 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12575 16235 12633 16241
rect 12575 16201 12587 16235
rect 12621 16232 12633 16235
rect 14734 16232 14740 16244
rect 12621 16204 14740 16232
rect 12621 16201 12633 16204
rect 12575 16195 12633 16201
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 12894 16164 12900 16176
rect 8956 16136 9260 16164
rect 12855 16136 12900 16164
rect 5442 16056 5448 16108
rect 5500 16096 5506 16108
rect 9122 16096 9128 16108
rect 5500 16068 9128 16096
rect 5500 16056 5506 16068
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 3970 15988 3976 16040
rect 4028 16028 4034 16040
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 4028 16000 4077 16028
rect 4028 15988 4034 16000
rect 4065 15997 4077 16000
rect 4111 15997 4123 16031
rect 4065 15991 4123 15997
rect 3050 15892 3056 15904
rect 3011 15864 3056 15892
rect 3050 15852 3056 15864
rect 3108 15852 3114 15904
rect 3973 15895 4031 15901
rect 3973 15861 3985 15895
rect 4019 15892 4031 15895
rect 4080 15892 4108 15991
rect 4890 15988 4896 16040
rect 4948 16028 4954 16040
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 4948 16000 5089 16028
rect 4948 15988 4954 16000
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5534 16028 5540 16040
rect 5495 16000 5540 16028
rect 5077 15991 5135 15997
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 5810 15960 5816 15972
rect 5771 15932 5816 15960
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 7374 15920 7380 15972
rect 7432 15960 7438 15972
rect 8036 15960 8064 15991
rect 8294 15960 8300 15972
rect 7432 15932 8064 15960
rect 8255 15932 8300 15960
rect 7432 15920 7438 15932
rect 8294 15920 8300 15932
rect 8352 15920 8358 15972
rect 9232 15960 9260 16136
rect 12894 16124 12900 16136
rect 12952 16124 12958 16176
rect 9490 16056 9496 16108
rect 9548 16096 9554 16108
rect 9766 16096 9772 16108
rect 9548 16068 9772 16096
rect 9548 16056 9554 16068
rect 9766 16056 9772 16068
rect 9824 16096 9830 16108
rect 11333 16099 11391 16105
rect 11333 16096 11345 16099
rect 9824 16068 11345 16096
rect 9824 16056 9830 16068
rect 10923 16037 10951 16068
rect 11333 16065 11345 16068
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 10908 16031 10966 16037
rect 10908 15997 10920 16031
rect 10954 15997 10966 16031
rect 10908 15991 10966 15997
rect 12504 16031 12562 16037
rect 12504 15997 12516 16031
rect 12550 16028 12562 16031
rect 12802 16028 12808 16040
rect 12550 16000 12808 16028
rect 12550 15997 12562 16000
rect 12504 15991 12562 15997
rect 12802 15988 12808 16000
rect 12860 16028 12866 16040
rect 13265 16031 13323 16037
rect 13265 16028 13277 16031
rect 12860 16000 13277 16028
rect 12860 15988 12866 16000
rect 13265 15997 13277 16000
rect 13311 15997 13323 16031
rect 13265 15991 13323 15997
rect 9446 15963 9504 15969
rect 9446 15960 9458 15963
rect 9232 15932 9458 15960
rect 9446 15929 9458 15932
rect 9492 15960 9504 15963
rect 9950 15960 9956 15972
rect 9492 15932 9956 15960
rect 9492 15929 9504 15932
rect 9446 15923 9504 15929
rect 9950 15920 9956 15932
rect 10008 15920 10014 15972
rect 5626 15892 5632 15904
rect 4019 15864 5632 15892
rect 4019 15861 4031 15864
rect 3973 15855 4031 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 10045 15895 10103 15901
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10594 15892 10600 15904
rect 10091 15864 10600 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 4890 15688 4896 15700
rect 4847 15660 4896 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 4890 15648 4896 15660
rect 4948 15648 4954 15700
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 6178 15688 6184 15700
rect 5316 15660 6184 15688
rect 5316 15648 5322 15660
rect 5546 15629 5574 15660
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6822 15688 6828 15700
rect 6735 15660 6828 15688
rect 6822 15648 6828 15660
rect 6880 15688 6886 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6880 15660 7021 15688
rect 6880 15648 6886 15660
rect 7009 15657 7021 15660
rect 7055 15657 7067 15691
rect 7009 15651 7067 15657
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7892 15660 7941 15688
rect 7892 15648 7898 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 7929 15651 7987 15657
rect 8018 15648 8024 15700
rect 8076 15688 8082 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 8076 15660 8309 15688
rect 8076 15648 8082 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 8297 15651 8355 15657
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 10008 15660 10057 15688
rect 10008 15648 10014 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 10045 15651 10103 15657
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 10652 15660 11652 15688
rect 10652 15648 10658 15660
rect 5531 15623 5589 15629
rect 5531 15589 5543 15623
rect 5577 15589 5589 15623
rect 7852 15620 7880 15648
rect 5531 15583 5589 15589
rect 5644 15592 7880 15620
rect 5258 15512 5264 15564
rect 5316 15552 5322 15564
rect 5644 15552 5672 15592
rect 11238 15580 11244 15632
rect 11296 15620 11302 15632
rect 11624 15629 11652 15660
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 11296 15592 11529 15620
rect 11296 15580 11302 15592
rect 11517 15589 11529 15592
rect 11563 15589 11575 15623
rect 11517 15583 11575 15589
rect 11609 15623 11667 15629
rect 11609 15589 11621 15623
rect 11655 15620 11667 15623
rect 11698 15620 11704 15632
rect 11655 15592 11704 15620
rect 11655 15589 11667 15592
rect 11609 15583 11667 15589
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 5316 15524 5672 15552
rect 5316 15512 5322 15524
rect 6730 15512 6736 15564
rect 6788 15552 6794 15564
rect 6917 15555 6975 15561
rect 6917 15552 6929 15555
rect 6788 15524 6929 15552
rect 6788 15512 6794 15524
rect 6917 15521 6929 15524
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15552 7527 15555
rect 8018 15552 8024 15564
rect 7515 15524 8024 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8202 15512 8208 15564
rect 8260 15552 8266 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 8260 15524 8493 15552
rect 8260 15512 8266 15524
rect 8481 15521 8493 15524
rect 8527 15521 8539 15555
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 8481 15515 8539 15521
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 12986 15552 12992 15564
rect 12947 15524 12992 15552
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5810 15484 5816 15496
rect 5215 15456 5816 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 3050 15376 3056 15428
rect 3108 15416 3114 15428
rect 7834 15416 7840 15428
rect 3108 15388 7840 15416
rect 3108 15376 3114 15388
rect 7834 15376 7840 15388
rect 7892 15416 7898 15428
rect 8665 15419 8723 15425
rect 8665 15416 8677 15419
rect 7892 15388 8677 15416
rect 7892 15376 7898 15388
rect 8665 15385 8677 15388
rect 8711 15385 8723 15419
rect 12066 15416 12072 15428
rect 12027 15388 12072 15416
rect 8665 15379 8723 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 6086 15348 6092 15360
rect 6047 15320 6092 15348
rect 6086 15308 6092 15320
rect 6144 15308 6150 15360
rect 10594 15348 10600 15360
rect 10555 15320 10600 15348
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13127 15351 13185 15357
rect 13127 15348 13139 15351
rect 12768 15320 13139 15348
rect 12768 15308 12774 15320
rect 13127 15317 13139 15320
rect 13173 15317 13185 15351
rect 13127 15311 13185 15317
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 8018 15144 8024 15156
rect 7979 15116 8024 15144
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 8260 15116 8401 15144
rect 8260 15104 8266 15116
rect 8389 15113 8401 15116
rect 8435 15113 8447 15147
rect 8846 15144 8852 15156
rect 8807 15116 8852 15144
rect 8389 15107 8447 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10008 15116 10149 15144
rect 10008 15104 10014 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10594 15144 10600 15156
rect 10555 15116 10600 15144
rect 10137 15107 10195 15113
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 11698 15144 11704 15156
rect 11659 15116 11704 15144
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 3200 15048 4154 15076
rect 3200 15036 3206 15048
rect 4126 14940 4154 15048
rect 4890 15036 4896 15088
rect 4948 15076 4954 15088
rect 10870 15076 10876 15088
rect 4948 15048 10876 15076
rect 4948 15036 4954 15048
rect 10870 15036 10876 15048
rect 10928 15036 10934 15088
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 12986 15076 12992 15088
rect 11204 15048 12992 15076
rect 11204 15036 11210 15048
rect 12986 15036 12992 15048
rect 13044 15036 13050 15088
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4798 15008 4804 15020
rect 4571 14980 4804 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4798 14968 4804 14980
rect 4856 15008 4862 15020
rect 6822 15008 6828 15020
rect 4856 14980 5580 15008
rect 6783 14980 6828 15008
rect 4856 14968 4862 14980
rect 5552 14952 5580 14980
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 8938 15008 8944 15020
rect 8352 14980 8944 15008
rect 8352 14968 8358 14980
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 10962 15008 10968 15020
rect 10827 14980 10968 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 10962 14968 10968 14980
rect 11020 15008 11026 15020
rect 13587 15011 13645 15017
rect 13587 15008 13599 15011
rect 11020 14980 13599 15008
rect 11020 14968 11026 14980
rect 13587 14977 13599 14980
rect 13633 14977 13645 15011
rect 13587 14971 13645 14977
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4126 14912 4905 14940
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5258 14940 5264 14952
rect 4939 14912 5264 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5534 14940 5540 14952
rect 5447 14912 5540 14940
rect 5534 14900 5540 14912
rect 5592 14940 5598 14952
rect 8018 14940 8024 14952
rect 5592 14912 8024 14940
rect 5592 14900 5598 14912
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12504 14943 12562 14949
rect 12504 14940 12516 14943
rect 12299 14912 12516 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12504 14909 12516 14912
rect 12550 14940 12562 14943
rect 12894 14940 12900 14952
rect 12550 14912 12900 14940
rect 12550 14909 12562 14912
rect 12504 14903 12562 14909
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 13484 14943 13542 14949
rect 13484 14940 13496 14943
rect 13412 14912 13496 14940
rect 13412 14900 13418 14912
rect 13484 14909 13496 14912
rect 13530 14940 13542 14943
rect 13530 14909 13543 14940
rect 13484 14903 13543 14909
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14872 6147 14875
rect 6178 14872 6184 14884
rect 6135 14844 6184 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 6178 14832 6184 14844
rect 6236 14872 6242 14884
rect 6641 14875 6699 14881
rect 6641 14872 6653 14875
rect 6236 14844 6653 14872
rect 6236 14832 6242 14844
rect 6641 14841 6653 14844
rect 6687 14872 6699 14875
rect 7187 14875 7245 14881
rect 7187 14872 7199 14875
rect 6687 14844 7199 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7187 14841 7199 14844
rect 7233 14872 7245 14875
rect 7650 14872 7656 14884
rect 7233 14844 7656 14872
rect 7233 14841 7245 14844
rect 7187 14835 7245 14841
rect 7650 14832 7656 14844
rect 7708 14872 7714 14884
rect 8846 14872 8852 14884
rect 7708 14844 8852 14872
rect 7708 14832 7714 14844
rect 8846 14832 8852 14844
rect 8904 14872 8910 14884
rect 9262 14875 9320 14881
rect 9262 14872 9274 14875
rect 8904 14844 9274 14872
rect 8904 14832 8910 14844
rect 9262 14841 9274 14844
rect 9308 14841 9320 14875
rect 9262 14835 9320 14841
rect 10873 14875 10931 14881
rect 10873 14841 10885 14875
rect 10919 14841 10931 14875
rect 10873 14835 10931 14841
rect 5258 14804 5264 14816
rect 5219 14776 5264 14804
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 9858 14804 9864 14816
rect 9819 14776 9864 14804
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10888 14804 10916 14835
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11425 14875 11483 14881
rect 11425 14872 11437 14875
rect 11112 14844 11437 14872
rect 11112 14832 11118 14844
rect 11425 14841 11437 14844
rect 11471 14841 11483 14875
rect 11425 14835 11483 14841
rect 13515 14816 13543 14903
rect 10652 14776 10916 14804
rect 10652 14764 10658 14776
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12575 14807 12633 14813
rect 12575 14804 12587 14807
rect 12032 14776 12587 14804
rect 12032 14764 12038 14776
rect 12575 14773 12587 14776
rect 12621 14773 12633 14807
rect 13515 14804 13544 14816
rect 13451 14776 13544 14804
rect 12575 14767 12633 14773
rect 13538 14764 13544 14776
rect 13596 14804 13602 14816
rect 13909 14807 13967 14813
rect 13909 14804 13921 14807
rect 13596 14776 13921 14804
rect 13596 14764 13602 14776
rect 13909 14773 13921 14776
rect 13955 14773 13967 14807
rect 13909 14767 13967 14773
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 5316 14572 5457 14600
rect 5316 14560 5322 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5445 14563 5503 14569
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 6788 14572 7389 14600
rect 6788 14560 6794 14572
rect 7377 14569 7389 14572
rect 7423 14569 7435 14603
rect 7834 14600 7840 14612
rect 7795 14572 7840 14600
rect 7377 14563 7435 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 8018 14600 8024 14612
rect 7979 14572 8024 14600
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8938 14600 8944 14612
rect 8899 14572 8944 14600
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9732 14572 9965 14600
rect 9732 14560 9738 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 11296 14572 11437 14600
rect 11296 14560 11302 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11425 14563 11483 14569
rect 6549 14535 6607 14541
rect 6549 14501 6561 14535
rect 6595 14532 6607 14535
rect 6638 14532 6644 14544
rect 6595 14504 6644 14532
rect 6595 14501 6607 14504
rect 6549 14495 6607 14501
rect 6638 14492 6644 14504
rect 6696 14532 6702 14544
rect 7742 14532 7748 14544
rect 6696 14504 7748 14532
rect 6696 14492 6702 14504
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 7852 14532 7880 14560
rect 7852 14504 8432 14532
rect 4890 14464 4896 14476
rect 4851 14436 4896 14464
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 7926 14464 7932 14476
rect 7887 14436 7932 14464
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 8404 14473 8432 14504
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10505 14535 10563 14541
rect 10505 14532 10517 14535
rect 9916 14504 10517 14532
rect 9916 14492 9922 14504
rect 10505 14501 10517 14504
rect 10551 14532 10563 14535
rect 11146 14532 11152 14544
rect 10551 14504 11152 14532
rect 10551 14501 10563 14504
rect 10505 14495 10563 14501
rect 11146 14492 11152 14504
rect 11204 14532 11210 14544
rect 12069 14535 12127 14541
rect 12069 14532 12081 14535
rect 11204 14504 12081 14532
rect 11204 14492 11210 14504
rect 12069 14501 12081 14504
rect 12115 14501 12127 14535
rect 12069 14495 12127 14501
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 8846 14464 8852 14476
rect 8435 14436 8852 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 8846 14424 8852 14436
rect 8904 14424 8910 14476
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11112 14436 11157 14464
rect 11112 14424 11118 14436
rect 6178 14356 6184 14408
rect 6236 14396 6242 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6236 14368 6469 14396
rect 6236 14356 6242 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6730 14396 6736 14408
rect 6691 14368 6736 14396
rect 6457 14359 6515 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 11606 14396 11612 14408
rect 10459 14368 11612 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14396 12035 14399
rect 12710 14396 12716 14408
rect 12023 14368 12716 14396
rect 12023 14365 12035 14368
rect 11977 14359 12035 14365
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 8294 14288 8300 14340
rect 8352 14328 8358 14340
rect 10502 14328 10508 14340
rect 8352 14300 10508 14328
rect 8352 14288 8358 14300
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 10870 14288 10876 14340
rect 10928 14328 10934 14340
rect 12066 14328 12072 14340
rect 10928 14300 12072 14328
rect 10928 14288 10934 14300
rect 12066 14288 12072 14300
rect 12124 14328 12130 14340
rect 12529 14331 12587 14337
rect 12529 14328 12541 14331
rect 12124 14300 12541 14328
rect 12124 14288 12130 14300
rect 12529 14297 12541 14300
rect 12575 14297 12587 14331
rect 12529 14291 12587 14297
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 5123 14263 5181 14269
rect 5123 14260 5135 14263
rect 4396 14232 5135 14260
rect 4396 14220 4402 14232
rect 5123 14229 5135 14232
rect 5169 14229 5181 14263
rect 5123 14223 5181 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 3007 14059 3065 14065
rect 3007 14025 3019 14059
rect 3053 14056 3065 14059
rect 6178 14056 6184 14068
rect 3053 14028 6184 14056
rect 3053 14025 3065 14028
rect 3007 14019 3065 14025
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6273 14059 6331 14065
rect 6273 14025 6285 14059
rect 6319 14056 6331 14059
rect 6638 14056 6644 14068
rect 6319 14028 6644 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7926 14056 7932 14068
rect 7887 14028 7932 14056
rect 7926 14016 7932 14028
rect 7984 14056 7990 14068
rect 8110 14056 8116 14068
rect 7984 14028 8116 14056
rect 7984 14016 7990 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 10045 14059 10103 14065
rect 10045 14025 10057 14059
rect 10091 14056 10103 14059
rect 10594 14056 10600 14068
rect 10091 14028 10600 14056
rect 10091 14025 10103 14028
rect 10045 14019 10103 14025
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11606 14056 11612 14068
rect 11519 14028 11612 14056
rect 11606 14016 11612 14028
rect 11664 14056 11670 14068
rect 11974 14056 11980 14068
rect 11664 14028 11980 14056
rect 11664 14016 11670 14028
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12710 14056 12716 14068
rect 12671 14028 12716 14056
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 4019 13991 4077 13997
rect 4019 13957 4031 13991
rect 4065 13988 4077 13991
rect 11164 13988 11192 14016
rect 11885 13991 11943 13997
rect 11885 13988 11897 13991
rect 4065 13960 6960 13988
rect 11164 13960 11897 13988
rect 4065 13957 4077 13960
rect 4019 13951 4077 13957
rect 6932 13932 6960 13960
rect 11885 13957 11897 13960
rect 11931 13957 11943 13991
rect 11885 13951 11943 13957
rect 4430 13920 4436 13932
rect 4391 13892 4436 13920
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13920 4951 13923
rect 5258 13920 5264 13932
rect 4939 13892 5264 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 6914 13920 6920 13932
rect 6827 13892 6920 13920
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 10870 13920 10876 13932
rect 10831 13892 10876 13920
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 2936 13855 2994 13861
rect 2936 13821 2948 13855
rect 2982 13821 2994 13855
rect 2936 13815 2994 13821
rect 3948 13855 4006 13861
rect 3948 13821 3960 13855
rect 3994 13852 4006 13855
rect 4448 13852 4476 13880
rect 3994 13824 4476 13852
rect 3994 13821 4006 13824
rect 3948 13815 4006 13821
rect 2951 13716 2979 13815
rect 4448 13796 4476 13824
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8168 13824 8401 13852
rect 8168 13812 8174 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8389 13815 8447 13821
rect 8496 13824 8861 13852
rect 4430 13744 4436 13796
rect 4488 13744 4494 13796
rect 4801 13787 4859 13793
rect 4801 13753 4813 13787
rect 4847 13784 4859 13787
rect 4890 13784 4896 13796
rect 4847 13756 4896 13784
rect 4847 13753 4859 13756
rect 4801 13747 4859 13753
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 5626 13744 5632 13796
rect 5684 13784 5690 13796
rect 5684 13756 6316 13784
rect 5684 13744 5690 13756
rect 3418 13716 3424 13728
rect 2951 13688 3424 13716
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 5258 13716 5264 13728
rect 5219 13688 5264 13716
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 5813 13719 5871 13725
rect 5813 13716 5825 13719
rect 5408 13688 5825 13716
rect 5408 13676 5414 13688
rect 5813 13685 5825 13688
rect 5859 13685 5871 13719
rect 6288 13716 6316 13756
rect 6638 13744 6644 13796
rect 6696 13784 6702 13796
rect 7009 13787 7067 13793
rect 7009 13784 7021 13787
rect 6696 13756 7021 13784
rect 6696 13744 6702 13756
rect 7009 13753 7021 13756
rect 7055 13753 7067 13787
rect 7009 13747 7067 13753
rect 8496 13716 8524 13824
rect 8849 13821 8861 13824
rect 8895 13852 8907 13855
rect 9401 13855 9459 13861
rect 9401 13852 9413 13855
rect 8895 13824 9413 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 9401 13821 9413 13824
rect 9447 13821 9459 13855
rect 9401 13815 9459 13821
rect 10226 13784 10232 13796
rect 10187 13756 10232 13784
rect 10226 13744 10232 13756
rect 10284 13744 10290 13796
rect 10321 13787 10379 13793
rect 10321 13753 10333 13787
rect 10367 13784 10379 13787
rect 10594 13784 10600 13796
rect 10367 13756 10600 13784
rect 10367 13753 10379 13756
rect 10321 13747 10379 13753
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 8662 13716 8668 13728
rect 6288 13688 8524 13716
rect 8623 13688 8668 13716
rect 5813 13679 5871 13685
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 6086 13512 6092 13524
rect 5920 13484 6092 13512
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 4341 13447 4399 13453
rect 4341 13444 4353 13447
rect 4120 13416 4353 13444
rect 4120 13404 4126 13416
rect 4341 13413 4353 13416
rect 4387 13444 4399 13447
rect 5350 13444 5356 13456
rect 4387 13416 5356 13444
rect 4387 13413 4399 13416
rect 4341 13407 4399 13413
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 5920 13453 5948 13484
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 6733 13515 6791 13521
rect 6733 13512 6745 13515
rect 6236 13484 6745 13512
rect 6236 13472 6242 13484
rect 6733 13481 6745 13484
rect 6779 13481 6791 13515
rect 6733 13475 6791 13481
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7101 13515 7159 13521
rect 7101 13512 7113 13515
rect 6972 13484 7113 13512
rect 6972 13472 6978 13484
rect 7101 13481 7113 13484
rect 7147 13481 7159 13515
rect 7101 13475 7159 13481
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 8812 13484 9996 13512
rect 8812 13472 8818 13484
rect 5905 13447 5963 13453
rect 5905 13413 5917 13447
rect 5951 13413 5963 13447
rect 7926 13444 7932 13456
rect 7887 13416 7932 13444
rect 5905 13407 5963 13413
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 9858 13444 9864 13456
rect 9819 13416 9864 13444
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 9968 13444 9996 13484
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10284 13484 10701 13512
rect 10284 13472 10290 13484
rect 10689 13481 10701 13484
rect 10735 13512 10747 13515
rect 11379 13515 11437 13521
rect 11379 13512 11391 13515
rect 10735 13484 11391 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 11379 13481 11391 13484
rect 11425 13481 11437 13515
rect 11379 13475 11437 13481
rect 9968 13416 11351 13444
rect 11323 13385 11351 13416
rect 11308 13379 11366 13385
rect 11308 13345 11320 13379
rect 11354 13376 11366 13379
rect 11974 13376 11980 13388
rect 11354 13348 11980 13376
rect 11354 13345 11366 13348
rect 11308 13339 11366 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 4338 13308 4344 13320
rect 4295 13280 4344 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4890 13308 4896 13320
rect 4851 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 5166 13268 5172 13320
rect 5224 13308 5230 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5224 13280 5825 13308
rect 5224 13268 5230 13280
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 8662 13308 8668 13320
rect 7699 13280 8668 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 10870 13308 10876 13320
rect 9815 13280 10876 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 6362 13240 6368 13252
rect 6323 13212 6368 13240
rect 6362 13200 6368 13212
rect 6420 13200 6426 13252
rect 6638 13200 6644 13252
rect 6696 13240 6702 13252
rect 8110 13240 8116 13252
rect 6696 13212 8116 13240
rect 6696 13200 6702 13212
rect 8110 13200 8116 13212
rect 8168 13240 8174 13252
rect 8849 13243 8907 13249
rect 8849 13240 8861 13243
rect 8168 13212 8861 13240
rect 8168 13200 8174 13212
rect 8849 13209 8861 13212
rect 8895 13209 8907 13243
rect 8849 13203 8907 13209
rect 10321 13243 10379 13249
rect 10321 13209 10333 13243
rect 10367 13240 10379 13243
rect 10502 13240 10508 13252
rect 10367 13212 10508 13240
rect 10367 13209 10379 13212
rect 10321 13203 10379 13209
rect 10502 13200 10508 13212
rect 10560 13200 10566 13252
rect 5258 13172 5264 13184
rect 5171 13144 5264 13172
rect 5258 13132 5264 13144
rect 5316 13172 5322 13184
rect 7926 13172 7932 13184
rect 5316 13144 7932 13172
rect 5316 13132 5322 13144
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 8570 13172 8576 13184
rect 8531 13144 8576 13172
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 3697 12971 3755 12977
rect 3697 12937 3709 12971
rect 3743 12968 3755 12971
rect 4338 12968 4344 12980
rect 3743 12940 4344 12968
rect 3743 12937 3755 12940
rect 3697 12931 3755 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 6144 12940 6193 12968
rect 6144 12928 6150 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 7653 12971 7711 12977
rect 7653 12937 7665 12971
rect 7699 12968 7711 12971
rect 7926 12968 7932 12980
rect 7699 12940 7932 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 8941 12971 8999 12977
rect 8941 12968 8953 12971
rect 8720 12940 8953 12968
rect 8720 12928 8726 12940
rect 8941 12937 8953 12940
rect 8987 12937 8999 12971
rect 10870 12968 10876 12980
rect 10831 12940 10876 12968
rect 8941 12931 8999 12937
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 4062 12900 4068 12912
rect 4023 12872 4068 12900
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 5166 12860 5172 12912
rect 5224 12900 5230 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 5224 12872 6561 12900
rect 5224 12860 5230 12872
rect 6549 12869 6561 12872
rect 6595 12869 6607 12903
rect 9858 12900 9864 12912
rect 6549 12863 6607 12869
rect 8680 12872 9864 12900
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12832 7343 12835
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7331 12804 7757 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 7745 12801 7757 12804
rect 7791 12832 7803 12835
rect 8018 12832 8024 12844
rect 7791 12804 8024 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 4208 12767 4266 12773
rect 4208 12733 4220 12767
rect 4254 12764 4266 12767
rect 4706 12764 4712 12776
rect 4254 12736 4712 12764
rect 4254 12733 4266 12736
rect 4208 12727 4266 12733
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 4295 12699 4353 12705
rect 4295 12665 4307 12699
rect 4341 12696 4353 12699
rect 5258 12696 5264 12708
rect 4341 12668 5264 12696
rect 4341 12665 4353 12668
rect 4295 12659 4353 12665
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 5350 12656 5356 12708
rect 5408 12696 5414 12708
rect 5905 12699 5963 12705
rect 5408 12668 5453 12696
rect 5408 12656 5414 12668
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 6362 12696 6368 12708
rect 5951 12668 6368 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 6362 12656 6368 12668
rect 6420 12696 6426 12708
rect 7374 12696 7380 12708
rect 6420 12668 7380 12696
rect 6420 12656 6426 12668
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 7926 12656 7932 12708
rect 7984 12696 7990 12708
rect 8066 12699 8124 12705
rect 8066 12696 8078 12699
rect 7984 12668 8078 12696
rect 7984 12656 7990 12668
rect 8066 12665 8078 12668
rect 8112 12665 8124 12699
rect 8066 12659 8124 12665
rect 4706 12628 4712 12640
rect 4667 12600 4712 12628
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5077 12631 5135 12637
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 5368 12628 5396 12656
rect 5123 12600 5396 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 8680 12637 8708 12872
rect 9858 12860 9864 12872
rect 9916 12900 9922 12912
rect 10505 12903 10563 12909
rect 10505 12900 10517 12903
rect 9916 12872 10517 12900
rect 9916 12860 9922 12872
rect 10505 12869 10517 12872
rect 10551 12869 10563 12903
rect 10505 12863 10563 12869
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9674 12832 9680 12844
rect 9447 12804 9680 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 13446 12832 13452 12844
rect 9824 12804 13452 12832
rect 9824 12792 9830 12804
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 11124 12767 11182 12773
rect 11124 12733 11136 12767
rect 11170 12764 11182 12767
rect 11514 12764 11520 12776
rect 11170 12736 11520 12764
rect 11170 12733 11182 12736
rect 11124 12727 11182 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 9585 12699 9643 12705
rect 9585 12665 9597 12699
rect 9631 12665 9643 12699
rect 9585 12659 9643 12665
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 8260 12600 8677 12628
rect 8260 12588 8266 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 8665 12591 8723 12597
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 9600 12628 9628 12659
rect 9674 12656 9680 12708
rect 9732 12696 9738 12708
rect 10226 12696 10232 12708
rect 9732 12668 9777 12696
rect 10187 12668 10232 12696
rect 9732 12656 9738 12668
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 9548 12600 9628 12628
rect 11195 12631 11253 12637
rect 9548 12588 9554 12600
rect 11195 12597 11207 12631
rect 11241 12628 11253 12631
rect 11330 12628 11336 12640
rect 11241 12600 11336 12628
rect 11241 12597 11253 12600
rect 11195 12591 11253 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 11974 12628 11980 12640
rect 11887 12600 11980 12628
rect 11974 12588 11980 12600
rect 12032 12628 12038 12640
rect 12618 12628 12624 12640
rect 12032 12600 12624 12628
rect 12032 12588 12038 12600
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 5031 12427 5089 12433
rect 5031 12393 5043 12427
rect 5077 12424 5089 12427
rect 5166 12424 5172 12436
rect 5077 12396 5172 12424
rect 5077 12393 5089 12396
rect 5031 12387 5089 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5353 12427 5411 12433
rect 5353 12424 5365 12427
rect 5316 12396 5365 12424
rect 5316 12384 5322 12396
rect 5353 12393 5365 12396
rect 5399 12393 5411 12427
rect 5353 12387 5411 12393
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 7926 12424 7932 12436
rect 7883 12396 7932 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 9876 12396 11468 12424
rect 6086 12356 6092 12368
rect 6047 12328 6092 12356
rect 6086 12316 6092 12328
rect 6144 12316 6150 12368
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 8202 12356 8208 12368
rect 7340 12328 8208 12356
rect 7340 12316 7346 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 9582 12356 9588 12368
rect 8628 12328 9588 12356
rect 8628 12316 8634 12328
rect 9582 12316 9588 12328
rect 9640 12356 9646 12368
rect 9876 12365 9904 12396
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 9640 12328 9873 12356
rect 9640 12316 9646 12328
rect 9861 12325 9873 12328
rect 9907 12325 9919 12359
rect 11330 12356 11336 12368
rect 11291 12328 11336 12356
rect 9861 12319 9919 12325
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 11440 12365 11468 12396
rect 11425 12359 11483 12365
rect 11425 12325 11437 12359
rect 11471 12356 11483 12359
rect 11974 12356 11980 12368
rect 11471 12328 11980 12356
rect 11471 12325 11483 12328
rect 11425 12319 11483 12325
rect 11974 12316 11980 12328
rect 12032 12316 12038 12368
rect 12856 12291 12914 12297
rect 12856 12257 12868 12291
rect 12902 12288 12914 12291
rect 13262 12288 13268 12300
rect 12902 12260 13268 12288
rect 12902 12257 12914 12260
rect 12856 12251 12914 12257
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6086 12220 6092 12232
rect 6043 12192 6092 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12220 6331 12223
rect 6730 12220 6736 12232
rect 6319 12192 6736 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 4890 12112 4896 12164
rect 4948 12152 4954 12164
rect 6288 12152 6316 12183
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 8110 12220 8116 12232
rect 8071 12192 8116 12220
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 9766 12220 9772 12232
rect 9679 12192 9772 12220
rect 9766 12180 9772 12192
rect 9824 12220 9830 12232
rect 12943 12223 13001 12229
rect 12943 12220 12955 12223
rect 9824 12192 12955 12220
rect 9824 12180 9830 12192
rect 12943 12189 12955 12192
rect 12989 12189 13001 12223
rect 12943 12183 13001 12189
rect 4948 12124 6316 12152
rect 8665 12155 8723 12161
rect 4948 12112 4954 12124
rect 8665 12121 8677 12155
rect 8711 12152 8723 12155
rect 10226 12152 10232 12164
rect 8711 12124 10232 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 10226 12112 10232 12124
rect 10284 12152 10290 12164
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 10284 12124 10333 12152
rect 10284 12112 10290 12124
rect 10321 12121 10333 12124
rect 10367 12121 10379 12155
rect 10321 12115 10379 12121
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 11885 12155 11943 12161
rect 11885 12152 11897 12155
rect 10560 12124 11897 12152
rect 10560 12112 10566 12124
rect 11885 12121 11897 12124
rect 11931 12121 11943 12155
rect 11885 12115 11943 12121
rect 4801 12087 4859 12093
rect 4801 12053 4813 12087
rect 4847 12084 4859 12087
rect 4982 12084 4988 12096
rect 4847 12056 4988 12084
rect 4847 12053 4859 12056
rect 4801 12047 4859 12053
rect 4982 12044 4988 12056
rect 5040 12084 5046 12096
rect 5442 12084 5448 12096
rect 5040 12056 5448 12084
rect 5040 12044 5046 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 4893 11883 4951 11889
rect 4893 11849 4905 11883
rect 4939 11880 4951 11883
rect 5534 11880 5540 11892
rect 4939 11852 5540 11880
rect 4939 11849 4951 11852
rect 4893 11843 4951 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 5902 11880 5908 11892
rect 5675 11852 5908 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 5644 11676 5672 11843
rect 5902 11840 5908 11852
rect 5960 11840 5966 11892
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6236 11852 6561 11880
rect 6236 11840 6242 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 6549 11843 6607 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7653 11883 7711 11889
rect 7653 11849 7665 11883
rect 7699 11880 7711 11883
rect 7926 11880 7932 11892
rect 7699 11852 7932 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 8662 11880 8668 11892
rect 8575 11852 8668 11880
rect 8662 11840 8668 11852
rect 8720 11880 8726 11892
rect 9674 11880 9680 11892
rect 8720 11852 9680 11880
rect 8720 11840 8726 11852
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 11149 11883 11207 11889
rect 11149 11849 11161 11883
rect 11195 11880 11207 11883
rect 11330 11880 11336 11892
rect 11195 11852 11336 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 12032 11852 12081 11880
rect 12032 11840 12038 11852
rect 12069 11849 12081 11852
rect 12115 11849 12127 11883
rect 12986 11880 12992 11892
rect 12947 11852 12992 11880
rect 12069 11843 12127 11849
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 9582 11812 9588 11824
rect 9543 11784 9588 11812
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 13262 11812 13268 11824
rect 13223 11784 13268 11812
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 6270 11744 6276 11756
rect 5803 11716 6276 11744
rect 5803 11688 5831 11716
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9180 11716 9781 11744
rect 9180 11704 9186 11716
rect 9769 11713 9781 11716
rect 9815 11744 9827 11747
rect 10502 11744 10508 11756
rect 9815 11716 10508 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11379 11747 11437 11753
rect 11379 11744 11391 11747
rect 10928 11716 11391 11744
rect 10928 11704 10934 11716
rect 11379 11713 11391 11716
rect 11425 11713 11437 11747
rect 11379 11707 11437 11713
rect 5803 11685 5816 11688
rect 5788 11679 5816 11685
rect 5788 11676 5800 11679
rect 4755 11648 5672 11676
rect 5723 11648 5800 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 5788 11645 5800 11648
rect 5788 11639 5816 11645
rect 5810 11636 5816 11639
rect 5868 11636 5874 11688
rect 7742 11676 7748 11688
rect 7703 11648 7748 11676
rect 7742 11636 7748 11648
rect 7800 11676 7806 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 7800 11648 8953 11676
rect 7800 11636 7806 11648
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 11276 11679 11334 11685
rect 11276 11676 11288 11679
rect 11204 11648 11288 11676
rect 11204 11636 11210 11648
rect 11276 11645 11288 11648
rect 11322 11676 11334 11679
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11322 11648 11713 11676
rect 11322 11645 11334 11648
rect 11276 11639 11334 11645
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 12504 11679 12562 11685
rect 12504 11676 12516 11679
rect 12216 11648 12516 11676
rect 12216 11636 12222 11648
rect 12504 11645 12516 11648
rect 12550 11676 12562 11679
rect 12986 11676 12992 11688
rect 12550 11648 12992 11676
rect 12550 11645 12562 11648
rect 12504 11639 12562 11645
rect 12986 11636 12992 11648
rect 13044 11636 13050 11688
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 5261 11611 5319 11617
rect 5261 11608 5273 11611
rect 5040 11580 5273 11608
rect 5040 11568 5046 11580
rect 5261 11577 5273 11580
rect 5307 11608 5319 11611
rect 7282 11608 7288 11620
rect 5307 11580 7288 11608
rect 5307 11577 5319 11580
rect 5261 11571 5319 11577
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8066 11611 8124 11617
rect 8066 11608 8078 11611
rect 7984 11580 8078 11608
rect 7984 11568 7990 11580
rect 8066 11577 8078 11580
rect 8112 11577 8124 11611
rect 8066 11571 8124 11577
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 9861 11611 9919 11617
rect 9364 11580 9720 11608
rect 9364 11568 9370 11580
rect 5859 11543 5917 11549
rect 5859 11509 5871 11543
rect 5905 11540 5917 11543
rect 6086 11540 6092 11552
rect 5905 11512 6092 11540
rect 5905 11509 5917 11512
rect 5859 11503 5917 11509
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9398 11540 9404 11552
rect 8904 11512 9404 11540
rect 8904 11500 8910 11512
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9692 11540 9720 11580
rect 9861 11577 9873 11611
rect 9907 11577 9919 11611
rect 10410 11608 10416 11620
rect 10371 11580 10416 11608
rect 9861 11571 9919 11577
rect 9876 11540 9904 11571
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 9692 11512 10701 11540
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 10689 11503 10747 11509
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 12575 11543 12633 11549
rect 12575 11540 12587 11543
rect 10836 11512 12587 11540
rect 10836 11500 10842 11512
rect 12575 11509 12587 11512
rect 12621 11509 12633 11543
rect 12575 11503 12633 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 5718 11336 5724 11348
rect 5679 11308 5724 11336
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 6086 11336 6092 11348
rect 6047 11308 6092 11336
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 6788 11308 7297 11336
rect 6788 11296 6794 11308
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 7285 11299 7343 11305
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9122 11336 9128 11348
rect 8904 11308 9128 11336
rect 8904 11296 8910 11308
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 9766 11336 9772 11348
rect 9539 11308 9772 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 11379 11339 11437 11345
rect 11379 11305 11391 11339
rect 11425 11336 11437 11339
rect 12066 11336 12072 11348
rect 11425 11308 12072 11336
rect 11425 11305 11437 11308
rect 11379 11299 11437 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 7009 11271 7067 11277
rect 4724 11240 6592 11268
rect 4724 11209 4752 11240
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11169 4767 11203
rect 4709 11163 4767 11169
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4724 11132 4752 11163
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 4856 11172 5273 11200
rect 4856 11160 4862 11172
rect 5261 11169 5273 11172
rect 5307 11200 5319 11203
rect 5902 11200 5908 11212
rect 5307 11172 5908 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 6564 11209 6592 11240
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 7742 11268 7748 11280
rect 7055 11240 7748 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 8158 11271 8216 11277
rect 8158 11268 8170 11271
rect 7984 11240 8170 11268
rect 7984 11228 7990 11240
rect 8158 11237 8170 11240
rect 8204 11237 8216 11271
rect 9858 11268 9864 11280
rect 9819 11240 9864 11268
rect 8158 11231 8216 11237
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 6638 11200 6644 11212
rect 6595 11172 6644 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 6822 11200 6828 11212
rect 6783 11172 6828 11200
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 10428 11200 10456 11228
rect 11276 11203 11334 11209
rect 11276 11200 11288 11203
rect 10428 11172 11288 11200
rect 11276 11169 11288 11172
rect 11322 11169 11334 11203
rect 11276 11163 11334 11169
rect 12320 11203 12378 11209
rect 12320 11169 12332 11203
rect 12366 11200 12378 11203
rect 12618 11200 12624 11212
rect 12366 11172 12624 11200
rect 12366 11169 12378 11172
rect 12320 11163 12378 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 4120 11104 4752 11132
rect 5445 11135 5503 11141
rect 4120 11092 4126 11104
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 5491 11104 7849 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 7837 11101 7849 11104
rect 7883 11132 7895 11135
rect 8202 11132 8208 11144
rect 7883 11104 8208 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 10226 11132 10232 11144
rect 9815 11104 10232 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10226 11092 10232 11104
rect 10284 11132 10290 11144
rect 11422 11132 11428 11144
rect 10284 11104 11428 11132
rect 10284 11092 10290 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 7745 11067 7803 11073
rect 7745 11033 7757 11067
rect 7791 11064 7803 11067
rect 8110 11064 8116 11076
rect 7791 11036 8116 11064
rect 7791 11033 7803 11036
rect 7745 11027 7803 11033
rect 8110 11024 8116 11036
rect 8168 11064 8174 11076
rect 12391 11067 12449 11073
rect 12391 11064 12403 11067
rect 8168 11036 12403 11064
rect 8168 11024 8174 11036
rect 12391 11033 12403 11036
rect 12437 11033 12449 11067
rect 12391 11027 12449 11033
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 4062 10792 4068 10804
rect 4023 10764 4068 10792
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 7926 10792 7932 10804
rect 7887 10764 7932 10792
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 8812 10764 9505 10792
rect 8812 10752 8818 10764
rect 9493 10761 9505 10764
rect 9539 10792 9551 10795
rect 9858 10792 9864 10804
rect 9539 10764 9864 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 11422 10792 11428 10804
rect 11383 10764 11428 10792
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 10778 10724 10784 10736
rect 8588 10696 10784 10724
rect 8588 10668 8616 10696
rect 10778 10684 10784 10696
rect 10836 10684 10842 10736
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 4396 10628 5549 10656
rect 4396 10616 4402 10628
rect 5537 10625 5549 10628
rect 5583 10656 5595 10659
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 5583 10628 7205 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 7193 10625 7205 10628
rect 7239 10656 7251 10659
rect 7650 10656 7656 10668
rect 7239 10628 7656 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 8570 10656 8576 10668
rect 8483 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8846 10656 8852 10668
rect 8807 10628 8852 10656
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 10410 10656 10416 10668
rect 10371 10628 10416 10656
rect 10410 10616 10416 10628
rect 10468 10656 10474 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 10468 10628 11805 10656
rect 10468 10616 10474 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 5258 10520 5264 10532
rect 4203 10492 5264 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5353 10523 5411 10529
rect 5353 10489 5365 10523
rect 5399 10520 5411 10523
rect 5718 10520 5724 10532
rect 5399 10492 5724 10520
rect 5399 10489 5411 10492
rect 5353 10483 5411 10489
rect 5718 10480 5724 10492
rect 5776 10480 5782 10532
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 6917 10523 6975 10529
rect 6917 10520 6929 10523
rect 6788 10492 6929 10520
rect 6788 10480 6794 10492
rect 6917 10489 6929 10492
rect 6963 10489 6975 10523
rect 6917 10483 6975 10489
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7064 10492 7109 10520
rect 7064 10480 7070 10492
rect 8662 10480 8668 10532
rect 8720 10520 8726 10532
rect 9953 10523 10011 10529
rect 8720 10492 8765 10520
rect 8720 10480 8726 10492
rect 9953 10489 9965 10523
rect 9999 10520 10011 10523
rect 10134 10520 10140 10532
rect 9999 10492 10140 10520
rect 9999 10489 10011 10492
rect 9953 10483 10011 10489
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 10229 10523 10287 10529
rect 10229 10489 10241 10523
rect 10275 10489 10287 10523
rect 10229 10483 10287 10489
rect 6365 10455 6423 10461
rect 6365 10421 6377 10455
rect 6411 10452 6423 10455
rect 6638 10452 6644 10464
rect 6411 10424 6644 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8680 10452 8708 10480
rect 8435 10424 8708 10452
rect 10244 10452 10272 10483
rect 10594 10452 10600 10464
rect 10244 10424 10600 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 10594 10412 10600 10424
rect 10652 10452 10658 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 10652 10424 11069 10452
rect 10652 10412 10658 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 12618 10452 12624 10464
rect 12579 10424 12624 10452
rect 11057 10415 11115 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 5258 10248 5264 10260
rect 5219 10220 5264 10248
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 6822 10248 6828 10260
rect 5408 10220 6828 10248
rect 5408 10208 5414 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 7984 10220 8109 10248
rect 7984 10208 7990 10220
rect 5902 10189 5908 10192
rect 5899 10180 5908 10189
rect 5863 10152 5908 10180
rect 5899 10143 5908 10152
rect 5902 10140 5908 10143
rect 5960 10140 5966 10192
rect 7466 10180 7472 10192
rect 7427 10152 7472 10180
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 8081 10180 8109 10220
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 8260 10220 8309 10248
rect 8260 10208 8266 10220
rect 8297 10217 8309 10220
rect 8343 10217 8355 10251
rect 8297 10211 8355 10217
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8628 10220 8677 10248
rect 8628 10208 8634 10220
rect 8665 10217 8677 10220
rect 8711 10217 8723 10251
rect 10594 10248 10600 10260
rect 10555 10220 10600 10248
rect 8665 10211 8723 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 9766 10180 9772 10192
rect 8081 10152 9772 10180
rect 9766 10140 9772 10152
rect 9824 10180 9830 10192
rect 9998 10183 10056 10189
rect 9998 10180 10010 10183
rect 9824 10152 10010 10180
rect 9824 10140 9830 10152
rect 9998 10149 10010 10152
rect 10044 10149 10056 10183
rect 9998 10143 10056 10149
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 10192 10152 11437 10180
rect 10192 10140 10198 10152
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 11425 10143 11483 10149
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 4522 10112 4528 10124
rect 3568 10084 4528 10112
rect 3568 10072 3574 10084
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 7006 10112 7012 10124
rect 6503 10084 7012 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 7006 10072 7012 10084
rect 7064 10112 7070 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 7064 10084 7113 10112
rect 7064 10072 7070 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 6914 10044 6920 10056
rect 5583 10016 6920 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7374 10044 7380 10056
rect 7287 10016 7380 10044
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7650 10044 7656 10056
rect 7611 10016 7656 10044
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 4430 9936 4436 9988
rect 4488 9976 4494 9988
rect 6822 9976 6828 9988
rect 4488 9948 6828 9976
rect 4488 9936 4494 9948
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 7392 9976 7420 10004
rect 9033 9979 9091 9985
rect 9033 9976 9045 9979
rect 7392 9948 9045 9976
rect 9033 9945 9045 9948
rect 9079 9945 9091 9979
rect 9033 9939 9091 9945
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 4522 9704 4528 9716
rect 4483 9676 4528 9704
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 9766 9704 9772 9716
rect 6696 9676 8984 9704
rect 9727 9676 9772 9704
rect 6696 9664 6702 9676
rect 5905 9639 5963 9645
rect 5905 9605 5917 9639
rect 5951 9636 5963 9639
rect 7466 9636 7472 9648
rect 5951 9608 7472 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 7466 9596 7472 9608
rect 7524 9636 7530 9648
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7524 9608 7849 9636
rect 7524 9596 7530 9608
rect 7837 9605 7849 9608
rect 7883 9605 7895 9639
rect 7837 9599 7895 9605
rect 7558 9568 7564 9580
rect 7116 9540 7564 9568
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 4203 9472 4997 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4985 9469 4997 9472
rect 5031 9500 5043 9503
rect 5442 9500 5448 9512
rect 5031 9472 5448 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7116 9509 7144 9540
rect 7558 9528 7564 9540
rect 7616 9568 7622 9580
rect 7616 9540 8432 9568
rect 7616 9528 7622 9540
rect 8404 9512 8432 9540
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 7064 9472 7113 9500
rect 7064 9460 7070 9472
rect 7101 9469 7113 9472
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 8386 9500 8392 9512
rect 8299 9472 8392 9500
rect 7285 9463 7343 9469
rect 4893 9435 4951 9441
rect 4893 9401 4905 9435
rect 4939 9432 4951 9435
rect 5347 9435 5405 9441
rect 5347 9432 5359 9435
rect 4939 9404 5359 9432
rect 4939 9401 4951 9404
rect 4893 9395 4951 9401
rect 5347 9401 5359 9404
rect 5393 9401 5405 9435
rect 5347 9395 5405 9401
rect 5368 9364 5396 9395
rect 6086 9392 6092 9444
rect 6144 9432 6150 9444
rect 6549 9435 6607 9441
rect 6549 9432 6561 9435
rect 6144 9404 6561 9432
rect 6144 9392 6150 9404
rect 6549 9401 6561 9404
rect 6595 9432 6607 9435
rect 7300 9432 7328 9463
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8846 9500 8852 9512
rect 8807 9472 8852 9500
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 8956 9500 8984 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9732 9540 10701 9568
rect 9732 9528 9738 9540
rect 10689 9537 10701 9540
rect 10735 9568 10747 9571
rect 11333 9571 11391 9577
rect 11333 9568 11345 9571
rect 10735 9540 11345 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 11333 9537 11345 9540
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 10229 9503 10287 9509
rect 10229 9500 10241 9503
rect 8956 9472 10241 9500
rect 10229 9469 10241 9472
rect 10275 9469 10287 9503
rect 10410 9500 10416 9512
rect 10371 9472 10416 9500
rect 10229 9463 10287 9469
rect 6595 9404 7328 9432
rect 8297 9435 8355 9441
rect 6595 9401 6607 9404
rect 6549 9395 6607 9401
rect 8297 9401 8309 9435
rect 8343 9432 8355 9435
rect 8864 9432 8892 9460
rect 8343 9404 8892 9432
rect 9125 9435 9183 9441
rect 8343 9401 8355 9404
rect 8297 9395 8355 9401
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 9582 9432 9588 9444
rect 9171 9404 9588 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 9582 9392 9588 9404
rect 9640 9392 9646 9444
rect 10244 9432 10272 9463
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10244 9404 10977 9432
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 5902 9364 5908 9376
rect 5368 9336 5908 9364
rect 5902 9324 5908 9336
rect 5960 9364 5966 9376
rect 6273 9367 6331 9373
rect 6273 9364 6285 9367
rect 5960 9336 6285 9364
rect 5960 9324 5966 9336
rect 6273 9333 6285 9336
rect 6319 9364 6331 9367
rect 6638 9364 6644 9376
rect 6319 9336 6644 9364
rect 6319 9333 6331 9336
rect 6273 9327 6331 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 6914 9364 6920 9376
rect 6875 9336 6920 9364
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 4764 9132 5181 9160
rect 4764 9120 4770 9132
rect 5169 9129 5181 9132
rect 5215 9160 5227 9163
rect 5258 9160 5264 9172
rect 5215 9132 5264 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 5442 9160 5448 9172
rect 5403 9132 5448 9160
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6457 9163 6515 9169
rect 6457 9129 6469 9163
rect 6503 9160 6515 9163
rect 6914 9160 6920 9172
rect 6503 9132 6920 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7156 9132 8753 9160
rect 7156 9120 7162 9132
rect 6638 9052 6644 9104
rect 6696 9092 6702 9104
rect 7463 9095 7521 9101
rect 7463 9092 7475 9095
rect 6696 9064 7475 9092
rect 6696 9052 6702 9064
rect 7463 9061 7475 9064
rect 7509 9092 7521 9095
rect 7926 9092 7932 9104
rect 7509 9064 7932 9092
rect 7509 9061 7521 9064
rect 7463 9055 7521 9061
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 8386 9092 8392 9104
rect 8347 9064 8392 9092
rect 8386 9052 8392 9064
rect 8444 9052 8450 9104
rect 8725 9092 8753 9132
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 9815 9163 9873 9169
rect 9815 9160 9827 9163
rect 9548 9132 9827 9160
rect 9548 9120 9554 9132
rect 9815 9129 9827 9132
rect 9861 9129 9873 9163
rect 9815 9123 9873 9129
rect 8725 9064 10732 9092
rect 4338 9024 4344 9036
rect 4299 8996 4344 9024
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 5534 9024 5540 9036
rect 5495 8996 5540 9024
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 6086 9024 6092 9036
rect 5859 8996 6092 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 5828 8956 5856 8987
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7006 9024 7012 9036
rect 6963 8996 7012 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9674 9024 9680 9036
rect 9732 9033 9738 9036
rect 10704 9033 10732 9064
rect 9732 9027 9770 9033
rect 8536 8996 9680 9024
rect 8536 8984 8542 8996
rect 9674 8984 9680 8996
rect 9758 8993 9770 9027
rect 9732 8987 9770 8993
rect 10689 9027 10747 9033
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 10778 9024 10784 9036
rect 10735 8996 10784 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 9732 8984 9738 8987
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 7098 8956 7104 8968
rect 4948 8928 5856 8956
rect 7059 8928 7104 8956
rect 4948 8916 4954 8928
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 8202 8956 8208 8968
rect 7248 8928 8208 8956
rect 7248 8916 7254 8928
rect 8202 8916 8208 8928
rect 8260 8956 8266 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8260 8928 8769 8956
rect 8260 8916 8266 8928
rect 8757 8925 8769 8928
rect 8803 8956 8815 8959
rect 10410 8956 10416 8968
rect 8803 8928 10416 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 10410 8916 10416 8928
rect 10468 8956 10474 8968
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 10468 8928 10517 8956
rect 10468 8916 10474 8928
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 7208 8888 7236 8916
rect 10226 8888 10232 8900
rect 5224 8860 7236 8888
rect 10139 8860 10232 8888
rect 5224 8848 5230 8860
rect 10226 8848 10232 8860
rect 10284 8888 10290 8900
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 10284 8860 10885 8888
rect 10284 8848 10290 8860
rect 10873 8857 10885 8860
rect 10919 8857 10931 8891
rect 10873 8851 10931 8857
rect 106 8780 112 8832
rect 164 8820 170 8832
rect 4479 8823 4537 8829
rect 4479 8820 4491 8823
rect 164 8792 4491 8820
rect 164 8780 170 8792
rect 4479 8789 4491 8792
rect 4525 8789 4537 8823
rect 8018 8820 8024 8832
rect 7979 8792 8024 8820
rect 4479 8783 4537 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4338 8616 4344 8628
rect 4299 8588 4344 8616
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 4856 8588 4997 8616
rect 4856 8576 4862 8588
rect 4985 8585 4997 8588
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 4709 8551 4767 8557
rect 4709 8517 4721 8551
rect 4755 8548 4767 8551
rect 4890 8548 4896 8560
rect 4755 8520 4896 8548
rect 4755 8517 4767 8520
rect 4709 8511 4767 8517
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 5000 8412 5028 8579
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 5592 8588 6193 8616
rect 5592 8576 5598 8588
rect 6181 8585 6193 8588
rect 6227 8616 6239 8619
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 6227 8588 9229 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 9217 8585 9229 8588
rect 9263 8616 9275 8619
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9263 8588 9505 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9674 8616 9680 8628
rect 9635 8588 9680 8616
rect 9493 8579 9551 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10778 8616 10784 8628
rect 10739 8588 10784 8616
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 7745 8551 7803 8557
rect 7745 8517 7757 8551
rect 7791 8548 7803 8551
rect 7926 8548 7932 8560
rect 7791 8520 7932 8548
rect 7791 8517 7803 8520
rect 7745 8511 7803 8517
rect 7926 8508 7932 8520
rect 7984 8508 7990 8560
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 5951 8452 7021 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7009 8449 7021 8452
rect 7055 8480 7067 8483
rect 7098 8480 7104 8492
rect 7055 8452 7104 8480
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8846 8480 8852 8492
rect 8159 8452 8852 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5000 8384 5181 8412
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5316 8384 5641 8412
rect 5316 8372 5322 8384
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 8202 8412 8208 8424
rect 8163 8384 8208 8412
rect 5629 8375 5687 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 8772 8421 8800 8452
rect 8846 8440 8852 8452
rect 8904 8480 8910 8492
rect 9306 8480 9312 8492
rect 8904 8452 9312 8480
rect 8904 8440 8910 8452
rect 9306 8440 9312 8452
rect 9364 8480 9370 8492
rect 9364 8452 10272 8480
rect 9364 8440 9370 8452
rect 10244 8424 10272 8452
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 9539 8384 9781 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 10226 8412 10232 8424
rect 10187 8384 10232 8412
rect 9769 8375 9827 8381
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 8904 8316 8953 8344
rect 8904 8304 8910 8316
rect 8941 8313 8953 8316
rect 8987 8313 8999 8347
rect 8941 8307 8999 8313
rect 7190 8276 7196 8288
rect 7151 8248 7196 8276
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 7006 8072 7012 8084
rect 5874 8044 7012 8072
rect 5874 8004 5902 8044
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 5092 7976 5902 8004
rect 6549 8007 6607 8013
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 5092 7945 5120 7976
rect 6549 7973 6561 8007
rect 6595 8004 6607 8007
rect 6730 8004 6736 8016
rect 6595 7976 6736 8004
rect 6595 7973 6607 7976
rect 6549 7967 6607 7973
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 8110 8004 8116 8016
rect 8071 7976 8116 8004
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 9766 7964 9772 8016
rect 9824 8004 9830 8016
rect 9998 8007 10056 8013
rect 9998 8004 10010 8007
rect 9824 7976 10010 8004
rect 9824 7964 9830 7976
rect 9998 7973 10010 7976
rect 10044 7973 10056 8007
rect 9998 7967 10056 7973
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4580 7908 5089 7936
rect 4580 7896 4586 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5258 7936 5264 7948
rect 5219 7908 5264 7936
rect 5077 7899 5135 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9640 7908 9689 7936
rect 9640 7896 9646 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 5534 7868 5540 7880
rect 5495 7840 5540 7868
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6196 7840 6469 7868
rect 5810 7692 5816 7744
rect 5868 7732 5874 7744
rect 6196 7741 6224 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 7098 7868 7104 7880
rect 7059 7840 7104 7868
rect 6457 7831 6515 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7616 7840 8033 7868
rect 7616 7828 7622 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 8754 7868 8760 7880
rect 8711 7840 8760 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 10376 7840 11437 7868
rect 10376 7828 10382 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 5868 7704 6193 7732
rect 5868 7692 5874 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 10594 7732 10600 7744
rect 10555 7704 10600 7732
rect 6181 7695 6239 7701
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 4522 7528 4528 7540
rect 4483 7500 4528 7528
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5258 7528 5264 7540
rect 4939 7500 5264 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 7745 7531 7803 7537
rect 7745 7497 7757 7531
rect 7791 7528 7803 7531
rect 8110 7528 8116 7540
rect 7791 7500 8116 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 10781 7531 10839 7537
rect 10781 7528 10793 7531
rect 9640 7500 10793 7528
rect 9640 7488 9646 7500
rect 10781 7497 10793 7500
rect 10827 7497 10839 7531
rect 10781 7491 10839 7497
rect 9125 7463 9183 7469
rect 9125 7429 9137 7463
rect 9171 7460 9183 7463
rect 9766 7460 9772 7472
rect 9171 7432 9772 7460
rect 9171 7429 9183 7432
rect 9125 7423 9183 7429
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 11103 7463 11161 7469
rect 11103 7429 11115 7463
rect 11149 7460 11161 7463
rect 12342 7460 12348 7472
rect 11149 7432 12348 7460
rect 11149 7429 11161 7432
rect 11103 7423 11161 7429
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 5592 7364 6837 7392
rect 5592 7352 5598 7364
rect 6825 7361 6837 7364
rect 6871 7392 6883 7395
rect 7006 7392 7012 7404
rect 6871 7364 7012 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 8846 7352 8852 7404
rect 8904 7392 8910 7404
rect 9214 7392 9220 7404
rect 8904 7364 9220 7392
rect 8904 7352 8910 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 5166 7324 5172 7336
rect 5127 7296 5172 7324
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5316 7296 5641 7324
rect 5316 7284 5322 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 11000 7327 11058 7333
rect 11000 7324 11012 7327
rect 8812 7296 11012 7324
rect 8812 7284 8818 7296
rect 11000 7293 11012 7296
rect 11046 7324 11058 7327
rect 11425 7327 11483 7333
rect 11425 7324 11437 7327
rect 11046 7296 11437 7324
rect 11046 7293 11058 7296
rect 11000 7287 11058 7293
rect 11425 7293 11437 7296
rect 11471 7293 11483 7327
rect 11425 7287 11483 7293
rect 5902 7256 5908 7268
rect 5863 7228 5908 7256
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 6273 7259 6331 7265
rect 6273 7225 6285 7259
rect 6319 7256 6331 7259
rect 6730 7256 6736 7268
rect 6319 7228 6736 7256
rect 6319 7225 6331 7228
rect 6273 7219 6331 7225
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 7187 7259 7245 7265
rect 7187 7225 7199 7259
rect 7233 7256 7245 7259
rect 8110 7256 8116 7268
rect 7233 7228 8116 7256
rect 7233 7225 7245 7228
rect 7187 7219 7245 7225
rect 6638 7188 6644 7200
rect 6551 7160 6644 7188
rect 6638 7148 6644 7160
rect 6696 7188 6702 7200
rect 7202 7188 7230 7219
rect 8110 7216 8116 7228
rect 8168 7256 8174 7268
rect 9579 7259 9637 7265
rect 9579 7256 9591 7259
rect 8168 7228 9591 7256
rect 8168 7216 8174 7228
rect 9579 7225 9591 7228
rect 9625 7256 9637 7259
rect 9766 7256 9772 7268
rect 9625 7228 9772 7256
rect 9625 7225 9637 7228
rect 9579 7219 9637 7225
rect 9766 7216 9772 7228
rect 9824 7256 9830 7268
rect 10413 7259 10471 7265
rect 10413 7256 10425 7259
rect 9824 7228 10425 7256
rect 9824 7216 9830 7228
rect 10413 7225 10425 7228
rect 10459 7225 10471 7259
rect 10413 7219 10471 7225
rect 6696 7160 7230 7188
rect 6696 7148 6702 7160
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 7616 7160 8401 7188
rect 7616 7148 7622 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 10134 7188 10140 7200
rect 10095 7160 10140 7188
rect 8389 7151 8447 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 4939 6987 4997 6993
rect 4939 6953 4951 6987
rect 4985 6984 4997 6987
rect 5810 6984 5816 6996
rect 4985 6956 5816 6984
rect 4985 6953 4997 6956
rect 4939 6947 4997 6953
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 5960 6956 7573 6984
rect 5960 6944 5966 6956
rect 7561 6953 7573 6956
rect 7607 6984 7619 6987
rect 8110 6984 8116 6996
rect 7607 6956 7788 6984
rect 8071 6956 8116 6984
rect 7607 6953 7619 6956
rect 7561 6947 7619 6953
rect 5258 6916 5264 6928
rect 5219 6888 5264 6916
rect 5258 6876 5264 6888
rect 5316 6876 5322 6928
rect 6175 6919 6233 6925
rect 6175 6885 6187 6919
rect 6221 6916 6233 6919
rect 6638 6916 6644 6928
rect 6221 6888 6644 6916
rect 6221 6885 6233 6888
rect 6175 6879 6233 6885
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 7006 6916 7012 6928
rect 6967 6888 7012 6916
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4836 6851 4894 6857
rect 4836 6848 4848 6851
rect 4672 6820 4848 6848
rect 4672 6808 4678 6820
rect 4836 6817 4848 6820
rect 4882 6817 4894 6851
rect 4836 6811 4894 6817
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 7760 6857 7788 6956
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 9214 6984 9220 6996
rect 9175 6956 9220 6984
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 10597 6987 10655 6993
rect 10597 6953 10609 6987
rect 10643 6984 10655 6987
rect 11422 6984 11428 6996
rect 10643 6956 11428 6984
rect 10643 6953 10655 6956
rect 10597 6947 10655 6953
rect 11422 6944 11428 6956
rect 11480 6984 11486 6996
rect 11480 6956 11652 6984
rect 11480 6944 11486 6956
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9998 6919 10056 6925
rect 9998 6916 10010 6919
rect 9824 6888 10010 6916
rect 9824 6876 9830 6888
rect 9998 6885 10010 6888
rect 10044 6885 10056 6919
rect 9998 6879 10056 6885
rect 10134 6876 10140 6928
rect 10192 6916 10198 6928
rect 10410 6916 10416 6928
rect 10192 6888 10416 6916
rect 10192 6876 10198 6888
rect 10410 6876 10416 6888
rect 10468 6916 10474 6928
rect 11624 6925 11652 6956
rect 10873 6919 10931 6925
rect 10873 6916 10885 6919
rect 10468 6888 10885 6916
rect 10468 6876 10474 6888
rect 10873 6885 10885 6888
rect 10919 6885 10931 6919
rect 10873 6879 10931 6885
rect 11609 6919 11667 6925
rect 11609 6885 11621 6919
rect 11655 6885 11667 6919
rect 11609 6879 11667 6885
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 5224 6820 5641 6848
rect 5224 6808 5230 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9858 6848 9864 6860
rect 9723 6820 9864 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6086 6780 6092 6792
rect 5859 6752 6092 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 11514 6780 11520 6792
rect 11475 6752 11520 6780
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 6730 6644 6736 6656
rect 6643 6616 6736 6644
rect 6730 6604 6736 6616
rect 6788 6644 6794 6656
rect 7006 6644 7012 6656
rect 6788 6616 7012 6644
rect 6788 6604 6794 6616
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 8665 6647 8723 6653
rect 8665 6613 8677 6647
rect 8711 6644 8723 6647
rect 8754 6644 8760 6656
rect 8711 6616 8760 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 4798 6440 4804 6452
rect 4672 6412 4804 6440
rect 4672 6400 4678 6412
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 7248 6412 8401 6440
rect 7248 6400 7254 6412
rect 8389 6409 8401 6412
rect 8435 6409 8447 6443
rect 9766 6440 9772 6452
rect 9727 6412 9772 6440
rect 8389 6403 8447 6409
rect 6641 6375 6699 6381
rect 6641 6341 6653 6375
rect 6687 6372 6699 6375
rect 7929 6375 7987 6381
rect 7929 6372 7941 6375
rect 6687 6344 7941 6372
rect 6687 6341 6699 6344
rect 6641 6335 6699 6341
rect 7929 6341 7941 6344
rect 7975 6372 7987 6375
rect 8110 6372 8116 6384
rect 7975 6344 8116 6372
rect 7975 6341 7987 6344
rect 7929 6335 7987 6341
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 8404 6304 8432 6403
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 11422 6440 11428 6452
rect 11383 6412 11428 6440
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8404 6276 8677 6304
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8938 6304 8944 6316
rect 8899 6276 8944 6304
rect 8665 6267 8723 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10318 6304 10324 6316
rect 10183 6276 10324 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 5772 6239 5830 6245
rect 5772 6236 5784 6239
rect 3384 6208 5784 6236
rect 3384 6196 3390 6208
rect 5772 6205 5784 6208
rect 5818 6236 5830 6239
rect 6178 6236 6184 6248
rect 5818 6208 6184 6236
rect 5818 6205 5830 6208
rect 5772 6199 5830 6205
rect 6178 6196 6184 6208
rect 6236 6196 6242 6248
rect 5859 6171 5917 6177
rect 5859 6137 5871 6171
rect 5905 6168 5917 6171
rect 6914 6168 6920 6180
rect 5905 6140 6920 6168
rect 5905 6137 5917 6140
rect 5859 6131 5917 6137
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7558 6168 7564 6180
rect 7064 6140 7109 6168
rect 7519 6140 7564 6168
rect 7064 6128 7070 6140
rect 7558 6128 7564 6140
rect 7616 6128 7622 6180
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 8812 6140 8857 6168
rect 8812 6128 8818 6140
rect 10410 6128 10416 6180
rect 10468 6168 10474 6180
rect 10962 6168 10968 6180
rect 10468 6140 10513 6168
rect 10923 6140 10968 6168
rect 10468 6128 10474 6140
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 6086 6100 6092 6112
rect 5675 6072 6092 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6236 6072 6281 6100
rect 6236 6060 6242 6072
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11514 6100 11520 6112
rect 11112 6072 11520 6100
rect 11112 6060 11118 6072
rect 11514 6060 11520 6072
rect 11572 6100 11578 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11572 6072 11805 6100
rect 11572 6060 11578 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 6972 5868 7389 5896
rect 6972 5856 6978 5868
rect 7377 5865 7389 5868
rect 7423 5865 7435 5899
rect 8754 5896 8760 5908
rect 8715 5868 8760 5896
rect 7377 5859 7435 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9858 5896 9864 5908
rect 9819 5868 9864 5896
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 7006 5828 7012 5840
rect 5316 5800 6500 5828
rect 6967 5800 7012 5828
rect 5316 5788 5322 5800
rect 5626 5720 5632 5772
rect 5684 5760 5690 5772
rect 6472 5769 6500 5800
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 7098 5788 7104 5840
rect 7156 5828 7162 5840
rect 7745 5831 7803 5837
rect 7745 5828 7757 5831
rect 7156 5800 7757 5828
rect 7156 5788 7162 5800
rect 7745 5797 7757 5800
rect 7791 5797 7803 5831
rect 7745 5791 7803 5797
rect 7837 5831 7895 5837
rect 7837 5797 7849 5831
rect 7883 5828 7895 5831
rect 8018 5828 8024 5840
rect 7883 5800 8024 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 8938 5828 8944 5840
rect 8435 5800 8944 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 10229 5831 10287 5837
rect 10229 5797 10241 5831
rect 10275 5828 10287 5831
rect 10594 5828 10600 5840
rect 10275 5800 10600 5828
rect 10275 5797 10287 5800
rect 10229 5791 10287 5797
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5684 5732 6009 5760
rect 5684 5720 5690 5732
rect 5997 5729 6009 5732
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6546 5760 6552 5772
rect 6503 5732 6552 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 10962 5760 10968 5772
rect 10827 5732 10968 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 10962 5720 10968 5732
rect 11020 5760 11026 5772
rect 11676 5763 11734 5769
rect 11676 5760 11688 5763
rect 11020 5732 11688 5760
rect 11020 5720 11026 5732
rect 11676 5729 11688 5732
rect 11722 5760 11734 5763
rect 11974 5760 11980 5772
rect 11722 5732 11980 5760
rect 11722 5729 11734 5732
rect 11676 5723 11734 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 11747 5559 11805 5565
rect 11747 5525 11759 5559
rect 11793 5556 11805 5559
rect 13630 5556 13636 5568
rect 11793 5528 13636 5556
rect 11793 5525 11805 5528
rect 11747 5519 11805 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 5626 5352 5632 5364
rect 5587 5324 5632 5352
rect 5626 5312 5632 5324
rect 5684 5352 5690 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5684 5324 6377 5352
rect 5684 5312 5690 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6546 5352 6552 5364
rect 6507 5324 6552 5352
rect 6365 5315 6423 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7193 5355 7251 5361
rect 7193 5321 7205 5355
rect 7239 5352 7251 5355
rect 8018 5352 8024 5364
rect 7239 5324 8024 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9306 5352 9312 5364
rect 9171 5324 9312 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 6273 5287 6331 5293
rect 6273 5284 6285 5287
rect 5787 5256 6285 5284
rect 5787 5157 5815 5256
rect 6273 5253 6285 5256
rect 6319 5284 6331 5287
rect 6822 5284 6828 5296
rect 6319 5256 6828 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 7282 5244 7288 5296
rect 7340 5284 7346 5296
rect 8481 5287 8539 5293
rect 8481 5284 8493 5287
rect 7340 5256 8493 5284
rect 7340 5244 7346 5256
rect 8481 5253 8493 5256
rect 8527 5253 8539 5287
rect 8481 5247 8539 5253
rect 5859 5219 5917 5225
rect 5859 5185 5871 5219
rect 5905 5216 5917 5219
rect 8846 5216 8852 5228
rect 5905 5188 8852 5216
rect 5905 5185 5917 5188
rect 5859 5179 5917 5185
rect 8846 5176 8852 5188
rect 8904 5176 8910 5228
rect 9140 5216 9168 5315
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 10134 5312 10140 5364
rect 10192 5352 10198 5364
rect 10597 5355 10655 5361
rect 10597 5352 10609 5355
rect 10192 5324 10609 5352
rect 10192 5312 10198 5324
rect 10597 5321 10609 5324
rect 10643 5321 10655 5355
rect 10597 5315 10655 5321
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 11974 5352 11980 5364
rect 11747 5324 11980 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 12584 5324 12909 5352
rect 12584 5312 12590 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 10321 5219 10379 5225
rect 9140 5188 9720 5216
rect 5772 5151 5830 5157
rect 5772 5117 5784 5151
rect 5818 5117 5830 5151
rect 5772 5111 5830 5117
rect 6365 5151 6423 5157
rect 6365 5117 6377 5151
rect 6411 5148 6423 5151
rect 7650 5148 7656 5160
rect 6411 5120 7656 5148
rect 6411 5117 6423 5120
rect 6365 5111 6423 5117
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8570 5148 8576 5160
rect 8251 5120 8576 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 7561 5083 7619 5089
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 8220 5080 8248 5111
rect 8570 5108 8576 5120
rect 8628 5148 8634 5160
rect 9140 5148 9168 5188
rect 9398 5148 9404 5160
rect 8628 5120 9168 5148
rect 9359 5120 9404 5148
rect 8628 5108 8634 5120
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 9692 5157 9720 5188
rect 10321 5185 10333 5219
rect 10367 5216 10379 5219
rect 10594 5216 10600 5228
rect 10367 5188 10600 5216
rect 10367 5185 10379 5188
rect 10321 5179 10379 5185
rect 10594 5176 10600 5188
rect 10652 5176 10658 5228
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5117 9735 5151
rect 9677 5111 9735 5117
rect 10848 5151 10906 5157
rect 10848 5117 10860 5151
rect 10894 5117 10906 5151
rect 10848 5111 10906 5117
rect 8386 5080 8392 5092
rect 7607 5052 8248 5080
rect 8347 5052 8392 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 8481 5083 8539 5089
rect 8481 5049 8493 5083
rect 8527 5080 8539 5083
rect 10863 5080 10891 5111
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 12544 5157 12572 5312
rect 12488 5151 12572 5157
rect 12488 5148 12500 5151
rect 11388 5120 12500 5148
rect 11388 5108 11394 5120
rect 12488 5117 12500 5120
rect 12534 5120 12572 5151
rect 12534 5117 12546 5120
rect 12488 5111 12546 5117
rect 8527 5052 11376 5080
rect 8527 5049 8539 5052
rect 8481 5043 8539 5049
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8665 5015 8723 5021
rect 8665 5012 8677 5015
rect 7800 4984 8677 5012
rect 7800 4972 7806 4984
rect 8665 4981 8677 4984
rect 8711 4981 8723 5015
rect 9306 5012 9312 5024
rect 9267 4984 9312 5012
rect 8665 4975 8723 4981
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 10919 5015 10977 5021
rect 10919 4981 10931 5015
rect 10965 5012 10977 5015
rect 11146 5012 11152 5024
rect 10965 4984 11152 5012
rect 10965 4981 10977 4984
rect 10919 4975 10977 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11348 5021 11376 5052
rect 11514 5040 11520 5092
rect 11572 5080 11578 5092
rect 12575 5083 12633 5089
rect 12575 5080 12587 5083
rect 11572 5052 12587 5080
rect 11572 5040 11578 5052
rect 12575 5049 12587 5052
rect 12621 5049 12633 5083
rect 12575 5043 12633 5049
rect 11333 5015 11391 5021
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 13354 5012 13360 5024
rect 11379 4984 13360 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5224 4780 5273 4808
rect 5224 4768 5230 4780
rect 5261 4777 5273 4780
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4808 5414 4820
rect 7650 4808 7656 4820
rect 5408 4780 7230 4808
rect 7611 4780 7656 4808
rect 5408 4768 5414 4780
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 6641 4743 6699 4749
rect 6641 4740 6653 4743
rect 6236 4712 6653 4740
rect 6236 4700 6242 4712
rect 6641 4709 6653 4712
rect 6687 4709 6699 4743
rect 6641 4703 6699 4709
rect 5496 4675 5554 4681
rect 5496 4641 5508 4675
rect 5542 4672 5554 4675
rect 5902 4672 5908 4684
rect 5542 4644 5908 4672
rect 5542 4641 5554 4644
rect 5496 4635 5554 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 7202 4672 7230 4780
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 7892 4780 9321 4808
rect 7892 4768 7898 4780
rect 9309 4777 9321 4780
rect 9355 4808 9367 4811
rect 9398 4808 9404 4820
rect 9355 4780 9404 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 9732 4780 10041 4808
rect 9732 4768 9738 4780
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9824 4712 9873 4740
rect 9824 4700 9830 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 10013 4740 10041 4780
rect 10013 4712 12388 4740
rect 9861 4703 9919 4709
rect 12360 4684 12388 4712
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7202 4644 8033 4672
rect 8021 4641 8033 4644
rect 8067 4672 8079 4675
rect 8110 4672 8116 4684
rect 8067 4644 8116 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 11241 4675 11299 4681
rect 11241 4641 11253 4675
rect 11287 4672 11299 4675
rect 11330 4672 11336 4684
rect 11287 4644 11336 4672
rect 11287 4641 11299 4644
rect 11241 4635 11299 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 12342 4672 12348 4684
rect 12255 4644 12348 4672
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 13446 4672 13452 4684
rect 13407 4644 13452 4672
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 5583 4607 5641 4613
rect 5583 4573 5595 4607
rect 5629 4604 5641 4607
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5629 4576 6009 4604
rect 5629 4573 5641 4576
rect 5583 4567 5641 4573
rect 5997 4573 6009 4576
rect 6043 4604 6055 4607
rect 6549 4607 6607 4613
rect 6549 4604 6561 4607
rect 6043 4576 6561 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6549 4573 6561 4576
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 9398 4604 9404 4616
rect 8803 4576 9404 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 10134 4604 10140 4616
rect 9815 4576 10041 4604
rect 10095 4576 10140 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 7098 4536 7104 4548
rect 7059 4508 7104 4536
rect 7098 4496 7104 4508
rect 7156 4536 7162 4548
rect 7742 4536 7748 4548
rect 7156 4508 7748 4536
rect 7156 4496 7162 4508
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 10013 4536 10041 4576
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10689 4539 10747 4545
rect 10689 4536 10701 4539
rect 10013 4508 10701 4536
rect 10689 4505 10701 4508
rect 10735 4536 10747 4539
rect 10778 4536 10784 4548
rect 10735 4508 10784 4536
rect 10735 4505 10747 4508
rect 10689 4499 10747 4505
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 12529 4539 12587 4545
rect 12529 4505 12541 4539
rect 12575 4536 12587 4539
rect 13906 4536 13912 4548
rect 12575 4508 13912 4536
rect 12575 4505 12587 4508
rect 12529 4499 12587 4505
rect 13906 4496 13912 4508
rect 13964 4496 13970 4548
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 6273 4471 6331 4477
rect 6273 4468 6285 4471
rect 6236 4440 6285 4468
rect 6236 4428 6242 4440
rect 6273 4437 6285 4440
rect 6319 4437 6331 4471
rect 6273 4431 6331 4437
rect 11425 4471 11483 4477
rect 11425 4437 11437 4471
rect 11471 4468 11483 4471
rect 12250 4468 12256 4480
rect 11471 4440 12256 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 14182 4468 14188 4480
rect 13679 4440 14188 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 5077 4267 5135 4273
rect 5077 4233 5089 4267
rect 5123 4264 5135 4267
rect 5258 4264 5264 4276
rect 5123 4236 5264 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5258 4224 5264 4236
rect 5316 4224 5322 4276
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6270 4264 6276 4276
rect 6052 4236 6276 4264
rect 6052 4224 6058 4236
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 7929 4267 7987 4273
rect 7929 4233 7941 4267
rect 7975 4264 7987 4267
rect 8570 4264 8576 4276
rect 7975 4236 8576 4264
rect 7975 4233 7987 4236
rect 7929 4227 7987 4233
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 11330 4264 11336 4276
rect 11291 4236 11336 4264
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12342 4264 12348 4276
rect 12299 4236 12348 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 13446 4264 13452 4276
rect 13407 4236 13452 4264
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 4614 4196 4620 4208
rect 4575 4168 4620 4196
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 8168 4168 9597 4196
rect 8168 4156 8174 4168
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 9585 4159 9643 4165
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 9953 4199 10011 4205
rect 9953 4196 9965 4199
rect 9824 4168 9965 4196
rect 9824 4156 9830 4168
rect 9953 4165 9965 4168
rect 9999 4165 10011 4199
rect 9953 4159 10011 4165
rect 10410 4156 10416 4208
rect 10468 4196 10474 4208
rect 10781 4199 10839 4205
rect 10781 4196 10793 4199
rect 10468 4168 10793 4196
rect 10468 4156 10474 4168
rect 10781 4165 10793 4168
rect 10827 4196 10839 4199
rect 11054 4196 11060 4208
rect 10827 4168 11060 4196
rect 10827 4165 10839 4168
rect 10781 4159 10839 4165
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 6270 4128 6276 4140
rect 6231 4100 6276 4128
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 6696 4100 7205 4128
rect 6696 4088 6702 4100
rect 7193 4097 7205 4100
rect 7239 4128 7251 4131
rect 7558 4128 7564 4140
rect 7239 4100 7564 4128
rect 7239 4097 7251 4100
rect 7193 4091 7251 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 8202 4088 8208 4100
rect 8260 4128 8266 4140
rect 8260 4100 8753 4128
rect 8260 4088 8266 4100
rect 4224 4063 4282 4069
rect 4224 4029 4236 4063
rect 4270 4060 4282 4063
rect 4614 4060 4620 4072
rect 4270 4032 4620 4060
rect 4270 4029 4282 4032
rect 4224 4023 4282 4029
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 5166 4060 5172 4072
rect 5127 4032 5172 4060
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5316 4032 5641 4060
rect 5316 4020 5322 4032
rect 5629 4029 5641 4032
rect 5675 4029 5687 4063
rect 8386 4060 8392 4072
rect 8347 4032 8392 4060
rect 5629 4023 5687 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 5905 3995 5963 4001
rect 5905 3961 5917 3995
rect 5951 3992 5963 3995
rect 5994 3992 6000 4004
rect 5951 3964 6000 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 6914 3992 6920 4004
rect 6875 3964 6920 3992
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 8725 4001 8753 4100
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 10229 4131 10287 4137
rect 10229 4128 10241 4131
rect 8904 4100 10241 4128
rect 8904 4088 8910 4100
rect 10229 4097 10241 4100
rect 10275 4128 10287 4131
rect 11609 4131 11667 4137
rect 11609 4128 11621 4131
rect 10275 4100 11621 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 11609 4097 11621 4100
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 11238 4060 11244 4072
rect 10928 4032 11244 4060
rect 10928 4020 10934 4032
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 11756 4032 12449 4060
rect 11756 4020 11762 4032
rect 12437 4029 12449 4032
rect 12483 4060 12495 4063
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12483 4032 13001 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13608 4063 13666 4069
rect 13608 4029 13620 4063
rect 13654 4060 13666 4063
rect 13814 4060 13820 4072
rect 13654 4032 13820 4060
rect 13654 4029 13666 4032
rect 13608 4023 13666 4029
rect 13814 4020 13820 4032
rect 13872 4060 13878 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13872 4032 14013 4060
rect 13872 4020 13878 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3961 7067 3995
rect 7009 3955 7067 3961
rect 8710 3995 8768 4001
rect 8710 3961 8722 3995
rect 8756 3961 8768 3995
rect 8710 3955 8768 3961
rect 10321 3995 10379 4001
rect 10321 3961 10333 3995
rect 10367 3961 10379 3995
rect 10321 3955 10379 3961
rect 4295 3927 4353 3933
rect 4295 3893 4307 3927
rect 4341 3924 4353 3927
rect 6086 3924 6092 3936
rect 4341 3896 6092 3924
rect 4341 3893 4353 3896
rect 4295 3887 4353 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 6730 3924 6736 3936
rect 6687 3896 6736 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 6730 3884 6736 3896
rect 6788 3924 6794 3936
rect 7024 3924 7052 3955
rect 6788 3896 7052 3924
rect 9309 3927 9367 3933
rect 6788 3884 6794 3896
rect 9309 3893 9321 3927
rect 9355 3924 9367 3927
rect 9582 3924 9588 3936
rect 9355 3896 9588 3924
rect 9355 3893 9367 3896
rect 9309 3887 9367 3893
rect 9582 3884 9588 3896
rect 9640 3924 9646 3936
rect 10336 3924 10364 3955
rect 10686 3924 10692 3936
rect 9640 3896 10692 3924
rect 9640 3884 9646 3896
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 12710 3924 12716 3936
rect 12667 3896 12716 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13679 3927 13737 3933
rect 13679 3924 13691 3927
rect 13136 3896 13691 3924
rect 13136 3884 13142 3896
rect 13679 3893 13691 3896
rect 13725 3893 13737 3927
rect 13679 3887 13737 3893
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 7834 3720 7840 3732
rect 4632 3692 7840 3720
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4632 3593 4660 3692
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8444 3692 9045 3720
rect 8444 3680 8450 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 9033 3683 9091 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 10560 3692 11161 3720
rect 10560 3680 10566 3692
rect 11149 3689 11161 3692
rect 11195 3720 11207 3723
rect 11514 3720 11520 3732
rect 11195 3692 11520 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 5258 3652 5264 3664
rect 5000 3624 5264 3652
rect 5000 3596 5028 3624
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 6270 3661 6276 3664
rect 6267 3652 6276 3661
rect 6183 3624 6276 3652
rect 6267 3615 6276 3624
rect 6328 3652 6334 3664
rect 8202 3661 8208 3664
rect 8158 3655 8208 3661
rect 8158 3652 8170 3655
rect 6328 3624 8170 3652
rect 6270 3612 6276 3615
rect 6328 3612 6334 3624
rect 8158 3621 8170 3624
rect 8204 3621 8208 3655
rect 8158 3615 8208 3621
rect 8202 3612 8208 3615
rect 8260 3612 8266 3664
rect 9858 3652 9864 3664
rect 9771 3624 9864 3652
rect 9858 3612 9864 3624
rect 9916 3652 9922 3664
rect 11422 3652 11428 3664
rect 9916 3624 11428 3652
rect 9916 3612 9922 3624
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4120 3556 4629 3584
rect 4120 3544 4126 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 4893 3587 4951 3593
rect 4893 3553 4905 3587
rect 4939 3584 4951 3587
rect 4982 3584 4988 3596
rect 4939 3556 4988 3584
rect 4939 3553 4951 3556
rect 4893 3547 4951 3553
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3584 5135 3587
rect 6822 3584 6828 3596
rect 5123 3556 6828 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 6822 3544 6828 3556
rect 6880 3584 6886 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6880 3556 7113 3584
rect 6880 3544 6886 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3584 7895 3587
rect 8018 3584 8024 3596
rect 7883 3556 8024 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 8018 3544 8024 3556
rect 8076 3584 8082 3596
rect 9306 3584 9312 3596
rect 8076 3556 9312 3584
rect 8076 3544 8082 3556
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 13449 3587 13507 3593
rect 13449 3584 13461 3587
rect 13412 3556 13461 3584
rect 13412 3544 13418 3556
rect 13449 3553 13461 3556
rect 13495 3553 13507 3587
rect 13449 3547 13507 3553
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 5994 3516 6000 3528
rect 5951 3488 6000 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 10410 3516 10416 3528
rect 9815 3488 10272 3516
rect 10371 3488 10416 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 5350 3408 5356 3460
rect 5408 3448 5414 3460
rect 5445 3451 5503 3457
rect 5445 3448 5457 3451
rect 5408 3420 5457 3448
rect 5408 3408 5414 3420
rect 5445 3417 5457 3420
rect 5491 3448 5503 3451
rect 6178 3448 6184 3460
rect 5491 3420 6184 3448
rect 5491 3417 5503 3420
rect 5445 3411 5503 3417
rect 6178 3408 6184 3420
rect 6236 3448 6242 3460
rect 6825 3451 6883 3457
rect 6825 3448 6837 3451
rect 6236 3420 6837 3448
rect 6236 3408 6242 3420
rect 6825 3417 6837 3420
rect 6871 3417 6883 3451
rect 6825 3411 6883 3417
rect 5718 3380 5724 3392
rect 5679 3352 5724 3380
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 6914 3380 6920 3392
rect 6604 3352 6920 3380
rect 6604 3340 6610 3352
rect 6914 3340 6920 3352
rect 6972 3380 6978 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 6972 3352 7481 3380
rect 6972 3340 6978 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 8757 3383 8815 3389
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 9766 3380 9772 3392
rect 8803 3352 9772 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 9766 3340 9772 3352
rect 9824 3380 9830 3392
rect 10134 3380 10140 3392
rect 9824 3352 10140 3380
rect 9824 3340 9830 3352
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10244 3380 10272 3488
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11790 3516 11796 3528
rect 11379 3488 11796 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11790 3476 11796 3488
rect 11848 3516 11854 3528
rect 13078 3516 13084 3528
rect 11848 3488 13084 3516
rect 11848 3476 11854 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 10318 3408 10324 3460
rect 10376 3448 10382 3460
rect 11238 3448 11244 3460
rect 10376 3420 11244 3448
rect 10376 3408 10382 3420
rect 11238 3408 11244 3420
rect 11296 3448 11302 3460
rect 11885 3451 11943 3457
rect 11885 3448 11897 3451
rect 11296 3420 11897 3448
rect 11296 3408 11302 3420
rect 11885 3417 11897 3420
rect 11931 3417 11943 3451
rect 11885 3411 11943 3417
rect 11146 3380 11152 3392
rect 10244 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 15562 3380 15568 3392
rect 13679 3352 15568 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 4062 3176 4068 3188
rect 4023 3148 4068 3176
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4982 3176 4988 3188
rect 4943 3148 4988 3176
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3176 6334 3188
rect 6641 3179 6699 3185
rect 6641 3176 6653 3179
rect 6328 3148 6653 3176
rect 6328 3136 6334 3148
rect 6641 3145 6653 3148
rect 6687 3145 6699 3179
rect 6641 3139 6699 3145
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8202 3176 8208 3188
rect 8159 3148 8208 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8202 3136 8208 3148
rect 8260 3176 8266 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 8260 3148 8401 3176
rect 8260 3136 8266 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 9493 3179 9551 3185
rect 9493 3145 9505 3179
rect 9539 3176 9551 3179
rect 9858 3176 9864 3188
rect 9539 3148 9864 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10134 3176 10140 3188
rect 10095 3148 10140 3176
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12986 3176 12992 3188
rect 12947 3148 12992 3176
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13354 3176 13360 3188
rect 13315 3148 13360 3176
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 658 3068 664 3120
rect 716 3108 722 3120
rect 4295 3111 4353 3117
rect 716 3080 4154 3108
rect 716 3068 722 3080
rect 3212 2975 3270 2981
rect 3212 2941 3224 2975
rect 3258 2972 3270 2975
rect 4126 2972 4154 3080
rect 4295 3077 4307 3111
rect 4341 3108 4353 3111
rect 6546 3108 6552 3120
rect 4341 3080 6552 3108
rect 4341 3077 4353 3080
rect 4295 3071 4353 3077
rect 6546 3068 6552 3080
rect 6604 3068 6610 3120
rect 6730 3068 6736 3120
rect 6788 3108 6794 3120
rect 7745 3111 7803 3117
rect 7745 3108 7757 3111
rect 6788 3080 7757 3108
rect 6788 3068 6794 3080
rect 7745 3077 7757 3080
rect 7791 3077 7803 3111
rect 7745 3071 7803 3077
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 11149 3111 11207 3117
rect 11149 3108 11161 3111
rect 8352 3080 11161 3108
rect 8352 3068 8358 3080
rect 11149 3077 11161 3080
rect 11195 3077 11207 3111
rect 11149 3071 11207 3077
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 11572 3080 12633 3108
rect 11572 3068 11578 3080
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 12621 3071 12679 3077
rect 4522 3000 4528 3052
rect 4580 3040 4586 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 4580 3012 5273 3040
rect 4580 3000 4586 3012
rect 5261 3009 5273 3012
rect 5307 3040 5319 3043
rect 5718 3040 5724 3052
rect 5307 3012 5724 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 6638 3040 6644 3052
rect 5951 3012 6644 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 9398 3040 9404 3052
rect 8619 3012 9404 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10468 3012 10701 3040
rect 10468 3000 10474 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 13679 3043 13737 3049
rect 13679 3040 13691 3043
rect 10836 3012 13691 3040
rect 10836 3000 10842 3012
rect 13679 3009 13691 3012
rect 13725 3009 13737 3043
rect 13679 3003 13737 3009
rect 4224 2975 4282 2981
rect 4224 2972 4236 2975
rect 3258 2944 3740 2972
rect 4126 2944 4236 2972
rect 3258 2941 3270 2944
rect 3212 2935 3270 2941
rect 3712 2913 3740 2944
rect 4224 2941 4236 2944
rect 4270 2972 4282 2975
rect 12437 2975 12495 2981
rect 4270 2944 4752 2972
rect 4270 2941 4282 2944
rect 4224 2935 4282 2941
rect 3697 2907 3755 2913
rect 3697 2873 3709 2907
rect 3743 2904 3755 2907
rect 4614 2904 4620 2916
rect 3743 2876 4620 2904
rect 3743 2873 3755 2876
rect 3697 2867 3755 2873
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 3283 2839 3341 2845
rect 3283 2805 3295 2839
rect 3329 2836 3341 2839
rect 3510 2836 3516 2848
rect 3329 2808 3516 2836
rect 3329 2805 3341 2808
rect 3283 2799 3341 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 4724 2845 4752 2944
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12986 2972 12992 2984
rect 12483 2944 12992 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12986 2932 12992 2944
rect 13044 2932 13050 2984
rect 13592 2975 13650 2981
rect 13592 2972 13604 2975
rect 13096 2944 13604 2972
rect 5350 2904 5356 2916
rect 5311 2876 5356 2904
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 7187 2907 7245 2913
rect 7187 2873 7199 2907
rect 7233 2904 7245 2907
rect 8202 2904 8208 2916
rect 7233 2876 8208 2904
rect 7233 2873 7245 2876
rect 7187 2867 7245 2873
rect 8202 2864 8208 2876
rect 8260 2904 8266 2916
rect 8894 2907 8952 2913
rect 8894 2904 8906 2907
rect 8260 2876 8906 2904
rect 8260 2864 8266 2876
rect 8894 2873 8906 2876
rect 8940 2873 8952 2907
rect 10410 2904 10416 2916
rect 10371 2876 10416 2904
rect 8894 2867 8952 2873
rect 10410 2864 10416 2876
rect 10468 2864 10474 2916
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2873 10563 2907
rect 10505 2867 10563 2873
rect 11149 2907 11207 2913
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 13096 2904 13124 2944
rect 13592 2941 13604 2944
rect 13638 2972 13650 2975
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13638 2944 14013 2972
rect 13638 2941 13650 2944
rect 13592 2935 13650 2941
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 11195 2876 13124 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 8294 2836 8300 2848
rect 4755 2808 8300 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10520 2836 10548 2867
rect 10192 2808 10548 2836
rect 10192 2796 10198 2808
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 4522 2632 4528 2644
rect 4483 2604 4528 2632
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 6052 2604 6285 2632
rect 6052 2592 6058 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 6730 2632 6736 2644
rect 6691 2604 6736 2632
rect 6273 2595 6331 2601
rect 6730 2592 6736 2604
rect 6788 2632 6794 2644
rect 8018 2632 8024 2644
rect 6788 2604 7236 2632
rect 7979 2604 8024 2632
rect 6788 2592 6794 2604
rect 3510 2524 3516 2576
rect 3568 2564 3574 2576
rect 7208 2573 7236 2604
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2632 9646 2644
rect 9640 2604 9996 2632
rect 9640 2592 9646 2604
rect 7101 2567 7159 2573
rect 7101 2564 7113 2567
rect 3568 2536 7113 2564
rect 3568 2524 3574 2536
rect 1578 2456 1584 2508
rect 1636 2496 1642 2508
rect 3418 2496 3424 2508
rect 1636 2468 3424 2496
rect 1636 2456 1642 2468
rect 3418 2456 3424 2468
rect 3476 2496 3482 2508
rect 4316 2499 4374 2505
rect 4316 2496 4328 2499
rect 3476 2468 4328 2496
rect 3476 2456 3482 2468
rect 4316 2465 4328 2468
rect 4362 2496 4374 2499
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 4362 2468 4721 2496
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 4709 2465 4721 2468
rect 4755 2465 4767 2499
rect 4709 2459 4767 2465
rect 5905 2499 5963 2505
rect 5905 2465 5917 2499
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 4264 2400 5273 2428
rect 4264 2372 4292 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 4246 2320 4252 2372
rect 4304 2320 4310 2372
rect 5169 2363 5227 2369
rect 5169 2329 5181 2363
rect 5215 2360 5227 2363
rect 5920 2360 5948 2459
rect 6932 2428 6960 2536
rect 7101 2533 7113 2536
rect 7147 2533 7159 2567
rect 7101 2527 7159 2533
rect 7193 2567 7251 2573
rect 7193 2533 7205 2567
rect 7239 2533 7251 2567
rect 7742 2564 7748 2576
rect 7703 2536 7748 2564
rect 7193 2527 7251 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 9968 2573 9996 2604
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 12805 2635 12863 2641
rect 12805 2632 12817 2635
rect 10376 2604 12817 2632
rect 10376 2592 10382 2604
rect 12805 2601 12817 2604
rect 12851 2601 12863 2635
rect 12805 2595 12863 2601
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2533 10011 2567
rect 9953 2527 10011 2533
rect 10505 2567 10563 2573
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 11238 2564 11244 2576
rect 10551 2536 11244 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8628 2468 9137 2496
rect 8628 2456 8634 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 11146 2496 11152 2508
rect 11107 2468 11152 2496
rect 9125 2459 9183 2465
rect 11146 2456 11152 2468
rect 11204 2456 11210 2508
rect 11330 2496 11336 2508
rect 11291 2468 11336 2496
rect 11330 2456 11336 2468
rect 11388 2496 11394 2508
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11388 2468 11897 2496
rect 11388 2456 11394 2468
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 11885 2459 11943 2465
rect 12618 2456 12624 2468
rect 12676 2496 12682 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12676 2468 13185 2496
rect 12676 2456 12682 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 6932 2400 8401 2428
rect 8389 2397 8401 2400
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 9907 2400 10793 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10781 2397 10793 2400
rect 10827 2397 10839 2431
rect 10781 2391 10839 2397
rect 7558 2360 7564 2372
rect 5215 2332 7564 2360
rect 5215 2329 5227 2332
rect 5169 2323 5227 2329
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 9876 2360 9904 2391
rect 11517 2363 11575 2369
rect 11517 2360 11529 2363
rect 8173 2332 9904 2360
rect 10520 2332 11529 2360
rect 6086 2252 6092 2304
rect 6144 2292 6150 2304
rect 8173 2292 8201 2332
rect 6144 2264 8201 2292
rect 6144 2252 6150 2264
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 8757 2295 8815 2301
rect 8757 2292 8769 2295
rect 8720 2264 8769 2292
rect 8720 2252 8726 2264
rect 8757 2261 8769 2264
rect 8803 2261 8815 2295
rect 8757 2255 8815 2261
rect 9858 2252 9864 2304
rect 9916 2292 9922 2304
rect 10520 2292 10548 2332
rect 11517 2329 11529 2332
rect 11563 2329 11575 2363
rect 11517 2323 11575 2329
rect 9916 2264 10548 2292
rect 9916 2252 9922 2264
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 2866 76 2872 128
rect 2924 116 2930 128
rect 5074 116 5080 128
rect 2924 88 5080 116
rect 2924 76 2930 88
rect 5074 76 5080 88
rect 5132 76 5138 128
<< via1 >>
rect 296 39584 348 39636
rect 1400 39584 1452 39636
rect 2136 39584 2188 39636
rect 6920 39584 6972 39636
rect 8852 39584 8904 39636
rect 3424 39516 3476 39568
rect 8392 39244 8444 39296
rect 9220 39244 9272 39296
rect 1492 38972 1544 39024
rect 2412 38972 2464 39024
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 8576 37068 8628 37120
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 11520 36864 11572 36916
rect 5356 36728 5408 36780
rect 3056 36660 3108 36712
rect 7196 36660 7248 36712
rect 7656 36660 7708 36712
rect 8576 36703 8628 36712
rect 8576 36669 8585 36703
rect 8585 36669 8619 36703
rect 8619 36669 8628 36703
rect 8576 36660 8628 36669
rect 10232 36592 10284 36644
rect 7196 36524 7248 36576
rect 8300 36567 8352 36576
rect 8300 36533 8309 36567
rect 8309 36533 8343 36567
rect 8343 36533 8352 36567
rect 8300 36524 8352 36533
rect 11152 36524 11204 36576
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 10416 36320 10468 36372
rect 12624 36320 12676 36372
rect 6644 36252 6696 36304
rect 9680 36227 9732 36236
rect 9680 36193 9689 36227
rect 9689 36193 9723 36227
rect 9723 36193 9732 36227
rect 9680 36184 9732 36193
rect 11244 36227 11296 36236
rect 11244 36193 11253 36227
rect 11253 36193 11287 36227
rect 11287 36193 11296 36227
rect 11244 36184 11296 36193
rect 7196 36159 7248 36168
rect 7196 36125 7205 36159
rect 7205 36125 7239 36159
rect 7239 36125 7248 36159
rect 7196 36116 7248 36125
rect 7748 36091 7800 36100
rect 7748 36057 7757 36091
rect 7757 36057 7791 36091
rect 7791 36057 7800 36091
rect 7748 36048 7800 36057
rect 8576 35980 8628 36032
rect 9496 35980 9548 36032
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 7196 35776 7248 35828
rect 11060 35776 11112 35828
rect 12072 35776 12124 35828
rect 13728 35776 13780 35828
rect 7748 35751 7800 35760
rect 7748 35717 7757 35751
rect 7757 35717 7791 35751
rect 7791 35717 7800 35751
rect 7748 35708 7800 35717
rect 7840 35572 7892 35624
rect 9496 35572 9548 35624
rect 10232 35615 10284 35624
rect 10232 35581 10241 35615
rect 10241 35581 10275 35615
rect 10275 35581 10284 35615
rect 10232 35572 10284 35581
rect 12440 35615 12492 35624
rect 7012 35504 7064 35556
rect 7196 35547 7248 35556
rect 7196 35513 7205 35547
rect 7205 35513 7239 35547
rect 7239 35513 7248 35547
rect 7196 35504 7248 35513
rect 6644 35479 6696 35488
rect 6644 35445 6653 35479
rect 6653 35445 6687 35479
rect 6687 35445 6696 35479
rect 6644 35436 6696 35445
rect 12440 35581 12449 35615
rect 12449 35581 12483 35615
rect 12483 35581 12492 35615
rect 12440 35572 12492 35581
rect 8760 35479 8812 35488
rect 8760 35445 8769 35479
rect 8769 35445 8803 35479
rect 8803 35445 8812 35479
rect 8760 35436 8812 35445
rect 9680 35436 9732 35488
rect 10692 35436 10744 35488
rect 11244 35436 11296 35488
rect 12072 35436 12124 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 1768 35232 1820 35284
rect 7012 35207 7064 35216
rect 7012 35173 7021 35207
rect 7021 35173 7055 35207
rect 7055 35173 7064 35207
rect 7012 35164 7064 35173
rect 12808 35232 12860 35284
rect 14096 35232 14148 35284
rect 9864 35164 9916 35216
rect 6184 35096 6236 35148
rect 8576 35139 8628 35148
rect 8576 35105 8620 35139
rect 8620 35105 8628 35139
rect 11520 35139 11572 35148
rect 8576 35096 8628 35105
rect 11520 35105 11529 35139
rect 11529 35105 11563 35139
rect 11563 35105 11572 35139
rect 11520 35096 11572 35105
rect 12716 35139 12768 35148
rect 12716 35105 12725 35139
rect 12725 35105 12759 35139
rect 12759 35105 12768 35139
rect 12716 35096 12768 35105
rect 7932 35028 7984 35080
rect 9404 35028 9456 35080
rect 10508 35071 10560 35080
rect 10508 35037 10517 35071
rect 10517 35037 10551 35071
rect 10551 35037 10560 35071
rect 10508 35028 10560 35037
rect 5264 34935 5316 34944
rect 5264 34901 5273 34935
rect 5273 34901 5307 34935
rect 5307 34901 5316 34935
rect 5264 34892 5316 34901
rect 7196 34892 7248 34944
rect 10876 34935 10928 34944
rect 10876 34901 10885 34935
rect 10885 34901 10919 34935
rect 10919 34901 10928 34935
rect 10876 34892 10928 34901
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 6184 34731 6236 34740
rect 6184 34697 6193 34731
rect 6193 34697 6227 34731
rect 6227 34697 6236 34731
rect 6184 34688 6236 34697
rect 7012 34688 7064 34740
rect 8576 34731 8628 34740
rect 8576 34697 8585 34731
rect 8585 34697 8619 34731
rect 8619 34697 8628 34731
rect 8576 34688 8628 34697
rect 15752 34688 15804 34740
rect 7196 34620 7248 34672
rect 756 34484 808 34536
rect 4344 34484 4396 34536
rect 5540 34552 5592 34604
rect 7840 34552 7892 34604
rect 8760 34552 8812 34604
rect 10876 34620 10928 34672
rect 12164 34620 12216 34672
rect 10968 34595 11020 34604
rect 10968 34561 10977 34595
rect 10977 34561 11011 34595
rect 11011 34561 11020 34595
rect 10968 34552 11020 34561
rect 12256 34552 12308 34604
rect 5264 34484 5316 34536
rect 7380 34484 7432 34536
rect 12716 34552 12768 34604
rect 13912 34484 13964 34536
rect 6736 34416 6788 34468
rect 10048 34416 10100 34468
rect 9864 34391 9916 34400
rect 9864 34357 9873 34391
rect 9873 34357 9907 34391
rect 9907 34357 9916 34391
rect 9864 34348 9916 34357
rect 10324 34391 10376 34400
rect 10324 34357 10333 34391
rect 10333 34357 10367 34391
rect 10367 34357 10376 34391
rect 11520 34416 11572 34468
rect 12348 34416 12400 34468
rect 10324 34348 10376 34357
rect 11980 34348 12032 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 5356 34187 5408 34196
rect 5356 34153 5365 34187
rect 5365 34153 5399 34187
rect 5399 34153 5408 34187
rect 5356 34144 5408 34153
rect 6184 34187 6236 34196
rect 6184 34153 6193 34187
rect 6193 34153 6227 34187
rect 6227 34153 6236 34187
rect 6184 34144 6236 34153
rect 6644 34144 6696 34196
rect 7012 34187 7064 34196
rect 7012 34153 7021 34187
rect 7021 34153 7055 34187
rect 7055 34153 7064 34187
rect 7012 34144 7064 34153
rect 7380 34187 7432 34196
rect 7380 34153 7389 34187
rect 7389 34153 7423 34187
rect 7423 34153 7432 34187
rect 7380 34144 7432 34153
rect 9404 34187 9456 34196
rect 9404 34153 9413 34187
rect 9413 34153 9447 34187
rect 9447 34153 9456 34187
rect 9404 34144 9456 34153
rect 10048 34187 10100 34196
rect 10048 34153 10057 34187
rect 10057 34153 10091 34187
rect 10091 34153 10100 34187
rect 10048 34144 10100 34153
rect 7840 34076 7892 34128
rect 10508 34076 10560 34128
rect 11520 34119 11572 34128
rect 11520 34085 11529 34119
rect 11529 34085 11563 34119
rect 11563 34085 11572 34119
rect 11520 34076 11572 34085
rect 14740 34144 14792 34196
rect 11704 34076 11756 34128
rect 3516 34008 3568 34060
rect 4804 34051 4856 34060
rect 4804 34017 4848 34051
rect 4848 34017 4856 34051
rect 4804 34008 4856 34017
rect 13544 34008 13596 34060
rect 5816 33983 5868 33992
rect 5816 33949 5825 33983
rect 5825 33949 5859 33983
rect 5859 33949 5868 33983
rect 5816 33940 5868 33949
rect 7932 33983 7984 33992
rect 7932 33949 7941 33983
rect 7941 33949 7975 33983
rect 7975 33949 7984 33983
rect 7932 33940 7984 33949
rect 9772 33940 9824 33992
rect 8852 33872 8904 33924
rect 12072 33915 12124 33924
rect 12072 33881 12081 33915
rect 12081 33881 12115 33915
rect 12115 33881 12124 33915
rect 12072 33872 12124 33881
rect 5632 33847 5684 33856
rect 5632 33813 5641 33847
rect 5641 33813 5675 33847
rect 5675 33813 5684 33847
rect 5632 33804 5684 33813
rect 8668 33847 8720 33856
rect 8668 33813 8677 33847
rect 8677 33813 8711 33847
rect 8711 33813 8720 33847
rect 8668 33804 8720 33813
rect 10692 33804 10744 33856
rect 12532 33847 12584 33856
rect 12532 33813 12541 33847
rect 12541 33813 12575 33847
rect 12575 33813 12584 33847
rect 12532 33804 12584 33813
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6184 33600 6236 33652
rect 6736 33600 6788 33652
rect 7840 33643 7892 33652
rect 7840 33609 7849 33643
rect 7849 33609 7883 33643
rect 7883 33609 7892 33643
rect 7840 33600 7892 33609
rect 8300 33643 8352 33652
rect 8300 33609 8309 33643
rect 8309 33609 8343 33643
rect 8343 33609 8352 33643
rect 8300 33600 8352 33609
rect 10048 33643 10100 33652
rect 10048 33609 10057 33643
rect 10057 33609 10091 33643
rect 10091 33609 10100 33643
rect 10048 33600 10100 33609
rect 11704 33643 11756 33652
rect 11704 33609 11713 33643
rect 11713 33609 11747 33643
rect 11747 33609 11756 33643
rect 11704 33600 11756 33609
rect 5816 33464 5868 33516
rect 7932 33464 7984 33516
rect 4068 33439 4120 33448
rect 4068 33405 4077 33439
rect 4077 33405 4111 33439
rect 4111 33405 4120 33439
rect 4068 33396 4120 33405
rect 5080 33396 5132 33448
rect 5264 33396 5316 33448
rect 10324 33532 10376 33584
rect 5356 33328 5408 33380
rect 4804 33303 4856 33312
rect 4804 33269 4813 33303
rect 4813 33269 4847 33303
rect 4847 33269 4856 33303
rect 4804 33260 4856 33269
rect 10692 33396 10744 33448
rect 5724 33328 5776 33380
rect 7012 33371 7064 33380
rect 7012 33337 7021 33371
rect 7021 33337 7055 33371
rect 7055 33337 7064 33371
rect 8668 33371 8720 33380
rect 7012 33328 7064 33337
rect 8668 33337 8677 33371
rect 8677 33337 8711 33371
rect 8711 33337 8720 33371
rect 8668 33328 8720 33337
rect 10048 33328 10100 33380
rect 12532 33507 12584 33516
rect 12532 33473 12541 33507
rect 12541 33473 12575 33507
rect 12575 33473 12584 33507
rect 12532 33464 12584 33473
rect 12808 33507 12860 33516
rect 12808 33473 12817 33507
rect 12817 33473 12851 33507
rect 12851 33473 12860 33507
rect 12808 33464 12860 33473
rect 5816 33260 5868 33312
rect 11428 33303 11480 33312
rect 11428 33269 11437 33303
rect 11437 33269 11471 33303
rect 11471 33269 11480 33303
rect 11428 33260 11480 33269
rect 13544 33303 13596 33312
rect 13544 33269 13553 33303
rect 13553 33269 13587 33303
rect 13587 33269 13596 33303
rect 13544 33260 13596 33269
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 4068 33056 4120 33108
rect 5632 33056 5684 33108
rect 8852 33099 8904 33108
rect 8852 33065 8861 33099
rect 8861 33065 8895 33099
rect 8895 33065 8904 33099
rect 8852 33056 8904 33065
rect 11520 33099 11572 33108
rect 11520 33065 11529 33099
rect 11529 33065 11563 33099
rect 11563 33065 11572 33099
rect 11520 33056 11572 33065
rect 6184 32988 6236 33040
rect 8024 33031 8076 33040
rect 8024 32997 8033 33031
rect 8033 32997 8067 33031
rect 8067 32997 8076 33031
rect 8024 32988 8076 32997
rect 10324 33031 10376 33040
rect 10324 32997 10333 33031
rect 10333 32997 10367 33031
rect 10367 32997 10376 33031
rect 10324 32988 10376 32997
rect 10968 32988 11020 33040
rect 11428 32988 11480 33040
rect 12072 32988 12124 33040
rect 12256 32988 12308 33040
rect 12808 32988 12860 33040
rect 4252 32920 4304 32972
rect 5172 32920 5224 32972
rect 13544 32920 13596 32972
rect 5080 32852 5132 32904
rect 5632 32852 5684 32904
rect 5908 32852 5960 32904
rect 7932 32895 7984 32904
rect 7932 32861 7941 32895
rect 7941 32861 7975 32895
rect 7975 32861 7984 32895
rect 7932 32852 7984 32861
rect 8208 32895 8260 32904
rect 8208 32861 8217 32895
rect 8217 32861 8251 32895
rect 8251 32861 8260 32895
rect 8208 32852 8260 32861
rect 9680 32852 9732 32904
rect 12072 32852 12124 32904
rect 4896 32784 4948 32836
rect 8576 32784 8628 32836
rect 5816 32716 5868 32768
rect 7012 32759 7064 32768
rect 7012 32725 7021 32759
rect 7021 32725 7055 32759
rect 7055 32725 7064 32759
rect 7012 32716 7064 32725
rect 7380 32759 7432 32768
rect 7380 32725 7389 32759
rect 7389 32725 7423 32759
rect 7423 32725 7432 32759
rect 7380 32716 7432 32725
rect 9772 32716 9824 32768
rect 9956 32759 10008 32768
rect 9956 32725 9965 32759
rect 9965 32725 9999 32759
rect 9999 32725 10008 32759
rect 9956 32716 10008 32725
rect 10048 32716 10100 32768
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 8024 32512 8076 32564
rect 9864 32555 9916 32564
rect 9864 32521 9873 32555
rect 9873 32521 9907 32555
rect 9907 32521 9916 32555
rect 9864 32512 9916 32521
rect 10324 32512 10376 32564
rect 11428 32512 11480 32564
rect 12072 32555 12124 32564
rect 12072 32521 12081 32555
rect 12081 32521 12115 32555
rect 12115 32521 12124 32555
rect 12072 32512 12124 32521
rect 12164 32512 12216 32564
rect 5172 32444 5224 32496
rect 7564 32444 7616 32496
rect 9680 32444 9732 32496
rect 4252 32351 4304 32360
rect 4252 32317 4270 32351
rect 4270 32317 4304 32351
rect 4252 32308 4304 32317
rect 5632 32308 5684 32360
rect 5816 32376 5868 32428
rect 10048 32419 10100 32428
rect 10048 32385 10057 32419
rect 10057 32385 10091 32419
rect 10091 32385 10100 32419
rect 10048 32376 10100 32385
rect 10968 32376 11020 32428
rect 6000 32308 6052 32360
rect 7380 32351 7432 32360
rect 7380 32317 7389 32351
rect 7389 32317 7423 32351
rect 7423 32317 7432 32351
rect 7380 32308 7432 32317
rect 12164 32308 12216 32360
rect 5908 32283 5960 32292
rect 5908 32249 5917 32283
rect 5917 32249 5951 32283
rect 5951 32249 5960 32283
rect 5908 32240 5960 32249
rect 4528 32172 4580 32224
rect 6184 32172 6236 32224
rect 7104 32172 7156 32224
rect 9864 32172 9916 32224
rect 13544 32172 13596 32224
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 5908 31968 5960 32020
rect 8116 31968 8168 32020
rect 9680 31968 9732 32020
rect 9956 32011 10008 32020
rect 9956 31977 9965 32011
rect 9965 31977 9999 32011
rect 9999 31977 10008 32011
rect 9956 31968 10008 31977
rect 12532 31968 12584 32020
rect 572 31900 624 31952
rect 6000 31943 6052 31952
rect 6000 31909 6009 31943
rect 6009 31909 6043 31943
rect 6043 31909 6052 31943
rect 6000 31900 6052 31909
rect 7012 31943 7064 31952
rect 7012 31909 7021 31943
rect 7021 31909 7055 31943
rect 7055 31909 7064 31943
rect 7012 31900 7064 31909
rect 7932 31900 7984 31952
rect 3976 31875 4028 31884
rect 3976 31841 3985 31875
rect 3985 31841 4019 31875
rect 4019 31841 4028 31875
rect 3976 31832 4028 31841
rect 5632 31832 5684 31884
rect 5816 31875 5868 31884
rect 5816 31841 5825 31875
rect 5825 31841 5859 31875
rect 5859 31841 5868 31875
rect 5816 31832 5868 31841
rect 8576 31832 8628 31884
rect 9680 31875 9732 31884
rect 4528 31764 4580 31816
rect 6552 31764 6604 31816
rect 6736 31696 6788 31748
rect 9680 31841 9689 31875
rect 9689 31841 9723 31875
rect 9723 31841 9732 31875
rect 9680 31832 9732 31841
rect 11152 31832 11204 31884
rect 11336 31832 11388 31884
rect 4160 31628 4212 31680
rect 8484 31628 8536 31680
rect 9496 31628 9548 31680
rect 10876 31628 10928 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 6552 31467 6604 31476
rect 6552 31433 6561 31467
rect 6561 31433 6595 31467
rect 6595 31433 6604 31467
rect 6552 31424 6604 31433
rect 7012 31467 7064 31476
rect 7012 31433 7021 31467
rect 7021 31433 7055 31467
rect 7055 31433 7064 31467
rect 7012 31424 7064 31433
rect 9680 31424 9732 31476
rect 8116 31356 8168 31408
rect 8208 31331 8260 31340
rect 8208 31297 8217 31331
rect 8217 31297 8251 31331
rect 8251 31297 8260 31331
rect 8208 31288 8260 31297
rect 10968 31288 11020 31340
rect 12256 31288 12308 31340
rect 5908 31220 5960 31272
rect 9036 31263 9088 31272
rect 9036 31229 9045 31263
rect 9045 31229 9079 31263
rect 9079 31229 9088 31263
rect 9036 31220 9088 31229
rect 9496 31263 9548 31272
rect 9496 31229 9505 31263
rect 9505 31229 9539 31263
rect 9539 31229 9548 31263
rect 9496 31220 9548 31229
rect 3976 31152 4028 31204
rect 5356 31152 5408 31204
rect 5816 31152 5868 31204
rect 7288 31152 7340 31204
rect 7748 31152 7800 31204
rect 9772 31195 9824 31204
rect 9772 31161 9781 31195
rect 9781 31161 9815 31195
rect 9815 31161 9824 31195
rect 9772 31152 9824 31161
rect 10876 31195 10928 31204
rect 10876 31161 10885 31195
rect 10885 31161 10919 31195
rect 10919 31161 10928 31195
rect 10876 31152 10928 31161
rect 4896 31127 4948 31136
rect 4896 31093 4905 31127
rect 4905 31093 4939 31127
rect 4939 31093 4948 31127
rect 4896 31084 4948 31093
rect 5632 31084 5684 31136
rect 6736 31084 6788 31136
rect 8576 31084 8628 31136
rect 9496 31084 9548 31136
rect 11336 31084 11388 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 8300 30880 8352 30932
rect 8760 30880 8812 30932
rect 10048 30923 10100 30932
rect 10048 30889 10057 30923
rect 10057 30889 10091 30923
rect 10091 30889 10100 30923
rect 10048 30880 10100 30889
rect 10876 30880 10928 30932
rect 10968 30923 11020 30932
rect 10968 30889 10977 30923
rect 10977 30889 11011 30923
rect 11011 30889 11020 30923
rect 10968 30880 11020 30889
rect 4896 30812 4948 30864
rect 7840 30855 7892 30864
rect 7840 30821 7849 30855
rect 7849 30821 7883 30855
rect 7883 30821 7892 30855
rect 7840 30812 7892 30821
rect 11612 30855 11664 30864
rect 11612 30821 11621 30855
rect 11621 30821 11655 30855
rect 11655 30821 11664 30855
rect 11612 30812 11664 30821
rect 12256 30812 12308 30864
rect 6092 30744 6144 30796
rect 6460 30787 6512 30796
rect 6460 30753 6469 30787
rect 6469 30753 6503 30787
rect 6503 30753 6512 30787
rect 6460 30744 6512 30753
rect 6920 30744 6972 30796
rect 3976 30676 4028 30728
rect 5356 30719 5408 30728
rect 5356 30685 5365 30719
rect 5365 30685 5399 30719
rect 5399 30685 5408 30719
rect 5356 30676 5408 30685
rect 8024 30676 8076 30728
rect 8208 30719 8260 30728
rect 8208 30685 8217 30719
rect 8217 30685 8251 30719
rect 8251 30685 8260 30719
rect 8208 30676 8260 30685
rect 8576 30676 8628 30728
rect 8760 30676 8812 30728
rect 10876 30676 10928 30728
rect 11520 30719 11572 30728
rect 11520 30685 11529 30719
rect 11529 30685 11563 30719
rect 11563 30685 11572 30719
rect 11520 30676 11572 30685
rect 6920 30608 6972 30660
rect 9036 30651 9088 30660
rect 9036 30617 9045 30651
rect 9045 30617 9079 30651
rect 9079 30617 9088 30651
rect 9036 30608 9088 30617
rect 5908 30540 5960 30592
rect 6184 30540 6236 30592
rect 7104 30583 7156 30592
rect 7104 30549 7113 30583
rect 7113 30549 7147 30583
rect 7147 30549 7156 30583
rect 7104 30540 7156 30549
rect 7748 30540 7800 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 3976 30336 4028 30388
rect 4896 30336 4948 30388
rect 7748 30379 7800 30388
rect 7748 30345 7757 30379
rect 7757 30345 7791 30379
rect 7791 30345 7800 30379
rect 7748 30336 7800 30345
rect 8024 30379 8076 30388
rect 8024 30345 8033 30379
rect 8033 30345 8067 30379
rect 8067 30345 8076 30379
rect 8024 30336 8076 30345
rect 9312 30336 9364 30388
rect 10876 30379 10928 30388
rect 10876 30345 10885 30379
rect 10885 30345 10919 30379
rect 10919 30345 10928 30379
rect 10876 30336 10928 30345
rect 11520 30379 11572 30388
rect 11520 30345 11529 30379
rect 11529 30345 11563 30379
rect 11563 30345 11572 30379
rect 11520 30336 11572 30345
rect 11612 30268 11664 30320
rect 5356 30243 5408 30252
rect 5356 30209 5365 30243
rect 5365 30209 5399 30243
rect 5399 30209 5408 30243
rect 5356 30200 5408 30209
rect 9772 30200 9824 30252
rect 7012 30132 7064 30184
rect 8576 30132 8628 30184
rect 5080 30107 5132 30116
rect 5080 30073 5089 30107
rect 5089 30073 5123 30107
rect 5123 30073 5132 30107
rect 5080 30064 5132 30073
rect 5908 30064 5960 30116
rect 6460 30064 6512 30116
rect 7104 30107 7156 30116
rect 7104 30073 7113 30107
rect 7113 30073 7147 30107
rect 7147 30073 7156 30107
rect 7104 30064 7156 30073
rect 7472 29996 7524 30048
rect 8300 29996 8352 30048
rect 10048 30064 10100 30116
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 5080 29792 5132 29844
rect 5356 29792 5408 29844
rect 7840 29835 7892 29844
rect 7840 29801 7849 29835
rect 7849 29801 7883 29835
rect 7883 29801 7892 29835
rect 7840 29792 7892 29801
rect 8024 29792 8076 29844
rect 9772 29792 9824 29844
rect 11520 29792 11572 29844
rect 4068 29724 4120 29776
rect 6552 29724 6604 29776
rect 7104 29724 7156 29776
rect 10048 29724 10100 29776
rect 12440 29724 12492 29776
rect 12256 29699 12308 29708
rect 12256 29665 12265 29699
rect 12265 29665 12299 29699
rect 12299 29665 12308 29699
rect 12256 29656 12308 29665
rect 3056 29588 3108 29640
rect 4620 29588 4672 29640
rect 6644 29631 6696 29640
rect 6644 29597 6653 29631
rect 6653 29597 6687 29631
rect 6687 29597 6696 29631
rect 6644 29588 6696 29597
rect 9772 29631 9824 29640
rect 9772 29597 9781 29631
rect 9781 29597 9815 29631
rect 9815 29597 9824 29631
rect 9772 29588 9824 29597
rect 12440 29588 12492 29640
rect 5356 29563 5408 29572
rect 5356 29529 5365 29563
rect 5365 29529 5399 29563
rect 5399 29529 5408 29563
rect 5356 29520 5408 29529
rect 4988 29452 5040 29504
rect 6092 29452 6144 29504
rect 10416 29452 10468 29504
rect 10784 29452 10836 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 4252 29248 4304 29300
rect 12256 29248 12308 29300
rect 4620 29180 4672 29232
rect 5080 29180 5132 29232
rect 6552 29223 6604 29232
rect 6552 29189 6561 29223
rect 6561 29189 6595 29223
rect 6595 29189 6604 29223
rect 6552 29180 6604 29189
rect 8300 29180 8352 29232
rect 4988 29155 5040 29164
rect 4988 29121 4997 29155
rect 4997 29121 5031 29155
rect 5031 29121 5040 29155
rect 4988 29112 5040 29121
rect 5356 29155 5408 29164
rect 5356 29121 5365 29155
rect 5365 29121 5399 29155
rect 5399 29121 5408 29155
rect 5356 29112 5408 29121
rect 10876 29155 10928 29164
rect 10876 29121 10885 29155
rect 10885 29121 10919 29155
rect 10919 29121 10928 29155
rect 10876 29112 10928 29121
rect 3056 28951 3108 28960
rect 3056 28917 3065 28951
rect 3065 28917 3099 28951
rect 3099 28917 3108 28951
rect 3056 28908 3108 28917
rect 4804 28976 4856 29028
rect 4344 28908 4396 28960
rect 4528 28908 4580 28960
rect 4712 28951 4764 28960
rect 4712 28917 4721 28951
rect 4721 28917 4755 28951
rect 4755 28917 4764 28951
rect 4712 28908 4764 28917
rect 5632 28908 5684 28960
rect 6920 29044 6972 29096
rect 7288 29087 7340 29096
rect 7288 29053 7297 29087
rect 7297 29053 7331 29087
rect 7331 29053 7340 29087
rect 7288 29044 7340 29053
rect 8300 28976 8352 29028
rect 6644 28908 6696 28960
rect 8024 28951 8076 28960
rect 8024 28917 8033 28951
rect 8033 28917 8067 28951
rect 8067 28917 8076 28951
rect 8024 28908 8076 28917
rect 10048 28908 10100 28960
rect 12256 29044 12308 29096
rect 13728 29044 13780 29096
rect 10416 29019 10468 29028
rect 10416 28985 10425 29019
rect 10425 28985 10459 29019
rect 10459 28985 10468 29019
rect 10416 28976 10468 28985
rect 11520 28976 11572 29028
rect 10692 28908 10744 28960
rect 13360 28908 13412 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 4620 28747 4672 28756
rect 4620 28713 4629 28747
rect 4629 28713 4663 28747
rect 4663 28713 4672 28747
rect 4620 28704 4672 28713
rect 6644 28704 6696 28756
rect 9772 28704 9824 28756
rect 13360 28704 13412 28756
rect 4068 28636 4120 28688
rect 4712 28679 4764 28688
rect 4712 28645 4721 28679
rect 4721 28645 4755 28679
rect 4755 28645 4764 28679
rect 4712 28636 4764 28645
rect 7012 28679 7064 28688
rect 7012 28645 7021 28679
rect 7021 28645 7055 28679
rect 7055 28645 7064 28679
rect 7012 28636 7064 28645
rect 8760 28679 8812 28688
rect 8760 28645 8769 28679
rect 8769 28645 8803 28679
rect 8803 28645 8812 28679
rect 8760 28636 8812 28645
rect 11152 28636 11204 28688
rect 12440 28679 12492 28688
rect 12440 28645 12449 28679
rect 12449 28645 12483 28679
rect 12483 28645 12492 28679
rect 12440 28636 12492 28645
rect 4804 28611 4856 28620
rect 4804 28577 4813 28611
rect 4813 28577 4847 28611
rect 4847 28577 4856 28611
rect 4804 28568 4856 28577
rect 6276 28500 6328 28552
rect 6644 28568 6696 28620
rect 7288 28611 7340 28620
rect 7288 28577 7297 28611
rect 7297 28577 7331 28611
rect 7331 28577 7340 28611
rect 7288 28568 7340 28577
rect 8116 28611 8168 28620
rect 8116 28577 8125 28611
rect 8125 28577 8159 28611
rect 8159 28577 8168 28611
rect 8116 28568 8168 28577
rect 8484 28611 8536 28620
rect 8484 28577 8493 28611
rect 8493 28577 8527 28611
rect 8527 28577 8536 28611
rect 8484 28568 8536 28577
rect 10876 28611 10928 28620
rect 10876 28577 10885 28611
rect 10885 28577 10919 28611
rect 10919 28577 10928 28611
rect 13268 28611 13320 28620
rect 10876 28568 10928 28577
rect 13268 28577 13277 28611
rect 13277 28577 13311 28611
rect 13311 28577 13320 28611
rect 13268 28568 13320 28577
rect 10324 28500 10376 28552
rect 12624 28364 12676 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 4804 28160 4856 28212
rect 6276 28203 6328 28212
rect 6276 28169 6285 28203
rect 6285 28169 6319 28203
rect 6319 28169 6328 28203
rect 6276 28160 6328 28169
rect 8300 28203 8352 28212
rect 8300 28169 8309 28203
rect 8309 28169 8343 28203
rect 8343 28169 8352 28203
rect 8300 28160 8352 28169
rect 8484 28160 8536 28212
rect 10692 28160 10744 28212
rect 11152 28203 11204 28212
rect 11152 28169 11161 28203
rect 11161 28169 11195 28203
rect 11195 28169 11204 28203
rect 11152 28160 11204 28169
rect 12348 28160 12400 28212
rect 13268 28160 13320 28212
rect 4068 28092 4120 28144
rect 6092 28092 6144 28144
rect 7472 28092 7524 28144
rect 5540 28024 5592 28076
rect 3976 27956 4028 28008
rect 4988 27999 5040 28008
rect 4988 27965 4997 27999
rect 4997 27965 5031 27999
rect 5031 27965 5040 27999
rect 4988 27956 5040 27965
rect 5080 27956 5132 28008
rect 8116 28024 8168 28076
rect 9680 28024 9732 28076
rect 7196 27956 7248 28008
rect 8484 27999 8536 28008
rect 5080 27820 5132 27872
rect 7012 27888 7064 27940
rect 8484 27965 8493 27999
rect 8493 27965 8527 27999
rect 8527 27965 8536 27999
rect 8484 27956 8536 27965
rect 8576 27888 8628 27940
rect 7472 27820 7524 27872
rect 8300 27820 8352 27872
rect 10048 27956 10100 28008
rect 10232 27999 10284 28008
rect 10232 27965 10241 27999
rect 10241 27965 10275 27999
rect 10275 27965 10284 27999
rect 10232 27956 10284 27965
rect 8852 27888 8904 27940
rect 9864 27888 9916 27940
rect 10600 27931 10652 27940
rect 10600 27897 10603 27931
rect 10603 27897 10637 27931
rect 10637 27897 10652 27931
rect 10600 27888 10652 27897
rect 10508 27820 10560 27872
rect 12716 27863 12768 27872
rect 12716 27829 12725 27863
rect 12725 27829 12759 27863
rect 12759 27829 12768 27863
rect 12716 27820 12768 27829
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4988 27616 5040 27668
rect 7012 27659 7064 27668
rect 7012 27625 7021 27659
rect 7021 27625 7055 27659
rect 7055 27625 7064 27659
rect 7012 27616 7064 27625
rect 8024 27659 8076 27668
rect 8024 27625 8033 27659
rect 8033 27625 8067 27659
rect 8067 27625 8076 27659
rect 8024 27616 8076 27625
rect 8484 27616 8536 27668
rect 10416 27616 10468 27668
rect 12624 27659 12676 27668
rect 6184 27548 6236 27600
rect 10048 27548 10100 27600
rect 10876 27548 10928 27600
rect 11704 27591 11756 27600
rect 11704 27557 11713 27591
rect 11713 27557 11747 27591
rect 11747 27557 11756 27591
rect 11704 27548 11756 27557
rect 12624 27625 12633 27659
rect 12633 27625 12667 27659
rect 12667 27625 12676 27659
rect 12624 27616 12676 27625
rect 4068 27480 4120 27532
rect 4160 27523 4212 27532
rect 4160 27489 4169 27523
rect 4169 27489 4203 27523
rect 4203 27489 4212 27523
rect 4160 27480 4212 27489
rect 5540 27480 5592 27532
rect 6000 27523 6052 27532
rect 6000 27489 6009 27523
rect 6009 27489 6043 27523
rect 6043 27489 6052 27523
rect 6000 27480 6052 27489
rect 7932 27523 7984 27532
rect 7932 27489 7941 27523
rect 7941 27489 7975 27523
rect 7975 27489 7984 27523
rect 7932 27480 7984 27489
rect 8576 27480 8628 27532
rect 12440 27480 12492 27532
rect 13084 27523 13136 27532
rect 13084 27489 13093 27523
rect 13093 27489 13127 27523
rect 13127 27489 13136 27523
rect 13084 27480 13136 27489
rect 6184 27412 6236 27464
rect 10140 27412 10192 27464
rect 10784 27412 10836 27464
rect 11612 27455 11664 27464
rect 11612 27421 11621 27455
rect 11621 27421 11655 27455
rect 11655 27421 11664 27455
rect 11612 27412 11664 27421
rect 10232 27344 10284 27396
rect 5080 27319 5132 27328
rect 5080 27285 5089 27319
rect 5089 27285 5123 27319
rect 5123 27285 5132 27319
rect 5080 27276 5132 27285
rect 6644 27319 6696 27328
rect 6644 27285 6653 27319
rect 6653 27285 6687 27319
rect 6687 27285 6696 27319
rect 6644 27276 6696 27285
rect 10324 27276 10376 27328
rect 11796 27276 11848 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 4160 27115 4212 27124
rect 4160 27081 4169 27115
rect 4169 27081 4203 27115
rect 4203 27081 4212 27115
rect 5908 27115 5960 27124
rect 4160 27072 4212 27081
rect 5908 27081 5917 27115
rect 5917 27081 5951 27115
rect 5951 27081 5960 27115
rect 5908 27072 5960 27081
rect 6184 27115 6236 27124
rect 6184 27081 6193 27115
rect 6193 27081 6227 27115
rect 6227 27081 6236 27115
rect 6184 27072 6236 27081
rect 6644 27072 6696 27124
rect 10048 27115 10100 27124
rect 10048 27081 10057 27115
rect 10057 27081 10091 27115
rect 10091 27081 10100 27115
rect 10048 27072 10100 27081
rect 11704 27072 11756 27124
rect 11796 27072 11848 27124
rect 13084 27115 13136 27124
rect 13084 27081 13093 27115
rect 13093 27081 13127 27115
rect 13127 27081 13136 27115
rect 13084 27072 13136 27081
rect 5448 27004 5500 27056
rect 7932 27004 7984 27056
rect 11244 27004 11296 27056
rect 12808 27004 12860 27056
rect 4712 26936 4764 26988
rect 6000 26936 6052 26988
rect 7288 26936 7340 26988
rect 10232 26936 10284 26988
rect 10876 26936 10928 26988
rect 12072 26936 12124 26988
rect 4988 26911 5040 26920
rect 4988 26877 4997 26911
rect 4997 26877 5031 26911
rect 5031 26877 5040 26911
rect 4988 26868 5040 26877
rect 5080 26800 5132 26852
rect 6092 26800 6144 26852
rect 10600 26843 10652 26852
rect 10600 26809 10609 26843
rect 10609 26809 10643 26843
rect 10643 26809 10652 26843
rect 10600 26800 10652 26809
rect 11244 26800 11296 26852
rect 5724 26732 5776 26784
rect 7840 26775 7892 26784
rect 7840 26741 7849 26775
rect 7849 26741 7883 26775
rect 7883 26741 7892 26775
rect 7840 26732 7892 26741
rect 8576 26732 8628 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 10140 26528 10192 26580
rect 10600 26528 10652 26580
rect 10968 26528 11020 26580
rect 11520 26571 11572 26580
rect 4068 26460 4120 26512
rect 8392 26460 8444 26512
rect 10324 26460 10376 26512
rect 10692 26503 10744 26512
rect 10692 26469 10701 26503
rect 10701 26469 10735 26503
rect 10735 26469 10744 26503
rect 10692 26460 10744 26469
rect 11244 26503 11296 26512
rect 11244 26469 11253 26503
rect 11253 26469 11287 26503
rect 11287 26469 11296 26503
rect 11244 26460 11296 26469
rect 11520 26537 11529 26571
rect 11529 26537 11563 26571
rect 11563 26537 11572 26571
rect 11520 26528 11572 26537
rect 4896 26435 4948 26444
rect 4896 26401 4905 26435
rect 4905 26401 4939 26435
rect 4939 26401 4948 26435
rect 4896 26392 4948 26401
rect 6460 26392 6512 26444
rect 6920 26392 6972 26444
rect 7380 26392 7432 26444
rect 8024 26435 8076 26444
rect 8024 26401 8033 26435
rect 8033 26401 8067 26435
rect 8067 26401 8076 26435
rect 8024 26392 8076 26401
rect 8576 26435 8628 26444
rect 8576 26401 8585 26435
rect 8585 26401 8619 26435
rect 8619 26401 8628 26435
rect 8576 26392 8628 26401
rect 12072 26435 12124 26444
rect 12072 26401 12116 26435
rect 12116 26401 12124 26435
rect 12072 26392 12124 26401
rect 7104 26367 7156 26376
rect 7104 26333 7113 26367
rect 7113 26333 7147 26367
rect 7147 26333 7156 26367
rect 7104 26324 7156 26333
rect 8760 26367 8812 26376
rect 8760 26333 8769 26367
rect 8769 26333 8803 26367
rect 8803 26333 8812 26367
rect 8760 26324 8812 26333
rect 10784 26324 10836 26376
rect 7564 26256 7616 26308
rect 8392 26256 8444 26308
rect 4988 26188 5040 26240
rect 5356 26188 5408 26240
rect 5540 26188 5592 26240
rect 9312 26231 9364 26240
rect 9312 26197 9321 26231
rect 9321 26197 9355 26231
rect 9355 26197 9364 26231
rect 9312 26188 9364 26197
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4896 26027 4948 26036
rect 4896 25993 4905 26027
rect 4905 25993 4939 26027
rect 4939 25993 4948 26027
rect 4896 25984 4948 25993
rect 6460 26027 6512 26036
rect 6460 25993 6469 26027
rect 6469 25993 6503 26027
rect 6503 25993 6512 26027
rect 6460 25984 6512 25993
rect 8852 25984 8904 26036
rect 10600 25984 10652 26036
rect 10692 25984 10744 26036
rect 11980 25984 12032 26036
rect 12072 26027 12124 26036
rect 12072 25993 12081 26027
rect 12081 25993 12115 26027
rect 12115 25993 12124 26027
rect 12072 25984 12124 25993
rect 6092 25848 6144 25900
rect 5540 25823 5592 25832
rect 5540 25789 5549 25823
rect 5549 25789 5583 25823
rect 5583 25789 5592 25823
rect 5540 25780 5592 25789
rect 9312 25823 9364 25832
rect 5080 25644 5132 25696
rect 5632 25712 5684 25764
rect 9312 25789 9321 25823
rect 9321 25789 9355 25823
rect 9355 25789 9364 25823
rect 9312 25780 9364 25789
rect 9772 25780 9824 25832
rect 11244 25780 11296 25832
rect 9404 25712 9456 25764
rect 8576 25644 8628 25696
rect 10048 25644 10100 25696
rect 10784 25644 10836 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 5356 25483 5408 25492
rect 5356 25449 5365 25483
rect 5365 25449 5399 25483
rect 5399 25449 5408 25483
rect 5356 25440 5408 25449
rect 6000 25440 6052 25492
rect 7104 25483 7156 25492
rect 7104 25449 7113 25483
rect 7113 25449 7147 25483
rect 7147 25449 7156 25483
rect 7104 25440 7156 25449
rect 8760 25440 8812 25492
rect 9404 25483 9456 25492
rect 9404 25449 9413 25483
rect 9413 25449 9447 25483
rect 9447 25449 9456 25483
rect 9404 25440 9456 25449
rect 10048 25483 10100 25492
rect 10048 25449 10057 25483
rect 10057 25449 10091 25483
rect 10091 25449 10100 25483
rect 10048 25440 10100 25449
rect 10692 25440 10744 25492
rect 10784 25440 10836 25492
rect 5540 25347 5592 25356
rect 5540 25313 5549 25347
rect 5549 25313 5583 25347
rect 5583 25313 5592 25347
rect 5540 25304 5592 25313
rect 5908 25304 5960 25356
rect 6092 25347 6144 25356
rect 6092 25313 6101 25347
rect 6101 25313 6135 25347
rect 6135 25313 6144 25347
rect 6092 25304 6144 25313
rect 7288 25347 7340 25356
rect 7288 25313 7297 25347
rect 7297 25313 7331 25347
rect 7331 25313 7340 25347
rect 11244 25372 11296 25424
rect 7288 25304 7340 25313
rect 10876 25304 10928 25356
rect 12440 25304 12492 25356
rect 6184 25279 6236 25288
rect 6184 25245 6193 25279
rect 6193 25245 6227 25279
rect 6227 25245 6236 25279
rect 6184 25236 6236 25245
rect 4436 25143 4488 25152
rect 4436 25109 4445 25143
rect 4445 25109 4479 25143
rect 4479 25109 4488 25143
rect 4436 25100 4488 25109
rect 5172 25100 5224 25152
rect 6736 25100 6788 25152
rect 8024 25100 8076 25152
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 4436 24896 4488 24948
rect 7104 24828 7156 24880
rect 12256 24896 12308 24948
rect 8484 24828 8536 24880
rect 8852 24871 8904 24880
rect 8852 24837 8861 24871
rect 8861 24837 8895 24871
rect 8895 24837 8904 24871
rect 8852 24828 8904 24837
rect 4804 24760 4856 24812
rect 7012 24760 7064 24812
rect 8760 24760 8812 24812
rect 3976 24735 4028 24744
rect 3976 24701 3985 24735
rect 3985 24701 4019 24735
rect 4019 24701 4028 24735
rect 3976 24692 4028 24701
rect 5356 24735 5408 24744
rect 5356 24701 5362 24735
rect 5362 24701 5408 24735
rect 5356 24692 5408 24701
rect 5448 24692 5500 24744
rect 6736 24692 6788 24744
rect 7288 24692 7340 24744
rect 3148 24556 3200 24608
rect 4344 24667 4396 24676
rect 4344 24633 4353 24667
rect 4353 24633 4387 24667
rect 4387 24633 4396 24667
rect 4344 24624 4396 24633
rect 5172 24667 5224 24676
rect 5172 24633 5181 24667
rect 5181 24633 5215 24667
rect 5215 24633 5224 24667
rect 5172 24624 5224 24633
rect 5908 24667 5960 24676
rect 5908 24633 5917 24667
rect 5917 24633 5951 24667
rect 5951 24633 5960 24667
rect 5908 24624 5960 24633
rect 5080 24556 5132 24608
rect 8944 24624 8996 24676
rect 9404 24667 9456 24676
rect 9404 24633 9407 24667
rect 9407 24633 9441 24667
rect 9441 24633 9456 24667
rect 10876 24803 10928 24812
rect 10876 24769 10885 24803
rect 10885 24769 10919 24803
rect 10919 24769 10928 24803
rect 10876 24760 10928 24769
rect 11244 24803 11296 24812
rect 11244 24769 11253 24803
rect 11253 24769 11287 24803
rect 11287 24769 11296 24803
rect 11244 24760 11296 24769
rect 9404 24624 9456 24633
rect 8484 24599 8536 24608
rect 8484 24565 8493 24599
rect 8493 24565 8527 24599
rect 8527 24565 8536 24599
rect 8484 24556 8536 24565
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 2780 24216 2832 24268
rect 7288 24352 7340 24404
rect 8024 24352 8076 24404
rect 9772 24395 9824 24404
rect 9772 24361 9781 24395
rect 9781 24361 9815 24395
rect 9815 24361 9824 24395
rect 9772 24352 9824 24361
rect 9956 24352 10008 24404
rect 5356 24284 5408 24336
rect 4252 24259 4304 24268
rect 4252 24225 4261 24259
rect 4261 24225 4295 24259
rect 4295 24225 4304 24259
rect 4252 24216 4304 24225
rect 5724 24259 5776 24268
rect 5724 24225 5733 24259
rect 5733 24225 5767 24259
rect 5767 24225 5776 24259
rect 7104 24284 7156 24336
rect 8484 24284 8536 24336
rect 5724 24216 5776 24225
rect 7012 24259 7064 24268
rect 7012 24225 7021 24259
rect 7021 24225 7055 24259
rect 7055 24225 7064 24259
rect 7012 24216 7064 24225
rect 3976 24148 4028 24200
rect 4344 24148 4396 24200
rect 9312 24216 9364 24268
rect 9680 24259 9732 24268
rect 9680 24225 9689 24259
rect 9689 24225 9723 24259
rect 9723 24225 9732 24259
rect 9680 24216 9732 24225
rect 10140 24259 10192 24268
rect 10140 24225 10149 24259
rect 10149 24225 10183 24259
rect 10183 24225 10192 24259
rect 10140 24216 10192 24225
rect 11520 24216 11572 24268
rect 8852 24148 8904 24200
rect 8944 24148 8996 24200
rect 12440 24148 12492 24200
rect 3332 24080 3384 24132
rect 4436 24080 4488 24132
rect 4620 24080 4672 24132
rect 5816 24080 5868 24132
rect 6184 24080 6236 24132
rect 6644 24080 6696 24132
rect 7380 24080 7432 24132
rect 8576 24080 8628 24132
rect 10140 24080 10192 24132
rect 3148 24055 3200 24064
rect 3148 24021 3157 24055
rect 3157 24021 3191 24055
rect 3191 24021 3200 24055
rect 3148 24012 3200 24021
rect 4160 24012 4212 24064
rect 4344 24012 4396 24064
rect 6000 24012 6052 24064
rect 8760 24012 8812 24064
rect 10692 24055 10744 24064
rect 10692 24021 10701 24055
rect 10701 24021 10735 24055
rect 10735 24021 10744 24055
rect 10692 24012 10744 24021
rect 11428 24012 11480 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 2780 23851 2832 23860
rect 2780 23817 2789 23851
rect 2789 23817 2823 23851
rect 2823 23817 2832 23851
rect 2780 23808 2832 23817
rect 4620 23808 4672 23860
rect 4712 23851 4764 23860
rect 4712 23817 4721 23851
rect 4721 23817 4755 23851
rect 4755 23817 4764 23851
rect 6644 23851 6696 23860
rect 4712 23808 4764 23817
rect 6644 23817 6653 23851
rect 6653 23817 6687 23851
rect 6687 23817 6696 23851
rect 6644 23808 6696 23817
rect 7104 23808 7156 23860
rect 8208 23851 8260 23860
rect 8208 23817 8217 23851
rect 8217 23817 8251 23851
rect 8251 23817 8260 23851
rect 8208 23808 8260 23817
rect 9956 23808 10008 23860
rect 10140 23851 10192 23860
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 11520 23851 11572 23860
rect 11520 23817 11529 23851
rect 11529 23817 11563 23851
rect 11563 23817 11572 23851
rect 11520 23808 11572 23817
rect 3332 23783 3384 23792
rect 3332 23749 3341 23783
rect 3341 23749 3375 23783
rect 3375 23749 3384 23783
rect 3332 23740 3384 23749
rect 6920 23740 6972 23792
rect 7380 23783 7432 23792
rect 7380 23749 7389 23783
rect 7389 23749 7423 23783
rect 7423 23749 7432 23783
rect 7380 23740 7432 23749
rect 8300 23740 8352 23792
rect 5724 23672 5776 23724
rect 7012 23672 7064 23724
rect 7472 23715 7524 23724
rect 7472 23681 7481 23715
rect 7481 23681 7515 23715
rect 7515 23681 7524 23715
rect 9312 23740 9364 23792
rect 7472 23672 7524 23681
rect 11428 23672 11480 23724
rect 12072 23740 12124 23792
rect 3240 23647 3292 23656
rect 3240 23613 3249 23647
rect 3249 23613 3283 23647
rect 3283 23613 3292 23647
rect 3240 23604 3292 23613
rect 4068 23604 4120 23656
rect 4804 23647 4856 23656
rect 4804 23613 4813 23647
rect 4813 23613 4847 23647
rect 4847 23613 4856 23647
rect 4804 23604 4856 23613
rect 5080 23604 5132 23656
rect 4712 23536 4764 23588
rect 5816 23647 5868 23656
rect 5816 23613 5825 23647
rect 5825 23613 5859 23647
rect 5859 23613 5868 23647
rect 5816 23604 5868 23613
rect 5540 23536 5592 23588
rect 7564 23604 7616 23656
rect 4896 23511 4948 23520
rect 4896 23477 4905 23511
rect 4905 23477 4939 23511
rect 4939 23477 4948 23511
rect 4896 23468 4948 23477
rect 5172 23468 5224 23520
rect 8760 23536 8812 23588
rect 10692 23536 10744 23588
rect 11520 23536 11572 23588
rect 12440 23579 12492 23588
rect 12440 23545 12449 23579
rect 12449 23545 12483 23579
rect 12483 23545 12492 23579
rect 12440 23536 12492 23545
rect 7288 23468 7340 23520
rect 9312 23468 9364 23520
rect 9680 23511 9732 23520
rect 9680 23477 9689 23511
rect 9689 23477 9723 23511
rect 9723 23477 9732 23511
rect 9680 23468 9732 23477
rect 12256 23468 12308 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 4252 23264 4304 23316
rect 4988 23264 5040 23316
rect 5448 23264 5500 23316
rect 5724 23264 5776 23316
rect 6644 23264 6696 23316
rect 7472 23307 7524 23316
rect 7472 23273 7481 23307
rect 7481 23273 7515 23307
rect 7515 23273 7524 23307
rect 7472 23264 7524 23273
rect 8852 23264 8904 23316
rect 2228 23196 2280 23248
rect 3148 23196 3200 23248
rect 3976 23196 4028 23248
rect 6920 23196 6972 23248
rect 8300 23196 8352 23248
rect 12072 23264 12124 23316
rect 12440 23264 12492 23316
rect 10416 23196 10468 23248
rect 10692 23196 10744 23248
rect 2688 23128 2740 23180
rect 3516 23060 3568 23112
rect 4528 23128 4580 23180
rect 5080 23128 5132 23180
rect 5448 23171 5500 23180
rect 5448 23137 5457 23171
rect 5457 23137 5491 23171
rect 5491 23137 5500 23171
rect 5448 23128 5500 23137
rect 5540 23128 5592 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23128 7892 23180
rect 8484 23171 8536 23180
rect 8484 23137 8493 23171
rect 8493 23137 8527 23171
rect 8527 23137 8536 23171
rect 8484 23128 8536 23137
rect 11888 23171 11940 23180
rect 5172 23060 5224 23112
rect 6000 23060 6052 23112
rect 8760 23103 8812 23112
rect 5632 22992 5684 23044
rect 8760 23069 8769 23103
rect 8769 23069 8803 23103
rect 8803 23069 8812 23103
rect 8760 23060 8812 23069
rect 11336 23060 11388 23112
rect 11152 22992 11204 23044
rect 11888 23137 11897 23171
rect 11897 23137 11931 23171
rect 11931 23137 11940 23171
rect 11888 23128 11940 23137
rect 11980 23128 12032 23180
rect 12716 23128 12768 23180
rect 12072 22924 12124 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2228 22763 2280 22772
rect 2228 22729 2237 22763
rect 2237 22729 2271 22763
rect 2271 22729 2280 22763
rect 2228 22720 2280 22729
rect 4528 22720 4580 22772
rect 4804 22763 4856 22772
rect 4804 22729 4813 22763
rect 4813 22729 4847 22763
rect 4847 22729 4856 22763
rect 4804 22720 4856 22729
rect 5540 22720 5592 22772
rect 7288 22720 7340 22772
rect 7840 22720 7892 22772
rect 9404 22720 9456 22772
rect 11980 22763 12032 22772
rect 11980 22729 11989 22763
rect 11989 22729 12023 22763
rect 12023 22729 12032 22763
rect 11980 22720 12032 22729
rect 12808 22720 12860 22772
rect 4160 22652 4212 22704
rect 4436 22652 4488 22704
rect 5448 22652 5500 22704
rect 10968 22652 11020 22704
rect 11428 22652 11480 22704
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 2872 22516 2924 22568
rect 4160 22516 4212 22568
rect 8760 22584 8812 22636
rect 11152 22627 11204 22636
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 11336 22584 11388 22636
rect 3424 22491 3476 22500
rect 3424 22457 3433 22491
rect 3433 22457 3467 22491
rect 3467 22457 3476 22491
rect 3424 22448 3476 22457
rect 2504 22423 2556 22432
rect 2504 22389 2513 22423
rect 2513 22389 2547 22423
rect 2547 22389 2556 22423
rect 2504 22380 2556 22389
rect 2872 22423 2924 22432
rect 2872 22389 2881 22423
rect 2881 22389 2915 22423
rect 2915 22389 2924 22423
rect 2872 22380 2924 22389
rect 3884 22448 3936 22500
rect 4252 22448 4304 22500
rect 4804 22448 4856 22500
rect 5356 22448 5408 22500
rect 6736 22448 6788 22500
rect 6644 22380 6696 22432
rect 8484 22423 8536 22432
rect 8484 22389 8493 22423
rect 8493 22389 8527 22423
rect 8527 22389 8536 22423
rect 8484 22380 8536 22389
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 10324 22423 10376 22432
rect 10324 22389 10333 22423
rect 10333 22389 10367 22423
rect 10367 22389 10376 22423
rect 10324 22380 10376 22389
rect 10968 22491 11020 22500
rect 10968 22457 10977 22491
rect 10977 22457 11011 22491
rect 11011 22457 11020 22491
rect 10968 22448 11020 22457
rect 12256 22448 12308 22500
rect 12900 22516 12952 22568
rect 12808 22448 12860 22500
rect 11336 22380 11388 22432
rect 11428 22380 11480 22432
rect 12072 22380 12124 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 2688 22219 2740 22228
rect 2688 22185 2697 22219
rect 2697 22185 2731 22219
rect 2731 22185 2740 22219
rect 2688 22176 2740 22185
rect 3424 22219 3476 22228
rect 3424 22185 3433 22219
rect 3433 22185 3467 22219
rect 3467 22185 3476 22219
rect 3424 22176 3476 22185
rect 4896 22176 4948 22228
rect 5356 22219 5408 22228
rect 5356 22185 5365 22219
rect 5365 22185 5399 22219
rect 5399 22185 5408 22219
rect 5356 22176 5408 22185
rect 5632 22176 5684 22228
rect 6736 22176 6788 22228
rect 7012 22219 7064 22228
rect 7012 22185 7021 22219
rect 7021 22185 7055 22219
rect 7055 22185 7064 22219
rect 7012 22176 7064 22185
rect 8760 22176 8812 22228
rect 10968 22219 11020 22228
rect 10968 22185 10977 22219
rect 10977 22185 11011 22219
rect 11011 22185 11020 22219
rect 10968 22176 11020 22185
rect 6092 22108 6144 22160
rect 6644 22151 6696 22160
rect 6644 22117 6653 22151
rect 6653 22117 6687 22151
rect 6687 22117 6696 22151
rect 6644 22108 6696 22117
rect 9404 22108 9456 22160
rect 11612 22151 11664 22160
rect 11612 22117 11621 22151
rect 11621 22117 11655 22151
rect 11655 22117 11664 22151
rect 11612 22108 11664 22117
rect 11980 22108 12032 22160
rect 13452 22108 13504 22160
rect 3332 22040 3384 22092
rect 4988 22083 5040 22092
rect 4988 22049 4997 22083
rect 4997 22049 5031 22083
rect 5031 22049 5040 22083
rect 4988 22040 5040 22049
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 10324 22040 10376 22092
rect 8116 21972 8168 22024
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 12164 21972 12216 22024
rect 13084 22015 13136 22024
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 2504 21904 2556 21956
rect 7472 21904 7524 21956
rect 12072 21947 12124 21956
rect 12072 21913 12081 21947
rect 12081 21913 12115 21947
rect 12115 21913 12124 21947
rect 12072 21904 12124 21913
rect 12532 21904 12584 21956
rect 4896 21836 4948 21888
rect 10784 21836 10836 21888
rect 11336 21879 11388 21888
rect 11336 21845 11345 21879
rect 11345 21845 11379 21879
rect 11379 21845 11388 21879
rect 11336 21836 11388 21845
rect 11980 21836 12032 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 4988 21632 5040 21684
rect 5356 21632 5408 21684
rect 9404 21675 9456 21684
rect 9404 21641 9413 21675
rect 9413 21641 9447 21675
rect 9447 21641 9456 21675
rect 9404 21632 9456 21641
rect 11612 21632 11664 21684
rect 12164 21675 12216 21684
rect 12164 21641 12173 21675
rect 12173 21641 12207 21675
rect 12207 21641 12216 21675
rect 12164 21632 12216 21641
rect 13452 21675 13504 21684
rect 13452 21641 13461 21675
rect 13461 21641 13495 21675
rect 13495 21641 13504 21675
rect 13452 21632 13504 21641
rect 4436 21564 4488 21616
rect 6828 21564 6880 21616
rect 13084 21564 13136 21616
rect 4160 21496 4212 21548
rect 4988 21539 5040 21548
rect 4988 21505 4997 21539
rect 4997 21505 5031 21539
rect 5031 21505 5040 21539
rect 4988 21496 5040 21505
rect 6736 21496 6788 21548
rect 7196 21496 7248 21548
rect 12072 21496 12124 21548
rect 13268 21496 13320 21548
rect 7380 21471 7432 21480
rect 7380 21437 7389 21471
rect 7389 21437 7423 21471
rect 7423 21437 7432 21471
rect 7380 21428 7432 21437
rect 7932 21471 7984 21480
rect 7932 21437 7941 21471
rect 7941 21437 7975 21471
rect 7975 21437 7984 21471
rect 7932 21428 7984 21437
rect 9588 21471 9640 21480
rect 3332 21292 3384 21344
rect 4896 21360 4948 21412
rect 7472 21360 7524 21412
rect 9588 21437 9597 21471
rect 9597 21437 9631 21471
rect 9631 21437 9640 21471
rect 9588 21428 9640 21437
rect 9680 21428 9732 21480
rect 8484 21360 8536 21412
rect 8668 21403 8720 21412
rect 8668 21369 8677 21403
rect 8677 21369 8711 21403
rect 8711 21369 8720 21403
rect 8668 21360 8720 21369
rect 9404 21360 9456 21412
rect 10048 21360 10100 21412
rect 12532 21403 12584 21412
rect 12532 21369 12541 21403
rect 12541 21369 12575 21403
rect 12575 21369 12584 21403
rect 12532 21360 12584 21369
rect 12624 21403 12676 21412
rect 12624 21369 12633 21403
rect 12633 21369 12667 21403
rect 12667 21369 12676 21403
rect 12624 21360 12676 21369
rect 7564 21292 7616 21344
rect 11336 21292 11388 21344
rect 12440 21292 12492 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 1400 21088 1452 21140
rect 3424 21088 3476 21140
rect 7380 21088 7432 21140
rect 7472 21131 7524 21140
rect 7472 21097 7481 21131
rect 7481 21097 7515 21131
rect 7515 21097 7524 21131
rect 7932 21131 7984 21140
rect 7472 21088 7524 21097
rect 7932 21097 7941 21131
rect 7941 21097 7975 21131
rect 7975 21097 7984 21131
rect 7932 21088 7984 21097
rect 8116 21131 8168 21140
rect 8116 21097 8125 21131
rect 8125 21097 8159 21131
rect 8159 21097 8168 21131
rect 8116 21088 8168 21097
rect 8668 21088 8720 21140
rect 10048 21131 10100 21140
rect 10048 21097 10057 21131
rect 10057 21097 10091 21131
rect 10091 21097 10100 21131
rect 10048 21088 10100 21097
rect 12624 21088 12676 21140
rect 4252 21020 4304 21072
rect 4436 21020 4488 21072
rect 9680 21020 9732 21072
rect 10784 21020 10836 21072
rect 11704 21020 11756 21072
rect 4896 20995 4948 21004
rect 4896 20961 4905 20995
rect 4905 20961 4939 20995
rect 4939 20961 4948 20995
rect 4896 20952 4948 20961
rect 6184 20952 6236 21004
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 6552 20952 6604 21004
rect 7472 20952 7524 21004
rect 8024 20995 8076 21004
rect 8024 20961 8033 20995
rect 8033 20961 8067 20995
rect 8067 20961 8076 20995
rect 8024 20952 8076 20961
rect 8484 20995 8536 21004
rect 8484 20961 8493 20995
rect 8493 20961 8527 20995
rect 8527 20961 8536 20995
rect 8484 20952 8536 20961
rect 13268 20952 13320 21004
rect 9312 20884 9364 20936
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 11152 20884 11204 20936
rect 13176 20884 13228 20936
rect 12072 20859 12124 20868
rect 12072 20825 12081 20859
rect 12081 20825 12115 20859
rect 12115 20825 12124 20859
rect 12072 20816 12124 20825
rect 9588 20748 9640 20800
rect 10048 20748 10100 20800
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 11060 20748 11112 20800
rect 11520 20748 11572 20800
rect 12532 20748 12584 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 4436 20544 4488 20596
rect 4896 20544 4948 20596
rect 5724 20587 5776 20596
rect 5724 20553 5733 20587
rect 5733 20553 5767 20587
rect 5767 20553 5776 20587
rect 5724 20544 5776 20553
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 4988 20519 5040 20528
rect 4988 20485 4997 20519
rect 4997 20485 5031 20519
rect 5031 20485 5040 20519
rect 4988 20476 5040 20485
rect 8024 20544 8076 20596
rect 9404 20544 9456 20596
rect 11704 20587 11756 20596
rect 11704 20553 11713 20587
rect 11713 20553 11747 20587
rect 11747 20553 11756 20587
rect 11704 20544 11756 20553
rect 11980 20544 12032 20596
rect 13268 20587 13320 20596
rect 13268 20553 13277 20587
rect 13277 20553 13311 20587
rect 13311 20553 13320 20587
rect 13268 20544 13320 20553
rect 13912 20587 13964 20596
rect 13912 20553 13921 20587
rect 13921 20553 13955 20587
rect 13955 20553 13964 20587
rect 13912 20544 13964 20553
rect 11152 20476 11204 20528
rect 5724 20340 5776 20392
rect 7380 20383 7432 20392
rect 7380 20349 7389 20383
rect 7389 20349 7423 20383
rect 7423 20349 7432 20383
rect 7380 20340 7432 20349
rect 8668 20408 8720 20460
rect 10968 20408 11020 20460
rect 9680 20340 9732 20392
rect 12348 20383 12400 20392
rect 4528 20315 4580 20324
rect 4528 20281 4537 20315
rect 4537 20281 4571 20315
rect 4571 20281 4580 20315
rect 4528 20272 4580 20281
rect 9404 20272 9456 20324
rect 5356 20204 5408 20256
rect 6184 20204 6236 20256
rect 12348 20349 12357 20383
rect 12357 20349 12391 20383
rect 12391 20349 12400 20383
rect 12348 20340 12400 20349
rect 12716 20340 12768 20392
rect 13912 20340 13964 20392
rect 10968 20272 11020 20324
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 112 19932 164 19984
rect 2964 19864 3016 19916
rect 4988 19932 5040 19984
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 6276 19864 6328 19916
rect 7748 20000 7800 20052
rect 8300 20000 8352 20052
rect 9680 20000 9732 20052
rect 12164 20000 12216 20052
rect 7564 19932 7616 19984
rect 10416 19975 10468 19984
rect 10416 19941 10425 19975
rect 10425 19941 10459 19975
rect 10459 19941 10468 19975
rect 10416 19932 10468 19941
rect 10876 19932 10928 19984
rect 11060 19975 11112 19984
rect 11060 19941 11069 19975
rect 11069 19941 11103 19975
rect 11103 19941 11112 19975
rect 11060 19932 11112 19941
rect 7748 19864 7800 19916
rect 8484 19864 8536 19916
rect 10232 19864 10284 19916
rect 4988 19839 5040 19848
rect 4988 19805 4997 19839
rect 4997 19805 5031 19839
rect 5031 19805 5040 19839
rect 7840 19839 7892 19848
rect 4988 19796 5040 19805
rect 6000 19728 6052 19780
rect 6828 19771 6880 19780
rect 6828 19737 6837 19771
rect 6837 19737 6871 19771
rect 6871 19737 6880 19771
rect 6828 19728 6880 19737
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 5264 19703 5316 19712
rect 5264 19669 5273 19703
rect 5273 19669 5307 19703
rect 5307 19669 5316 19703
rect 6092 19703 6144 19712
rect 5264 19660 5316 19669
rect 6092 19669 6101 19703
rect 6101 19669 6135 19703
rect 6135 19669 6144 19703
rect 6092 19660 6144 19669
rect 8668 19660 8720 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 2964 19499 3016 19508
rect 2964 19465 2973 19499
rect 2973 19465 3007 19499
rect 3007 19465 3016 19499
rect 2964 19456 3016 19465
rect 4712 19456 4764 19508
rect 10968 19499 11020 19508
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 5264 19431 5316 19440
rect 5264 19397 5273 19431
rect 5273 19397 5307 19431
rect 5307 19397 5316 19431
rect 5264 19388 5316 19397
rect 6276 19431 6328 19440
rect 6276 19397 6285 19431
rect 6285 19397 6319 19431
rect 6319 19397 6328 19431
rect 6276 19388 6328 19397
rect 6092 19320 6144 19372
rect 5172 19295 5224 19304
rect 5172 19261 5181 19295
rect 5181 19261 5215 19295
rect 5215 19261 5224 19295
rect 5172 19252 5224 19261
rect 6828 19295 6880 19304
rect 4896 19184 4948 19236
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 7748 19252 7800 19304
rect 10968 19465 10977 19499
rect 10977 19465 11011 19499
rect 11011 19465 11020 19499
rect 10968 19456 11020 19465
rect 8300 19388 8352 19440
rect 8668 19295 8720 19304
rect 8668 19261 8677 19295
rect 8677 19261 8711 19295
rect 8711 19261 8720 19295
rect 8668 19252 8720 19261
rect 9864 19252 9916 19304
rect 10232 19252 10284 19304
rect 6920 19184 6972 19236
rect 10692 19184 10744 19236
rect 5448 19116 5500 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 9312 19116 9364 19168
rect 9864 19116 9916 19168
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 4160 18912 4212 18964
rect 5816 18955 5868 18964
rect 5816 18921 5825 18955
rect 5825 18921 5859 18955
rect 5859 18921 5868 18955
rect 5816 18912 5868 18921
rect 6092 18955 6144 18964
rect 6092 18921 6101 18955
rect 6101 18921 6135 18955
rect 6135 18921 6144 18955
rect 6092 18912 6144 18921
rect 8300 18912 8352 18964
rect 6828 18844 6880 18896
rect 10416 18955 10468 18964
rect 10416 18921 10425 18955
rect 10425 18921 10459 18955
rect 10459 18921 10468 18955
rect 10416 18912 10468 18921
rect 4988 18819 5040 18828
rect 4988 18785 4997 18819
rect 4997 18785 5031 18819
rect 5031 18785 5040 18819
rect 4988 18776 5040 18785
rect 5172 18776 5224 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 6920 18776 6972 18828
rect 7380 18776 7432 18828
rect 7564 18776 7616 18828
rect 8484 18776 8536 18828
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10692 18819 10744 18828
rect 10692 18785 10701 18819
rect 10701 18785 10735 18819
rect 10735 18785 10744 18819
rect 10692 18776 10744 18785
rect 4068 18708 4120 18760
rect 6184 18708 6236 18760
rect 8208 18708 8260 18760
rect 9588 18708 9640 18760
rect 11520 18708 11572 18760
rect 4804 18683 4856 18692
rect 4804 18649 4813 18683
rect 4813 18649 4847 18683
rect 4847 18649 4856 18683
rect 4804 18640 4856 18649
rect 5448 18572 5500 18624
rect 7380 18572 7432 18624
rect 7472 18572 7524 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 8852 18368 8904 18420
rect 9404 18368 9456 18420
rect 9772 18368 9824 18420
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 4068 18300 4120 18352
rect 4804 18343 4856 18352
rect 4804 18309 4813 18343
rect 4813 18309 4847 18343
rect 4847 18309 4856 18343
rect 4804 18300 4856 18309
rect 6276 18343 6328 18352
rect 6276 18309 6285 18343
rect 6285 18309 6319 18343
rect 6319 18309 6328 18343
rect 6276 18300 6328 18309
rect 7380 18300 7432 18352
rect 7748 18300 7800 18352
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 5816 18232 5868 18284
rect 5908 18232 5960 18284
rect 9680 18232 9732 18284
rect 4804 18096 4856 18148
rect 7012 18164 7064 18216
rect 7472 18164 7524 18216
rect 7380 18139 7432 18148
rect 7380 18105 7389 18139
rect 7389 18105 7423 18139
rect 7423 18105 7432 18139
rect 8484 18164 8536 18216
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 9864 18300 9916 18352
rect 7380 18096 7432 18105
rect 4068 18028 4120 18080
rect 4528 18028 4580 18080
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5080 18028 5132 18037
rect 5816 18028 5868 18080
rect 9312 18096 9364 18148
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 6184 17824 6236 17876
rect 7012 17867 7064 17876
rect 7012 17833 7021 17867
rect 7021 17833 7055 17867
rect 7055 17833 7064 17867
rect 7012 17824 7064 17833
rect 7196 17824 7248 17876
rect 9404 17867 9456 17876
rect 9404 17833 9413 17867
rect 9413 17833 9447 17867
rect 9447 17833 9456 17867
rect 9404 17824 9456 17833
rect 9772 17824 9824 17876
rect 6920 17756 6972 17808
rect 9864 17756 9916 17808
rect 10324 17824 10376 17876
rect 11428 17824 11480 17876
rect 11520 17799 11572 17808
rect 11520 17765 11529 17799
rect 11529 17765 11563 17799
rect 11563 17765 11572 17799
rect 11520 17756 11572 17765
rect 5080 17688 5132 17740
rect 7564 17731 7616 17740
rect 7564 17697 7573 17731
rect 7573 17697 7607 17731
rect 7607 17697 7616 17731
rect 7564 17688 7616 17697
rect 7932 17731 7984 17740
rect 7932 17697 7941 17731
rect 7941 17697 7975 17731
rect 7975 17697 7984 17731
rect 7932 17688 7984 17697
rect 9588 17688 9640 17740
rect 3056 17620 3108 17672
rect 7656 17620 7708 17672
rect 8024 17663 8076 17672
rect 8024 17629 8033 17663
rect 8033 17629 8067 17663
rect 8067 17629 8076 17663
rect 8024 17620 8076 17629
rect 12808 17620 12860 17672
rect 4436 17552 4488 17604
rect 12716 17552 12768 17604
rect 4804 17527 4856 17536
rect 4804 17493 4813 17527
rect 4813 17493 4847 17527
rect 4847 17493 4856 17527
rect 4804 17484 4856 17493
rect 5724 17484 5776 17536
rect 12164 17484 12216 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 5080 17280 5132 17332
rect 7380 17323 7432 17332
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 8300 17280 8352 17332
rect 7840 17212 7892 17264
rect 4528 17144 4580 17196
rect 7932 17144 7984 17196
rect 4068 17076 4120 17128
rect 5632 17076 5684 17128
rect 7380 17076 7432 17128
rect 7656 17076 7708 17128
rect 9128 17119 9180 17128
rect 9128 17085 9137 17119
rect 9137 17085 9171 17119
rect 9171 17085 9180 17119
rect 9128 17076 9180 17085
rect 6920 17008 6972 17060
rect 9772 17280 9824 17332
rect 11520 17280 11572 17332
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 10784 17076 10836 17128
rect 10876 17119 10928 17128
rect 10876 17085 10920 17119
rect 10920 17085 10928 17119
rect 10876 17076 10928 17085
rect 12256 17076 12308 17128
rect 12072 17008 12124 17060
rect 12532 17051 12584 17060
rect 12532 17017 12541 17051
rect 12541 17017 12575 17051
rect 12575 17017 12584 17051
rect 12532 17008 12584 17017
rect 3976 16940 4028 16992
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 7564 16940 7616 16992
rect 11244 16940 11296 16992
rect 12164 16940 12216 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 4896 16736 4948 16788
rect 3056 16600 3108 16652
rect 7288 16736 7340 16788
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 9588 16736 9640 16788
rect 11428 16736 11480 16788
rect 6736 16600 6788 16652
rect 8300 16668 8352 16720
rect 10692 16711 10744 16720
rect 10692 16677 10701 16711
rect 10701 16677 10735 16711
rect 10735 16677 10744 16711
rect 10692 16668 10744 16677
rect 10784 16668 10836 16720
rect 12164 16668 12216 16720
rect 12808 16711 12860 16720
rect 12808 16677 12817 16711
rect 12817 16677 12851 16711
rect 12851 16677 12860 16711
rect 12808 16668 12860 16677
rect 7380 16600 7432 16652
rect 8024 16600 8076 16652
rect 5448 16575 5500 16584
rect 5448 16541 5457 16575
rect 5457 16541 5491 16575
rect 5491 16541 5500 16575
rect 5448 16532 5500 16541
rect 9680 16532 9732 16584
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 11060 16575 11112 16584
rect 11060 16541 11069 16575
rect 11069 16541 11103 16575
rect 11103 16541 11112 16575
rect 11060 16532 11112 16541
rect 12900 16532 12952 16584
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 3148 16396 3200 16405
rect 4804 16396 4856 16448
rect 5540 16396 5592 16448
rect 5908 16396 5960 16448
rect 7656 16396 7708 16448
rect 9312 16396 9364 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 7380 16235 7432 16244
rect 7380 16201 7389 16235
rect 7389 16201 7423 16235
rect 7423 16201 7432 16235
rect 7380 16192 7432 16201
rect 8300 16192 8352 16244
rect 8852 16192 8904 16244
rect 6736 16124 6788 16176
rect 7840 16124 7892 16176
rect 8116 16124 8168 16176
rect 10600 16192 10652 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 14740 16192 14792 16244
rect 12900 16167 12952 16176
rect 5448 16056 5500 16108
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 3976 15988 4028 16040
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 4896 15988 4948 16040
rect 5540 16031 5592 16040
rect 5540 15997 5549 16031
rect 5549 15997 5583 16031
rect 5583 15997 5592 16031
rect 5540 15988 5592 15997
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 5816 15963 5868 15972
rect 5816 15929 5825 15963
rect 5825 15929 5859 15963
rect 5859 15929 5868 15963
rect 5816 15920 5868 15929
rect 7380 15920 7432 15972
rect 8300 15963 8352 15972
rect 8300 15929 8309 15963
rect 8309 15929 8343 15963
rect 8343 15929 8352 15963
rect 8300 15920 8352 15929
rect 12900 16133 12909 16167
rect 12909 16133 12943 16167
rect 12943 16133 12952 16167
rect 12900 16124 12952 16133
rect 9496 16056 9548 16108
rect 9772 16056 9824 16108
rect 12808 15988 12860 16040
rect 9956 15920 10008 15972
rect 5632 15852 5684 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 4896 15648 4948 15700
rect 5264 15648 5316 15700
rect 6184 15648 6236 15700
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 7840 15648 7892 15700
rect 8024 15648 8076 15700
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 9956 15648 10008 15700
rect 10600 15648 10652 15700
rect 5264 15512 5316 15564
rect 11244 15580 11296 15632
rect 11704 15580 11756 15632
rect 6736 15512 6788 15564
rect 8024 15512 8076 15564
rect 8208 15512 8260 15564
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 5816 15444 5868 15496
rect 3056 15376 3108 15428
rect 7840 15376 7892 15428
rect 12072 15419 12124 15428
rect 12072 15385 12081 15419
rect 12081 15385 12115 15419
rect 12115 15385 12124 15419
rect 12072 15376 12124 15385
rect 6092 15351 6144 15360
rect 6092 15317 6101 15351
rect 6101 15317 6135 15351
rect 6135 15317 6144 15351
rect 6092 15308 6144 15317
rect 10600 15351 10652 15360
rect 10600 15317 10609 15351
rect 10609 15317 10643 15351
rect 10643 15317 10652 15351
rect 10600 15308 10652 15317
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 12716 15308 12768 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 8208 15104 8260 15156
rect 8852 15147 8904 15156
rect 8852 15113 8861 15147
rect 8861 15113 8895 15147
rect 8895 15113 8904 15147
rect 8852 15104 8904 15113
rect 9956 15104 10008 15156
rect 10600 15147 10652 15156
rect 10600 15113 10609 15147
rect 10609 15113 10643 15147
rect 10643 15113 10652 15147
rect 10600 15104 10652 15113
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 3148 15036 3200 15088
rect 4896 15036 4948 15088
rect 10876 15036 10928 15088
rect 11152 15036 11204 15088
rect 12992 15079 13044 15088
rect 12992 15045 13001 15079
rect 13001 15045 13035 15079
rect 13035 15045 13044 15079
rect 12992 15036 13044 15045
rect 4804 14968 4856 15020
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 8300 14968 8352 15020
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 10968 14968 11020 15020
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5264 14900 5316 14909
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 8024 14900 8076 14952
rect 12900 14900 12952 14952
rect 13360 14900 13412 14952
rect 6184 14832 6236 14884
rect 7656 14832 7708 14884
rect 8852 14832 8904 14884
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 10600 14764 10652 14816
rect 11060 14832 11112 14884
rect 11980 14764 12032 14816
rect 13544 14764 13596 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 5264 14560 5316 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 6736 14560 6788 14612
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 9680 14560 9732 14612
rect 11244 14560 11296 14612
rect 6644 14492 6696 14544
rect 7748 14492 7800 14544
rect 4896 14467 4948 14476
rect 4896 14433 4905 14467
rect 4905 14433 4939 14467
rect 4939 14433 4948 14467
rect 4896 14424 4948 14433
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 9864 14492 9916 14544
rect 11152 14492 11204 14544
rect 8852 14424 8904 14476
rect 11060 14467 11112 14476
rect 11060 14433 11069 14467
rect 11069 14433 11103 14467
rect 11103 14433 11112 14467
rect 11060 14424 11112 14433
rect 6184 14356 6236 14408
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 11612 14356 11664 14408
rect 12716 14356 12768 14408
rect 8300 14288 8352 14340
rect 10508 14288 10560 14340
rect 10876 14288 10928 14340
rect 12072 14288 12124 14340
rect 4344 14220 4396 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 6184 14016 6236 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 7932 14059 7984 14068
rect 7932 14025 7941 14059
rect 7941 14025 7975 14059
rect 7975 14025 7984 14059
rect 7932 14016 7984 14025
rect 8116 14016 8168 14068
rect 10600 14016 10652 14068
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 11612 14059 11664 14068
rect 11612 14025 11621 14059
rect 11621 14025 11655 14059
rect 11655 14025 11664 14059
rect 11612 14016 11664 14025
rect 11980 14016 12032 14068
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 5264 13880 5316 13932
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 8116 13812 8168 13864
rect 4436 13744 4488 13796
rect 4896 13744 4948 13796
rect 5632 13744 5684 13796
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 5356 13676 5408 13728
rect 6644 13744 6696 13796
rect 10232 13787 10284 13796
rect 10232 13753 10241 13787
rect 10241 13753 10275 13787
rect 10275 13753 10284 13787
rect 10232 13744 10284 13753
rect 10600 13744 10652 13796
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 4068 13404 4120 13456
rect 5356 13404 5408 13456
rect 6092 13472 6144 13524
rect 6184 13472 6236 13524
rect 6920 13472 6972 13524
rect 8760 13472 8812 13524
rect 7932 13447 7984 13456
rect 7932 13413 7941 13447
rect 7941 13413 7975 13447
rect 7975 13413 7984 13447
rect 7932 13404 7984 13413
rect 9864 13447 9916 13456
rect 9864 13413 9873 13447
rect 9873 13413 9907 13447
rect 9907 13413 9916 13447
rect 9864 13404 9916 13413
rect 10232 13472 10284 13524
rect 11980 13336 12032 13388
rect 4344 13268 4396 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 5172 13268 5224 13320
rect 8668 13268 8720 13320
rect 10876 13268 10928 13320
rect 6368 13243 6420 13252
rect 6368 13209 6377 13243
rect 6377 13209 6411 13243
rect 6411 13209 6420 13243
rect 6368 13200 6420 13209
rect 6644 13200 6696 13252
rect 8116 13200 8168 13252
rect 10508 13200 10560 13252
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 7932 13132 7984 13184
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 4344 12928 4396 12980
rect 6092 12928 6144 12980
rect 7932 12928 7984 12980
rect 8668 12928 8720 12980
rect 10876 12971 10928 12980
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 4068 12903 4120 12912
rect 4068 12869 4077 12903
rect 4077 12869 4111 12903
rect 4111 12869 4120 12903
rect 4068 12860 4120 12869
rect 5172 12860 5224 12912
rect 8024 12792 8076 12844
rect 4712 12724 4764 12776
rect 5264 12699 5316 12708
rect 5264 12665 5273 12699
rect 5273 12665 5307 12699
rect 5307 12665 5316 12699
rect 5264 12656 5316 12665
rect 5356 12699 5408 12708
rect 5356 12665 5365 12699
rect 5365 12665 5399 12699
rect 5399 12665 5408 12699
rect 5356 12656 5408 12665
rect 6368 12656 6420 12708
rect 7380 12656 7432 12708
rect 7932 12656 7984 12708
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 8208 12588 8260 12640
rect 9864 12860 9916 12912
rect 9680 12792 9732 12844
rect 9772 12792 9824 12844
rect 13452 12792 13504 12844
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 9496 12588 9548 12640
rect 9680 12699 9732 12708
rect 9680 12665 9689 12699
rect 9689 12665 9723 12699
rect 9723 12665 9732 12699
rect 10232 12699 10284 12708
rect 9680 12656 9732 12665
rect 10232 12665 10241 12699
rect 10241 12665 10275 12699
rect 10275 12665 10284 12699
rect 10232 12656 10284 12665
rect 11336 12588 11388 12640
rect 11980 12631 12032 12640
rect 11980 12597 11989 12631
rect 11989 12597 12023 12631
rect 12023 12597 12032 12631
rect 11980 12588 12032 12597
rect 12624 12588 12676 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 5172 12384 5224 12436
rect 5264 12384 5316 12436
rect 7932 12384 7984 12436
rect 6092 12359 6144 12368
rect 6092 12325 6101 12359
rect 6101 12325 6135 12359
rect 6135 12325 6144 12359
rect 6092 12316 6144 12325
rect 7288 12316 7340 12368
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 8576 12316 8628 12368
rect 9588 12316 9640 12368
rect 11336 12359 11388 12368
rect 11336 12325 11345 12359
rect 11345 12325 11379 12359
rect 11379 12325 11388 12359
rect 11336 12316 11388 12325
rect 11980 12316 12032 12368
rect 13268 12248 13320 12300
rect 6092 12180 6144 12232
rect 4896 12112 4948 12164
rect 6736 12180 6788 12232
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 10232 12112 10284 12164
rect 10508 12112 10560 12164
rect 4988 12044 5040 12096
rect 5448 12044 5500 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 5540 11840 5592 11892
rect 5908 11840 5960 11892
rect 6184 11840 6236 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 7932 11840 7984 11892
rect 8668 11883 8720 11892
rect 8668 11849 8677 11883
rect 8677 11849 8711 11883
rect 8711 11849 8720 11883
rect 8668 11840 8720 11849
rect 9680 11840 9732 11892
rect 11336 11840 11388 11892
rect 11980 11840 12032 11892
rect 12992 11883 13044 11892
rect 12992 11849 13001 11883
rect 13001 11849 13035 11883
rect 13035 11849 13044 11883
rect 12992 11840 13044 11849
rect 9588 11815 9640 11824
rect 9588 11781 9597 11815
rect 9597 11781 9631 11815
rect 9631 11781 9640 11815
rect 9588 11772 9640 11781
rect 13268 11815 13320 11824
rect 13268 11781 13277 11815
rect 13277 11781 13311 11815
rect 13311 11781 13320 11815
rect 13268 11772 13320 11781
rect 6276 11747 6328 11756
rect 6276 11713 6285 11747
rect 6285 11713 6319 11747
rect 6319 11713 6328 11747
rect 6276 11704 6328 11713
rect 9128 11704 9180 11756
rect 10508 11704 10560 11756
rect 10876 11704 10928 11756
rect 5816 11679 5868 11688
rect 5816 11645 5834 11679
rect 5834 11645 5868 11679
rect 5816 11636 5868 11645
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 11152 11636 11204 11688
rect 12164 11636 12216 11688
rect 12992 11636 13044 11688
rect 4988 11568 5040 11620
rect 7288 11568 7340 11620
rect 7932 11568 7984 11620
rect 9312 11568 9364 11620
rect 6092 11500 6144 11552
rect 8852 11500 8904 11552
rect 9404 11500 9456 11552
rect 10416 11611 10468 11620
rect 10416 11577 10425 11611
rect 10425 11577 10459 11611
rect 10459 11577 10468 11611
rect 10416 11568 10468 11577
rect 10784 11500 10836 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 6736 11296 6788 11348
rect 8852 11296 8904 11348
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 9772 11296 9824 11348
rect 12072 11296 12124 11348
rect 4068 11092 4120 11144
rect 4804 11160 4856 11212
rect 5908 11160 5960 11212
rect 7748 11228 7800 11280
rect 7932 11228 7984 11280
rect 9864 11271 9916 11280
rect 9864 11237 9873 11271
rect 9873 11237 9907 11271
rect 9907 11237 9916 11271
rect 9864 11228 9916 11237
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 6644 11160 6696 11212
rect 6828 11203 6880 11212
rect 6828 11169 6837 11203
rect 6837 11169 6871 11203
rect 6871 11169 6880 11203
rect 6828 11160 6880 11169
rect 12624 11160 12676 11212
rect 8208 11092 8260 11144
rect 10232 11092 10284 11144
rect 11428 11092 11480 11144
rect 8116 11024 8168 11076
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 4068 10795 4120 10804
rect 4068 10761 4077 10795
rect 4077 10761 4111 10795
rect 4111 10761 4120 10795
rect 4068 10752 4120 10761
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 7932 10795 7984 10804
rect 7932 10761 7941 10795
rect 7941 10761 7975 10795
rect 7975 10761 7984 10795
rect 7932 10752 7984 10761
rect 8760 10752 8812 10804
rect 9864 10752 9916 10804
rect 11428 10795 11480 10804
rect 11428 10761 11437 10795
rect 11437 10761 11471 10795
rect 11471 10761 11480 10795
rect 11428 10752 11480 10761
rect 10784 10684 10836 10736
rect 4344 10616 4396 10668
rect 7656 10616 7708 10668
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 5264 10523 5316 10532
rect 5264 10489 5273 10523
rect 5273 10489 5307 10523
rect 5307 10489 5316 10523
rect 5264 10480 5316 10489
rect 5724 10480 5776 10532
rect 6736 10480 6788 10532
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7012 10480 7064 10489
rect 8668 10523 8720 10532
rect 8668 10489 8677 10523
rect 8677 10489 8711 10523
rect 8711 10489 8720 10523
rect 8668 10480 8720 10489
rect 10140 10523 10192 10532
rect 10140 10489 10149 10523
rect 10149 10489 10183 10523
rect 10183 10489 10192 10523
rect 10140 10480 10192 10489
rect 6644 10412 6696 10464
rect 10600 10412 10652 10464
rect 12624 10455 12676 10464
rect 12624 10421 12633 10455
rect 12633 10421 12667 10455
rect 12667 10421 12676 10455
rect 12624 10412 12676 10421
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 5356 10208 5408 10260
rect 6828 10251 6880 10260
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 7932 10208 7984 10260
rect 5908 10183 5960 10192
rect 5908 10149 5911 10183
rect 5911 10149 5945 10183
rect 5945 10149 5960 10183
rect 5908 10140 5960 10149
rect 7472 10183 7524 10192
rect 7472 10149 7481 10183
rect 7481 10149 7515 10183
rect 7515 10149 7524 10183
rect 7472 10140 7524 10149
rect 8208 10208 8260 10260
rect 8576 10208 8628 10260
rect 10600 10251 10652 10260
rect 10600 10217 10609 10251
rect 10609 10217 10643 10251
rect 10643 10217 10652 10251
rect 10600 10208 10652 10217
rect 9772 10140 9824 10192
rect 10140 10140 10192 10192
rect 3516 10072 3568 10124
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 7012 10072 7064 10124
rect 6920 10004 6972 10056
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 4436 9936 4488 9988
rect 6828 9936 6880 9988
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 6644 9664 6696 9716
rect 9772 9707 9824 9716
rect 7472 9596 7524 9648
rect 5448 9460 5500 9512
rect 7012 9460 7064 9512
rect 7564 9528 7616 9580
rect 8392 9503 8444 9512
rect 6092 9392 6144 9444
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 9772 9673 9781 9707
rect 9781 9673 9815 9707
rect 9815 9673 9824 9707
rect 9772 9664 9824 9673
rect 9680 9528 9732 9580
rect 10416 9503 10468 9512
rect 9588 9392 9640 9444
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 5908 9324 5960 9376
rect 6644 9324 6696 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 4712 9120 4764 9172
rect 5264 9120 5316 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 6920 9120 6972 9172
rect 7104 9120 7156 9172
rect 6644 9052 6696 9104
rect 7932 9052 7984 9104
rect 8392 9095 8444 9104
rect 8392 9061 8401 9095
rect 8401 9061 8435 9095
rect 8435 9061 8444 9095
rect 8392 9052 8444 9061
rect 9496 9120 9548 9172
rect 4344 9027 4396 9036
rect 4344 8993 4353 9027
rect 4353 8993 4387 9027
rect 4387 8993 4396 9027
rect 4344 8984 4396 8993
rect 5540 9027 5592 9036
rect 5540 8993 5549 9027
rect 5549 8993 5583 9027
rect 5583 8993 5592 9027
rect 5540 8984 5592 8993
rect 4896 8916 4948 8968
rect 6092 8984 6144 9036
rect 7012 8984 7064 9036
rect 8484 8984 8536 9036
rect 9680 9027 9732 9036
rect 9680 8993 9724 9027
rect 9724 8993 9732 9027
rect 9680 8984 9732 8993
rect 10784 8984 10836 9036
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 7196 8916 7248 8968
rect 8208 8916 8260 8968
rect 10416 8916 10468 8968
rect 5172 8848 5224 8900
rect 10232 8891 10284 8900
rect 10232 8857 10241 8891
rect 10241 8857 10275 8891
rect 10275 8857 10284 8891
rect 10232 8848 10284 8857
rect 112 8780 164 8832
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4344 8619 4396 8628
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 4804 8576 4856 8628
rect 4896 8508 4948 8560
rect 5540 8576 5592 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 7932 8508 7984 8560
rect 7104 8440 7156 8492
rect 5264 8372 5316 8424
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 8852 8440 8904 8492
rect 9312 8440 9364 8492
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 8852 8304 8904 8356
rect 7196 8279 7248 8288
rect 7196 8245 7205 8279
rect 7205 8245 7239 8279
rect 7239 8245 7248 8279
rect 7196 8236 7248 8245
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 7012 8032 7064 8084
rect 4528 7896 4580 7948
rect 6736 7964 6788 8016
rect 8116 8007 8168 8016
rect 8116 7973 8125 8007
rect 8125 7973 8159 8007
rect 8159 7973 8168 8007
rect 8116 7964 8168 7973
rect 9772 7964 9824 8016
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 9588 7896 9640 7948
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 5816 7692 5868 7744
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7564 7828 7616 7880
rect 8760 7828 8812 7880
rect 10324 7828 10376 7880
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 5264 7488 5316 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 9588 7488 9640 7540
rect 9772 7420 9824 7472
rect 12348 7420 12400 7472
rect 5540 7352 5592 7404
rect 7012 7352 7064 7404
rect 8852 7352 8904 7404
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5172 7284 5224 7293
rect 5264 7284 5316 7336
rect 8760 7284 8812 7336
rect 5908 7259 5960 7268
rect 5908 7225 5917 7259
rect 5917 7225 5951 7259
rect 5951 7225 5960 7259
rect 5908 7216 5960 7225
rect 6736 7216 6788 7268
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 8116 7216 8168 7268
rect 9772 7216 9824 7268
rect 6644 7148 6696 7157
rect 7564 7148 7616 7200
rect 10140 7191 10192 7200
rect 10140 7157 10149 7191
rect 10149 7157 10183 7191
rect 10183 7157 10192 7191
rect 10140 7148 10192 7157
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 5816 6944 5868 6996
rect 5908 6944 5960 6996
rect 8116 6987 8168 6996
rect 5264 6919 5316 6928
rect 5264 6885 5273 6919
rect 5273 6885 5307 6919
rect 5307 6885 5316 6919
rect 5264 6876 5316 6885
rect 6644 6876 6696 6928
rect 7012 6919 7064 6928
rect 7012 6885 7021 6919
rect 7021 6885 7055 6919
rect 7055 6885 7064 6919
rect 7012 6876 7064 6885
rect 4620 6808 4672 6860
rect 5172 6808 5224 6860
rect 8116 6953 8125 6987
rect 8125 6953 8159 6987
rect 8159 6953 8168 6987
rect 8116 6944 8168 6953
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 11428 6944 11480 6996
rect 9772 6876 9824 6928
rect 10140 6876 10192 6928
rect 10416 6876 10468 6928
rect 9864 6808 9916 6860
rect 6092 6740 6144 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 7012 6604 7064 6656
rect 8760 6604 8812 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 4620 6400 4672 6452
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 7196 6400 7248 6452
rect 9772 6443 9824 6452
rect 8116 6332 8168 6384
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 11428 6443 11480 6452
rect 11428 6409 11437 6443
rect 11437 6409 11471 6443
rect 11471 6409 11480 6443
rect 11428 6400 11480 6409
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 3332 6196 3384 6248
rect 6184 6196 6236 6248
rect 6920 6171 6972 6180
rect 6920 6137 6929 6171
rect 6929 6137 6963 6171
rect 6963 6137 6972 6171
rect 6920 6128 6972 6137
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7564 6171 7616 6180
rect 7012 6128 7064 6137
rect 7564 6137 7573 6171
rect 7573 6137 7607 6171
rect 7607 6137 7616 6171
rect 7564 6128 7616 6137
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 8760 6128 8812 6137
rect 10416 6171 10468 6180
rect 10416 6137 10425 6171
rect 10425 6137 10459 6171
rect 10459 6137 10468 6171
rect 10968 6171 11020 6180
rect 10416 6128 10468 6137
rect 10968 6137 10977 6171
rect 10977 6137 11011 6171
rect 11011 6137 11020 6171
rect 10968 6128 11020 6137
rect 6092 6060 6144 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 11060 6060 11112 6112
rect 11520 6060 11572 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 6920 5856 6972 5908
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 5264 5788 5316 5840
rect 7012 5831 7064 5840
rect 5632 5720 5684 5772
rect 7012 5797 7021 5831
rect 7021 5797 7055 5831
rect 7055 5797 7064 5831
rect 7012 5788 7064 5797
rect 7104 5788 7156 5840
rect 8024 5788 8076 5840
rect 8944 5788 8996 5840
rect 10600 5788 10652 5840
rect 6552 5720 6604 5772
rect 10968 5720 11020 5772
rect 11980 5720 12032 5772
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 13636 5516 13688 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 8024 5312 8076 5364
rect 6828 5244 6880 5296
rect 7288 5244 7340 5296
rect 8852 5176 8904 5228
rect 9312 5312 9364 5364
rect 10140 5312 10192 5364
rect 11980 5312 12032 5364
rect 12532 5312 12584 5364
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 8576 5108 8628 5160
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 10600 5176 10652 5228
rect 8392 5083 8444 5092
rect 8392 5049 8401 5083
rect 8401 5049 8435 5083
rect 8435 5049 8444 5083
rect 8392 5040 8444 5049
rect 11336 5108 11388 5160
rect 7748 4972 7800 5024
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 11152 4972 11204 5024
rect 11520 5040 11572 5092
rect 13360 4972 13412 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 5172 4768 5224 4820
rect 5356 4768 5408 4820
rect 7656 4811 7708 4820
rect 6184 4700 6236 4752
rect 5908 4632 5960 4684
rect 7656 4777 7665 4811
rect 7665 4777 7699 4811
rect 7699 4777 7708 4811
rect 7656 4768 7708 4777
rect 7840 4768 7892 4820
rect 9404 4768 9456 4820
rect 9680 4768 9732 4820
rect 9772 4700 9824 4752
rect 8116 4632 8168 4684
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 11336 4632 11388 4684
rect 12348 4675 12400 4684
rect 12348 4641 12357 4675
rect 12357 4641 12391 4675
rect 12391 4641 12400 4675
rect 12348 4632 12400 4641
rect 13452 4675 13504 4684
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 9404 4564 9456 4616
rect 10140 4607 10192 4616
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 7748 4496 7800 4548
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10784 4496 10836 4548
rect 13912 4496 13964 4548
rect 6184 4428 6236 4480
rect 12256 4428 12308 4480
rect 14188 4428 14240 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 5264 4224 5316 4276
rect 6000 4224 6052 4276
rect 6276 4224 6328 4276
rect 8576 4224 8628 4276
rect 11336 4267 11388 4276
rect 11336 4233 11345 4267
rect 11345 4233 11379 4267
rect 11379 4233 11388 4267
rect 11336 4224 11388 4233
rect 12348 4224 12400 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 4620 4199 4672 4208
rect 4620 4165 4629 4199
rect 4629 4165 4663 4199
rect 4663 4165 4672 4199
rect 4620 4156 4672 4165
rect 8116 4156 8168 4208
rect 9772 4156 9824 4208
rect 10416 4156 10468 4208
rect 11060 4156 11112 4208
rect 6276 4131 6328 4140
rect 6276 4097 6285 4131
rect 6285 4097 6319 4131
rect 6319 4097 6328 4131
rect 6276 4088 6328 4097
rect 6644 4088 6696 4140
rect 7564 4088 7616 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 4620 4020 4672 4072
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 5264 4020 5316 4072
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 6000 3952 6052 4004
rect 6920 3995 6972 4004
rect 6920 3961 6929 3995
rect 6929 3961 6963 3995
rect 6963 3961 6972 3995
rect 6920 3952 6972 3961
rect 8852 4088 8904 4140
rect 10876 4020 10928 4072
rect 11244 4020 11296 4072
rect 11704 4020 11756 4072
rect 13820 4020 13872 4072
rect 6092 3884 6144 3936
rect 6736 3884 6788 3936
rect 9588 3884 9640 3936
rect 10692 3884 10744 3936
rect 12716 3884 12768 3936
rect 13084 3884 13136 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 4068 3544 4120 3596
rect 7840 3680 7892 3732
rect 8392 3680 8444 3732
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 10508 3680 10560 3732
rect 11520 3680 11572 3732
rect 5264 3612 5316 3664
rect 6276 3655 6328 3664
rect 6276 3621 6279 3655
rect 6279 3621 6313 3655
rect 6313 3621 6328 3655
rect 6276 3612 6328 3621
rect 8208 3612 8260 3664
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 11428 3655 11480 3664
rect 9864 3612 9916 3621
rect 11428 3621 11437 3655
rect 11437 3621 11471 3655
rect 11471 3621 11480 3655
rect 11428 3612 11480 3621
rect 4988 3544 5040 3596
rect 6828 3544 6880 3596
rect 8024 3544 8076 3596
rect 9312 3544 9364 3596
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 13360 3544 13412 3596
rect 6000 3476 6052 3528
rect 10416 3519 10468 3528
rect 5356 3408 5408 3460
rect 6184 3408 6236 3460
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 6552 3340 6604 3392
rect 6920 3340 6972 3392
rect 9772 3340 9824 3392
rect 10140 3340 10192 3392
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 11796 3476 11848 3528
rect 13084 3476 13136 3528
rect 10324 3408 10376 3460
rect 11244 3408 11296 3460
rect 11152 3340 11204 3392
rect 15568 3340 15620 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 4068 3179 4120 3188
rect 4068 3145 4077 3179
rect 4077 3145 4111 3179
rect 4111 3145 4120 3179
rect 4068 3136 4120 3145
rect 4988 3179 5040 3188
rect 4988 3145 4997 3179
rect 4997 3145 5031 3179
rect 5031 3145 5040 3179
rect 4988 3136 5040 3145
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 8208 3136 8260 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12992 3179 13044 3188
rect 12992 3145 13001 3179
rect 13001 3145 13035 3179
rect 13035 3145 13044 3179
rect 12992 3136 13044 3145
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 664 3068 716 3120
rect 6552 3068 6604 3120
rect 6736 3068 6788 3120
rect 8300 3068 8352 3120
rect 11520 3068 11572 3120
rect 4528 3000 4580 3052
rect 5724 3000 5776 3052
rect 6644 3000 6696 3052
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 9404 3000 9456 3052
rect 10416 3000 10468 3052
rect 10784 3000 10836 3052
rect 4620 2864 4672 2916
rect 3516 2796 3568 2848
rect 12992 2932 13044 2984
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 8208 2864 8260 2916
rect 10416 2907 10468 2916
rect 10416 2873 10425 2907
rect 10425 2873 10459 2907
rect 10459 2873 10468 2907
rect 10416 2864 10468 2873
rect 8300 2796 8352 2848
rect 10140 2796 10192 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 6000 2592 6052 2644
rect 6736 2635 6788 2644
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 8024 2635 8076 2644
rect 6736 2592 6788 2601
rect 3516 2524 3568 2576
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 1584 2456 1636 2508
rect 3424 2456 3476 2508
rect 4252 2320 4304 2372
rect 7748 2567 7800 2576
rect 7748 2533 7757 2567
rect 7757 2533 7791 2567
rect 7791 2533 7800 2567
rect 7748 2524 7800 2533
rect 10324 2592 10376 2644
rect 11244 2524 11296 2576
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 11152 2499 11204 2508
rect 11152 2465 11161 2499
rect 11161 2465 11195 2499
rect 11195 2465 11204 2499
rect 11152 2456 11204 2465
rect 11336 2499 11388 2508
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 7564 2320 7616 2372
rect 6092 2252 6144 2304
rect 8668 2252 8720 2304
rect 9864 2252 9916 2304
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 2872 76 2924 128
rect 5080 76 5132 128
<< metal2 >>
rect 294 39636 350 40000
rect 846 39658 902 40000
rect 294 39584 296 39636
rect 348 39584 350 39636
rect 294 39520 350 39584
rect 768 39630 902 39658
rect 1490 39658 1546 40000
rect 768 34542 796 39630
rect 846 39520 902 39630
rect 1400 39636 1452 39642
rect 1400 39578 1452 39584
rect 1490 39630 1808 39658
rect 756 34536 808 34542
rect 756 34478 808 34484
rect 570 33144 626 33153
rect 570 33079 626 33088
rect 584 31958 612 33079
rect 572 31952 624 31958
rect 572 31894 624 31900
rect 1412 21146 1440 39578
rect 1490 39520 1546 39630
rect 1492 39024 1544 39030
rect 1492 38966 1544 38972
rect 1504 27577 1532 38966
rect 1780 35290 1808 39630
rect 2134 39636 2190 40000
rect 2686 39658 2742 40000
rect 2134 39584 2136 39636
rect 2188 39584 2190 39636
rect 2134 39520 2190 39584
rect 2424 39630 2742 39658
rect 2424 39030 2452 39630
rect 2686 39520 2742 39630
rect 3330 39658 3386 40000
rect 3974 39658 4030 40000
rect 4526 39658 4582 40000
rect 5170 39658 5226 40000
rect 3330 39630 3556 39658
rect 3330 39520 3386 39630
rect 3424 39568 3476 39574
rect 3424 39510 3476 39516
rect 2412 39024 2464 39030
rect 2412 38966 2464 38972
rect 3056 36712 3108 36718
rect 3056 36654 3108 36660
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 3068 29646 3096 36654
rect 3056 29640 3108 29646
rect 3056 29582 3108 29588
rect 3068 28966 3096 29582
rect 3056 28960 3108 28966
rect 3056 28902 3108 28908
rect 1490 27568 1546 27577
rect 1490 27503 1546 27512
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2792 23866 2820 24210
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2228 23248 2280 23254
rect 2228 23190 2280 23196
rect 2240 22778 2268 23190
rect 2688 23180 2740 23186
rect 2688 23122 2740 23128
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2504 22432 2556 22438
rect 2504 22374 2556 22380
rect 2516 21962 2544 22374
rect 2700 22234 2728 23122
rect 2872 22568 2924 22574
rect 2870 22536 2872 22545
rect 2924 22536 2926 22545
rect 2870 22471 2926 22480
rect 2884 22438 2912 22471
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2504 21956 2556 21962
rect 2504 21898 2556 21904
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 110 20088 166 20097
rect 110 20023 166 20032
rect 124 19990 152 20023
rect 112 19984 164 19990
rect 112 19926 164 19932
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2976 19514 3004 19858
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 3068 18578 3096 28902
rect 3436 28665 3464 39510
rect 3528 34066 3556 39630
rect 3974 39630 4292 39658
rect 3974 39520 4030 39630
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3516 34060 3568 34066
rect 3516 34002 3568 34008
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 4080 33114 4108 33390
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 4080 32042 4108 33050
rect 4264 32978 4292 39630
rect 4526 39630 4936 39658
rect 4526 39520 4582 39630
rect 4344 34536 4396 34542
rect 4344 34478 4396 34484
rect 4252 32972 4304 32978
rect 4252 32914 4304 32920
rect 4252 32360 4304 32366
rect 4252 32302 4304 32308
rect 4080 32014 4200 32042
rect 3976 31884 4028 31890
rect 3976 31826 4028 31832
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3988 31210 4016 31826
rect 4172 31686 4200 32014
rect 4160 31680 4212 31686
rect 4160 31622 4212 31628
rect 3976 31204 4028 31210
rect 3976 31146 4028 31152
rect 3976 30728 4028 30734
rect 3976 30670 4028 30676
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3988 30394 4016 30670
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4068 29776 4120 29782
rect 4068 29718 4120 29724
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 4080 28694 4108 29718
rect 4264 29306 4292 32302
rect 4252 29300 4304 29306
rect 4252 29242 4304 29248
rect 4068 28688 4120 28694
rect 3422 28656 3478 28665
rect 4068 28630 4120 28636
rect 3422 28591 3478 28600
rect 3148 24608 3200 24614
rect 3148 24550 3200 24556
rect 3160 24070 3188 24550
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3148 24064 3200 24070
rect 3148 24006 3200 24012
rect 3160 23254 3188 24006
rect 3344 23798 3372 24074
rect 3332 23792 3384 23798
rect 3238 23760 3294 23769
rect 3332 23734 3384 23740
rect 3238 23695 3294 23704
rect 3252 23662 3280 23695
rect 3240 23656 3292 23662
rect 3240 23598 3292 23604
rect 3436 23474 3464 28591
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 4068 28144 4120 28150
rect 4068 28086 4120 28092
rect 3976 28008 4028 28014
rect 3976 27950 4028 27956
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3988 24750 4016 27950
rect 4080 27538 4108 28086
rect 4068 27532 4120 27538
rect 4068 27474 4120 27480
rect 4160 27532 4212 27538
rect 4160 27474 4212 27480
rect 4080 26518 4108 27474
rect 4172 27130 4200 27474
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4264 27010 4292 29242
rect 4356 28966 4384 34478
rect 4804 34060 4856 34066
rect 4804 34002 4856 34008
rect 4816 33318 4844 34002
rect 4804 33312 4856 33318
rect 4804 33254 4856 33260
rect 4528 32224 4580 32230
rect 4528 32166 4580 32172
rect 4540 31822 4568 32166
rect 4528 31816 4580 31822
rect 4528 31758 4580 31764
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4632 29238 4660 29582
rect 4620 29232 4672 29238
rect 4816 29209 4844 33254
rect 4908 32842 4936 39630
rect 5000 39630 5226 39658
rect 4896 32836 4948 32842
rect 4896 32778 4948 32784
rect 5000 32042 5028 39630
rect 5170 39520 5226 39630
rect 5814 39658 5870 40000
rect 6366 39658 6422 40000
rect 7010 39658 7066 40000
rect 7654 39658 7710 40000
rect 5814 39630 6040 39658
rect 5814 39520 5870 39630
rect 5356 36780 5408 36786
rect 5356 36722 5408 36728
rect 5264 34944 5316 34950
rect 5264 34886 5316 34892
rect 5276 34542 5304 34886
rect 5264 34536 5316 34542
rect 5264 34478 5316 34484
rect 5276 33454 5304 34478
rect 5368 34202 5396 36722
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5356 34196 5408 34202
rect 5356 34138 5408 34144
rect 5080 33448 5132 33454
rect 5080 33390 5132 33396
rect 5264 33448 5316 33454
rect 5264 33390 5316 33396
rect 5092 32910 5120 33390
rect 5368 33386 5396 34138
rect 5356 33380 5408 33386
rect 5408 33340 5488 33368
rect 5356 33322 5408 33328
rect 5172 32972 5224 32978
rect 5172 32914 5224 32920
rect 5080 32904 5132 32910
rect 5080 32846 5132 32852
rect 5184 32502 5212 32914
rect 5172 32496 5224 32502
rect 5172 32438 5224 32444
rect 5000 32014 5304 32042
rect 4896 31136 4948 31142
rect 4896 31078 4948 31084
rect 4908 30870 4936 31078
rect 4896 30864 4948 30870
rect 4896 30806 4948 30812
rect 4908 30394 4936 30806
rect 4896 30388 4948 30394
rect 4896 30330 4948 30336
rect 5080 30116 5132 30122
rect 5080 30058 5132 30064
rect 5092 29850 5120 30058
rect 5080 29844 5132 29850
rect 5080 29786 5132 29792
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 4620 29174 4672 29180
rect 4802 29200 4858 29209
rect 4344 28960 4396 28966
rect 4344 28902 4396 28908
rect 4528 28960 4580 28966
rect 4528 28902 4580 28908
rect 4172 26982 4292 27010
rect 4068 26512 4120 26518
rect 4068 26454 4120 26460
rect 3976 24744 4028 24750
rect 3976 24686 4028 24692
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3988 23474 4016 24142
rect 4172 24070 4200 26982
rect 4436 25152 4488 25158
rect 4436 25094 4488 25100
rect 4448 24954 4476 25094
rect 4436 24948 4488 24954
rect 4436 24890 4488 24896
rect 4344 24676 4396 24682
rect 4344 24618 4396 24624
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 3344 23446 3464 23474
rect 3896 23446 4016 23474
rect 3148 23248 3200 23254
rect 3148 23190 3200 23196
rect 3344 22098 3372 23446
rect 3516 23112 3568 23118
rect 3516 23054 3568 23060
rect 3424 22500 3476 22506
rect 3424 22442 3476 22448
rect 3436 22234 3464 22442
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3344 21350 3372 22034
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3068 18550 3280 18578
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3068 17338 3096 17614
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3068 15910 3096 16594
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15434 3096 15846
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 3160 15094 3188 16390
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3252 11801 3280 18550
rect 3238 11792 3294 11801
rect 3238 11727 3294 11736
rect 112 8832 164 8838
rect 112 8774 164 8780
rect 124 6769 152 8774
rect 110 6760 166 6769
rect 110 6695 166 6704
rect 3344 6254 3372 21286
rect 3424 21140 3476 21146
rect 3424 21082 3476 21088
rect 3436 13734 3464 21082
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3436 12345 3464 13670
rect 3422 12336 3478 12345
rect 3422 12271 3478 12280
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 664 3120 716 3126
rect 664 3062 716 3068
rect 386 82 442 480
rect 676 82 704 3062
rect 3436 2514 3464 11727
rect 3528 10130 3556 23054
rect 3896 22964 3924 23446
rect 3976 23248 4028 23254
rect 4080 23236 4108 23598
rect 4264 23322 4292 24210
rect 4356 24206 4384 24618
rect 4344 24200 4396 24206
rect 4344 24142 4396 24148
rect 4448 24138 4476 24890
rect 4436 24132 4488 24138
rect 4436 24074 4488 24080
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4252 23316 4304 23322
rect 4252 23258 4304 23264
rect 4028 23208 4108 23236
rect 3976 23190 4028 23196
rect 3896 22936 4016 22964
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3884 22500 3936 22506
rect 3988 22488 4016 22936
rect 4080 22658 4108 23208
rect 4160 22704 4212 22710
rect 4080 22652 4160 22658
rect 4080 22646 4212 22652
rect 4080 22630 4200 22646
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 3936 22460 4016 22488
rect 3884 22442 3936 22448
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 4172 21554 4200 22510
rect 4264 22506 4292 23258
rect 4252 22500 4304 22506
rect 4252 22442 4304 22448
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4252 21072 4304 21078
rect 4252 21014 4304 21020
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18970 4200 19246
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 4080 18358 4108 18702
rect 4068 18352 4120 18358
rect 3974 18320 4030 18329
rect 4068 18294 4120 18300
rect 3974 18255 4030 18264
rect 3988 18222 4016 18255
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 4080 17134 4108 18022
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3988 16046 4016 16934
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 4080 12918 4108 13398
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 4080 10810 4108 11086
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 4080 3194 4108 3538
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3528 2582 3556 2790
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 386 54 704 82
rect 1214 82 1270 480
rect 1596 82 1624 2450
rect 3974 2408 4030 2417
rect 4264 2378 4292 21014
rect 4356 18442 4384 24006
rect 4540 23474 4568 28902
rect 4632 28762 4660 29174
rect 5000 29170 5028 29446
rect 5080 29232 5132 29238
rect 5080 29174 5132 29180
rect 4802 29135 4858 29144
rect 4988 29164 5040 29170
rect 4988 29106 5040 29112
rect 4804 29028 4856 29034
rect 4804 28970 4856 28976
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 4724 28694 4752 28902
rect 4712 28688 4764 28694
rect 4712 28630 4764 28636
rect 4816 28626 4844 28970
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 4816 28218 4844 28562
rect 4804 28212 4856 28218
rect 4804 28154 4856 28160
rect 5092 28014 5120 29174
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 5080 28008 5132 28014
rect 5080 27950 5132 27956
rect 5000 27674 5028 27950
rect 5092 27878 5120 27950
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 5092 27334 5120 27814
rect 5080 27328 5132 27334
rect 5080 27270 5132 27276
rect 4712 26988 4764 26994
rect 4712 26930 4764 26936
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4632 23866 4660 24074
rect 4724 23866 4752 26930
rect 4988 26920 5040 26926
rect 4988 26862 5040 26868
rect 4896 26444 4948 26450
rect 4896 26386 4948 26392
rect 4908 26042 4936 26386
rect 5000 26246 5028 26862
rect 5092 26858 5120 27270
rect 5080 26852 5132 26858
rect 5080 26794 5132 26800
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 5092 26058 5120 26794
rect 4896 26036 4948 26042
rect 4896 25978 4948 25984
rect 5000 26030 5120 26058
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4724 23594 4752 23802
rect 4816 23662 4844 24754
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 4712 23588 4764 23594
rect 4712 23530 4764 23536
rect 4540 23446 4660 23474
rect 4528 23180 4580 23186
rect 4528 23122 4580 23128
rect 4540 22778 4568 23122
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4436 22704 4488 22710
rect 4540 22681 4568 22714
rect 4436 22646 4488 22652
rect 4526 22672 4582 22681
rect 4448 21622 4476 22646
rect 4526 22607 4582 22616
rect 4436 21616 4488 21622
rect 4436 21558 4488 21564
rect 4448 21078 4476 21558
rect 4436 21072 4488 21078
rect 4436 21014 4488 21020
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4448 20602 4476 20878
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4448 20312 4476 20538
rect 4528 20324 4580 20330
rect 4448 20284 4528 20312
rect 4528 20266 4580 20272
rect 4632 18612 4660 23446
rect 4724 19514 4752 23530
rect 4896 23520 4948 23526
rect 4802 23488 4858 23497
rect 5000 23497 5028 26030
rect 5080 25696 5132 25702
rect 5080 25638 5132 25644
rect 5092 24614 5120 25638
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 5184 24682 5212 25094
rect 5172 24676 5224 24682
rect 5172 24618 5224 24624
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4896 23462 4948 23468
rect 4986 23488 5042 23497
rect 4802 23423 4858 23432
rect 4816 22778 4844 23423
rect 4804 22772 4856 22778
rect 4804 22714 4856 22720
rect 4816 22506 4844 22714
rect 4908 22642 4936 23462
rect 4986 23423 5042 23432
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4908 22234 4936 22578
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 5000 22098 5028 23258
rect 5092 23186 5120 23598
rect 5184 23526 5212 24618
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5184 23118 5212 23462
rect 5172 23112 5224 23118
rect 5172 23054 5224 23060
rect 4988 22092 5040 22098
rect 4988 22034 5040 22040
rect 4896 21888 4948 21894
rect 4896 21830 4948 21836
rect 4908 21418 4936 21830
rect 5000 21690 5028 22034
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4896 21412 4948 21418
rect 4896 21354 4948 21360
rect 4908 21010 4936 21354
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4908 20602 4936 20946
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 5000 20534 5028 21490
rect 4988 20528 5040 20534
rect 5276 20505 5304 32014
rect 5356 31204 5408 31210
rect 5356 31146 5408 31152
rect 5368 30734 5396 31146
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 5368 30258 5396 30670
rect 5356 30252 5408 30258
rect 5356 30194 5408 30200
rect 5356 29844 5408 29850
rect 5356 29786 5408 29792
rect 5368 29578 5396 29786
rect 5356 29572 5408 29578
rect 5356 29514 5408 29520
rect 5368 29170 5396 29514
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 5460 27062 5488 33340
rect 5552 28082 5580 34546
rect 5816 33992 5868 33998
rect 5816 33934 5868 33940
rect 5632 33856 5684 33862
rect 5632 33798 5684 33804
rect 5644 33368 5672 33798
rect 5828 33522 5856 33934
rect 5816 33516 5868 33522
rect 5816 33458 5868 33464
rect 5724 33380 5776 33386
rect 5644 33340 5724 33368
rect 5644 33114 5672 33340
rect 5724 33322 5776 33328
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 5632 33108 5684 33114
rect 5632 33050 5684 33056
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5644 32366 5672 32846
rect 5828 32774 5856 33254
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 5816 32768 5868 32774
rect 5816 32710 5868 32716
rect 5828 32434 5856 32710
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 5632 32360 5684 32366
rect 5684 32320 5764 32348
rect 5632 32302 5684 32308
rect 5632 31884 5684 31890
rect 5632 31826 5684 31832
rect 5644 31142 5672 31826
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5632 28960 5684 28966
rect 5632 28902 5684 28908
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5552 26246 5580 27474
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5368 25498 5396 26182
rect 5552 25838 5580 26182
rect 5540 25832 5592 25838
rect 5540 25774 5592 25780
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 5552 25362 5580 25774
rect 5644 25770 5672 28902
rect 5736 26790 5764 32320
rect 5828 31890 5856 32370
rect 5920 32298 5948 32846
rect 6012 32450 6040 39630
rect 6366 39630 6868 39658
rect 6366 39520 6422 39630
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6644 36304 6696 36310
rect 6644 36246 6696 36252
rect 6656 35494 6684 36246
rect 6644 35488 6696 35494
rect 6644 35430 6696 35436
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6184 35148 6236 35154
rect 6184 35090 6236 35096
rect 6196 34746 6224 35090
rect 6184 34740 6236 34746
rect 6184 34682 6236 34688
rect 6196 34513 6224 34682
rect 6182 34504 6238 34513
rect 6182 34439 6238 34448
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6656 34202 6684 35430
rect 6736 34468 6788 34474
rect 6736 34410 6788 34416
rect 6184 34196 6236 34202
rect 6184 34138 6236 34144
rect 6644 34196 6696 34202
rect 6644 34138 6696 34144
rect 6196 33658 6224 34138
rect 6748 33658 6776 34410
rect 6184 33652 6236 33658
rect 6184 33594 6236 33600
rect 6736 33652 6788 33658
rect 6736 33594 6788 33600
rect 6196 33046 6224 33594
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6184 33040 6236 33046
rect 6184 32982 6236 32988
rect 6012 32422 6132 32450
rect 6000 32360 6052 32366
rect 6000 32302 6052 32308
rect 5908 32292 5960 32298
rect 5908 32234 5960 32240
rect 5920 32026 5948 32234
rect 5908 32020 5960 32026
rect 5908 31962 5960 31968
rect 6012 31958 6040 32302
rect 6000 31952 6052 31958
rect 6000 31894 6052 31900
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5828 31210 5856 31826
rect 5908 31272 5960 31278
rect 5908 31214 5960 31220
rect 5816 31204 5868 31210
rect 5816 31146 5868 31152
rect 5920 30598 5948 31214
rect 6104 30920 6132 32422
rect 6196 32230 6224 32982
rect 6184 32224 6236 32230
rect 6184 32166 6236 32172
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6564 31482 6592 31758
rect 6736 31748 6788 31754
rect 6736 31690 6788 31696
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6748 31142 6776 31690
rect 6736 31136 6788 31142
rect 6736 31078 6788 31084
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6012 30892 6132 30920
rect 5908 30592 5960 30598
rect 5908 30534 5960 30540
rect 5920 30122 5948 30534
rect 5908 30116 5960 30122
rect 5908 30058 5960 30064
rect 5920 27130 5948 30058
rect 6012 27538 6040 30892
rect 6092 30796 6144 30802
rect 6092 30738 6144 30744
rect 6460 30796 6512 30802
rect 6460 30738 6512 30744
rect 6104 29510 6132 30738
rect 6184 30592 6236 30598
rect 6184 30534 6236 30540
rect 6092 29504 6144 29510
rect 6092 29446 6144 29452
rect 6104 28150 6132 29446
rect 6092 28144 6144 28150
rect 6092 28086 6144 28092
rect 6196 27606 6224 30534
rect 6472 30122 6500 30738
rect 6460 30116 6512 30122
rect 6460 30058 6512 30064
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6552 29776 6604 29782
rect 6552 29718 6604 29724
rect 6564 29238 6592 29718
rect 6644 29640 6696 29646
rect 6644 29582 6696 29588
rect 6552 29232 6604 29238
rect 6552 29174 6604 29180
rect 6656 28966 6684 29582
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6656 28762 6684 28902
rect 6644 28756 6696 28762
rect 6644 28698 6696 28704
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6276 28552 6328 28558
rect 6276 28494 6328 28500
rect 6288 28218 6316 28494
rect 6276 28212 6328 28218
rect 6276 28154 6328 28160
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6184 27600 6236 27606
rect 6184 27542 6236 27548
rect 6000 27532 6052 27538
rect 6000 27474 6052 27480
rect 5908 27124 5960 27130
rect 5908 27066 5960 27072
rect 6012 26994 6040 27474
rect 6184 27464 6236 27470
rect 6184 27406 6236 27412
rect 6196 27130 6224 27406
rect 6656 27334 6684 28562
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6656 27130 6684 27270
rect 6184 27124 6236 27130
rect 6184 27066 6236 27072
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6000 26988 6052 26994
rect 6000 26930 6052 26936
rect 6092 26852 6144 26858
rect 6092 26794 6144 26800
rect 5724 26784 5776 26790
rect 5724 26726 5776 26732
rect 6104 25906 6132 26794
rect 6092 25900 6144 25906
rect 6092 25842 6144 25848
rect 5632 25764 5684 25770
rect 5632 25706 5684 25712
rect 5540 25356 5592 25362
rect 5540 25298 5592 25304
rect 5356 24744 5408 24750
rect 5356 24686 5408 24692
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 5368 24342 5396 24686
rect 5356 24336 5408 24342
rect 5356 24278 5408 24284
rect 5460 23322 5488 24686
rect 5540 23588 5592 23594
rect 5540 23530 5592 23536
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5552 23186 5580 23530
rect 5644 23474 5672 25706
rect 6000 25492 6052 25498
rect 6000 25434 6052 25440
rect 5908 25356 5960 25362
rect 6012 25344 6040 25434
rect 5960 25316 6040 25344
rect 5908 25298 5960 25304
rect 5908 24676 5960 24682
rect 5908 24618 5960 24624
rect 5724 24268 5776 24274
rect 5724 24210 5776 24216
rect 5736 23730 5764 24210
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5828 23662 5856 24074
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5644 23446 5856 23474
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5460 22710 5488 23122
rect 5552 22778 5580 23122
rect 5632 23044 5684 23050
rect 5632 22986 5684 22992
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 5356 22500 5408 22506
rect 5356 22442 5408 22448
rect 5368 22234 5396 22442
rect 5644 22234 5672 22986
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5368 21690 5396 22170
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5736 20602 5764 23258
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 4988 20470 5040 20476
rect 5262 20496 5318 20505
rect 5000 19990 5028 20470
rect 5262 20431 5318 20440
rect 5276 20210 5304 20431
rect 5736 20398 5764 20538
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5092 20182 5304 20210
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4908 19242 4936 19858
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 5000 18834 5028 19790
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 5092 18714 5120 20182
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 19446 5304 19654
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5184 18834 5212 19246
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 4804 18692 4856 18698
rect 5092 18686 5212 18714
rect 4804 18634 4856 18640
rect 4632 18584 4752 18612
rect 4356 18414 4660 18442
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4436 17604 4488 17610
rect 4436 17546 4488 17552
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4356 13326 4384 14214
rect 4448 13938 4476 17546
rect 4540 17202 4568 18022
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4356 12986 4384 13262
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4356 9042 4384 10610
rect 4448 9994 4476 13738
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4540 9722 4568 10066
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8634 4384 8978
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4540 7546 4568 7890
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4632 6866 4660 18414
rect 4724 12889 4752 18584
rect 4816 18358 4844 18634
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4816 17542 4844 18090
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5092 17746 5120 18022
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4816 16454 4844 17478
rect 5092 17338 5120 17682
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16794 4936 16934
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4908 16046 4936 16730
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4908 15706 4936 15982
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 4896 15088 4948 15094
rect 4896 15030 4948 15036
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4710 12880 4766 12889
rect 4710 12815 4766 12824
rect 4712 12776 4764 12782
rect 4710 12744 4712 12753
rect 4764 12744 4766 12753
rect 4710 12679 4766 12688
rect 4724 12646 4752 12679
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4816 11336 4844 14962
rect 4908 14482 4936 15030
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4908 13814 4936 14418
rect 5184 13814 5212 18686
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5276 16998 5304 17818
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 15706 5304 16934
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5276 14958 5304 15506
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5264 14816 5316 14822
rect 5368 14804 5396 20198
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5460 18630 5488 19110
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5644 17134 5672 19110
rect 5828 18970 5856 23446
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5828 18290 5856 18906
rect 5920 18290 5948 24618
rect 6012 24070 6040 25316
rect 6092 25356 6144 25362
rect 6092 25298 6144 25304
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 6012 23118 6040 24006
rect 6104 23186 6132 25298
rect 6196 25294 6224 27066
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6460 26444 6512 26450
rect 6460 26386 6512 26392
rect 6472 26042 6500 26386
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6184 25288 6236 25294
rect 6184 25230 6236 25236
rect 6196 24138 6224 25230
rect 6748 25158 6776 31078
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6748 24750 6776 25094
rect 6736 24744 6788 24750
rect 6736 24686 6788 24692
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6184 24132 6236 24138
rect 6184 24074 6236 24080
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 23866 6684 24074
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6656 23322 6684 23802
rect 6644 23316 6696 23322
rect 6644 23258 6696 23264
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6104 22166 6132 23122
rect 6736 22500 6788 22506
rect 6736 22442 6788 22448
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6656 22166 6684 22374
rect 6748 22234 6776 22442
rect 6736 22228 6788 22234
rect 6840 22216 6868 39630
rect 6920 39636 6972 39642
rect 6920 39578 6972 39584
rect 7010 39630 7236 39658
rect 6932 30802 6960 39578
rect 7010 39520 7066 39630
rect 7208 36718 7236 39630
rect 7300 39630 7710 39658
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 7196 36576 7248 36582
rect 7196 36518 7248 36524
rect 7208 36174 7236 36518
rect 7196 36168 7248 36174
rect 7196 36110 7248 36116
rect 7208 35834 7236 36110
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 7012 35556 7064 35562
rect 7012 35498 7064 35504
rect 7196 35556 7248 35562
rect 7196 35498 7248 35504
rect 7024 35222 7052 35498
rect 7012 35216 7064 35222
rect 7012 35158 7064 35164
rect 7024 34746 7052 35158
rect 7208 34950 7236 35498
rect 7196 34944 7248 34950
rect 7196 34886 7248 34892
rect 7012 34740 7064 34746
rect 7012 34682 7064 34688
rect 7024 34202 7052 34682
rect 7208 34678 7236 34886
rect 7196 34672 7248 34678
rect 7196 34614 7248 34620
rect 7012 34196 7064 34202
rect 7012 34138 7064 34144
rect 7012 33380 7064 33386
rect 7012 33322 7064 33328
rect 7024 32774 7052 33322
rect 7012 32768 7064 32774
rect 7012 32710 7064 32716
rect 7024 31958 7052 32710
rect 7104 32224 7156 32230
rect 7104 32166 7156 32172
rect 7012 31952 7064 31958
rect 7012 31894 7064 31900
rect 7024 31482 7052 31894
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 6932 29102 6960 30602
rect 7116 30598 7144 32166
rect 7300 31328 7328 39630
rect 7654 39520 7710 39630
rect 8298 39658 8354 40000
rect 8298 39630 8708 39658
rect 8298 39520 8354 39630
rect 8392 39296 8444 39302
rect 8392 39238 8444 39244
rect 7656 36712 7708 36718
rect 7656 36654 7708 36660
rect 7380 34536 7432 34542
rect 7380 34478 7432 34484
rect 7392 34202 7420 34478
rect 7380 34196 7432 34202
rect 7380 34138 7432 34144
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7392 32366 7420 32710
rect 7564 32496 7616 32502
rect 7562 32464 7564 32473
rect 7616 32464 7618 32473
rect 7562 32399 7618 32408
rect 7380 32360 7432 32366
rect 7380 32302 7432 32308
rect 7300 31300 7420 31328
rect 7288 31204 7340 31210
rect 7288 31146 7340 31152
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 7012 30184 7064 30190
rect 7012 30126 7064 30132
rect 6920 29096 6972 29102
rect 6920 29038 6972 29044
rect 7024 28694 7052 30126
rect 7116 30122 7144 30534
rect 7104 30116 7156 30122
rect 7104 30058 7156 30064
rect 7116 29782 7144 30058
rect 7104 29776 7156 29782
rect 7104 29718 7156 29724
rect 7300 29102 7328 31146
rect 7288 29096 7340 29102
rect 7288 29038 7340 29044
rect 7012 28688 7064 28694
rect 7012 28630 7064 28636
rect 7300 28626 7328 29038
rect 7288 28620 7340 28626
rect 7288 28562 7340 28568
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 7012 27940 7064 27946
rect 7012 27882 7064 27888
rect 7024 27674 7052 27882
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 6932 23798 6960 26386
rect 7104 26376 7156 26382
rect 7104 26318 7156 26324
rect 7116 25498 7144 26318
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 7116 24886 7144 25434
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7024 24274 7052 24754
rect 7116 24342 7144 24822
rect 7104 24336 7156 24342
rect 7104 24278 7156 24284
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 6920 23792 6972 23798
rect 6918 23760 6920 23769
rect 6972 23760 6974 23769
rect 7024 23730 7052 24210
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 6918 23695 6974 23704
rect 7012 23724 7064 23730
rect 6932 23254 6960 23695
rect 7012 23666 7064 23672
rect 6920 23248 6972 23254
rect 6920 23190 6972 23196
rect 7024 22234 7052 23666
rect 7012 22228 7064 22234
rect 6840 22188 6960 22216
rect 6736 22170 6788 22176
rect 6092 22160 6144 22166
rect 6012 22120 6092 22148
rect 6012 19786 6040 22120
rect 6092 22102 6144 22108
rect 6644 22160 6696 22166
rect 6644 22102 6696 22108
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6840 21622 6868 22034
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6196 20262 6224 20946
rect 6564 20602 6592 20946
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6092 19712 6144 19718
rect 6092 19654 6144 19660
rect 6104 19378 6132 19654
rect 6288 19446 6316 19858
rect 6276 19440 6328 19446
rect 6276 19382 6328 19388
rect 6092 19372 6144 19378
rect 6288 19334 6316 19382
rect 6092 19314 6144 19320
rect 6104 18970 6132 19314
rect 6196 19306 6316 19334
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6196 18766 6224 19306
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 5998 18592 6054 18601
rect 5998 18527 6054 18536
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5828 18086 5856 18226
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5460 16114 5488 16526
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5552 16046 5580 16390
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5552 14958 5580 15982
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5368 14776 5580 14804
rect 5264 14758 5316 14764
rect 5276 14618 5304 14758
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5276 13938 5304 14554
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 4908 13802 5120 13814
rect 4896 13796 5120 13802
rect 4948 13786 5120 13796
rect 5184 13786 5488 13814
rect 4896 13738 4948 13744
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 12170 4936 13262
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11626 5028 12038
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 4816 11308 4936 11336
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4816 10810 4844 11154
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9178 4752 9862
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 8634 4844 10746
rect 4908 8974 4936 11308
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4908 8566 4936 8910
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4632 6458 4660 6802
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4632 4214 4660 4245
rect 4620 4208 4672 4214
rect 4618 4176 4620 4185
rect 4672 4176 4674 4185
rect 4618 4111 4674 4120
rect 4632 4078 4660 4111
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4618 3088 4674 3097
rect 4528 3052 4580 3058
rect 4618 3023 4674 3032
rect 4528 2994 4580 3000
rect 4540 2650 4568 2994
rect 4632 2922 4660 3023
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 3974 2343 4030 2352
rect 4252 2372 4304 2378
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 2318 2000 2374 2009
rect 2318 1935 2374 1944
rect 1214 54 1624 82
rect 2042 82 2098 480
rect 2332 82 2360 1935
rect 2042 54 2360 82
rect 2870 128 2926 480
rect 2870 76 2872 128
rect 2924 76 2926 128
rect 386 0 442 54
rect 1214 0 1270 54
rect 2042 0 2098 54
rect 2870 0 2926 76
rect 3698 82 3754 480
rect 3988 82 4016 2343
rect 4252 2314 4304 2320
rect 3698 54 4016 82
rect 4526 82 4582 480
rect 4816 82 4844 6394
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5000 3194 5028 3538
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5092 134 5120 13786
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5184 12918 5212 13262
rect 5276 13190 5304 13670
rect 5368 13462 5396 13670
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 5184 12442 5212 12854
rect 5368 12714 5396 13398
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5276 12442 5304 12650
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5460 12102 5488 13786
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5552 11898 5580 14776
rect 5644 13802 5672 15846
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5276 10266 5304 10474
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5184 7342 5212 8842
rect 5276 8430 5304 9114
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 7954 5304 8366
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5276 7546 5304 7890
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5276 7342 5304 7482
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5184 6866 5212 7278
rect 5276 6934 5304 7278
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5276 5846 5304 6870
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5184 4078 5212 4762
rect 5276 4282 5304 5782
rect 5368 4826 5396 10202
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5552 9042 5580 11834
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5552 8634 5580 8978
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5552 7410 5580 7822
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5644 5778 5672 13738
rect 5736 11354 5764 17478
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5920 16454 5948 16934
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5828 15502 5856 15914
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 14618 5856 15438
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5920 11898 5948 16390
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5736 10538 5764 11290
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5828 7834 5856 11630
rect 5920 11218 5948 11834
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5920 9382 5948 10134
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5736 7806 5856 7834
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5644 5370 5672 5714
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5276 4078 5304 4218
rect 5736 4154 5764 7806
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 7002 5856 7686
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 7002 5948 7210
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5908 4684 5960 4690
rect 6012 4672 6040 18527
rect 6196 17882 6224 18702
rect 6288 18358 6316 18770
rect 6276 18352 6328 18358
rect 6276 18294 6328 18300
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6748 16658 6776 21490
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6840 19310 6868 19722
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6840 18902 6868 19246
rect 6932 19242 6960 22188
rect 7012 22170 7064 22176
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6932 18834 6960 19178
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6932 17814 6960 18770
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7024 17882 7052 18158
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6748 16182 6776 16594
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 6104 13530 6132 15302
rect 6196 14890 6224 15642
rect 6748 15570 6776 16118
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6748 14618 6776 15506
rect 6840 15026 6868 15642
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 14074 6224 14350
rect 6656 14074 6684 14486
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6196 13530 6224 14010
rect 6656 13802 6684 14010
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6104 12986 6132 13466
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6104 12374 6132 12922
rect 6380 12714 6408 13194
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6092 12368 6144 12374
rect 6144 12328 6224 12356
rect 6092 12310 6144 12316
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6104 11558 6132 12174
rect 6196 11898 6224 12328
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6288 11665 6316 11698
rect 6274 11656 6330 11665
rect 6274 11591 6330 11600
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6104 11354 6132 11494
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6656 11218 6684 13194
rect 6748 12238 6776 14350
rect 6932 14056 6960 17002
rect 6840 14028 6960 14056
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6748 11354 6776 12174
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 10470 6684 11154
rect 6748 10538 6776 11290
rect 6840 11218 6868 14028
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6932 13530 6960 13874
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6656 9722 6684 10406
rect 6840 10266 6868 11154
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7024 10130 7052 10474
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6104 9042 6132 9386
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6656 9110 6684 9318
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6748 7274 6776 7958
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6656 6934 6684 7142
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 6118 6132 6734
rect 6748 6662 6776 7210
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6196 6118 6224 6190
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6104 5914 6132 6054
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6196 5148 6224 6054
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 5370 6592 5714
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6840 5302 6868 9930
rect 6932 9382 6960 9998
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9178 6960 9318
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7024 9042 7052 9454
rect 7116 9178 7144 23802
rect 7208 21554 7236 27950
rect 7288 26988 7340 26994
rect 7288 26930 7340 26936
rect 7300 25362 7328 26930
rect 7392 26450 7420 31300
rect 7472 30048 7524 30054
rect 7472 29990 7524 29996
rect 7484 28150 7512 29990
rect 7472 28144 7524 28150
rect 7472 28086 7524 28092
rect 7484 27878 7512 28086
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 7380 26444 7432 26450
rect 7380 26386 7432 26392
rect 7576 26314 7604 32399
rect 7668 28994 7696 36654
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 7748 36100 7800 36106
rect 7748 36042 7800 36048
rect 7760 35766 7788 36042
rect 7748 35760 7800 35766
rect 7748 35702 7800 35708
rect 7760 32892 7788 35702
rect 7840 35624 7892 35630
rect 7840 35566 7892 35572
rect 7852 34610 7880 35566
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 7840 34604 7892 34610
rect 7840 34546 7892 34552
rect 7840 34128 7892 34134
rect 7840 34070 7892 34076
rect 7852 33658 7880 34070
rect 7944 33998 7972 35022
rect 7932 33992 7984 33998
rect 7932 33934 7984 33940
rect 7840 33652 7892 33658
rect 7840 33594 7892 33600
rect 7944 33522 7972 33934
rect 8312 33658 8340 36518
rect 8300 33652 8352 33658
rect 8300 33594 8352 33600
rect 7932 33516 7984 33522
rect 7932 33458 7984 33464
rect 7944 33134 7972 33458
rect 7944 33106 8156 33134
rect 8024 33040 8076 33046
rect 8024 32982 8076 32988
rect 7932 32904 7984 32910
rect 7760 32864 7932 32892
rect 7932 32846 7984 32852
rect 7944 31958 7972 32846
rect 8036 32570 8064 32982
rect 8024 32564 8076 32570
rect 8024 32506 8076 32512
rect 8128 32026 8156 33106
rect 8208 32904 8260 32910
rect 8208 32846 8260 32852
rect 8116 32020 8168 32026
rect 8116 31962 8168 31968
rect 7932 31952 7984 31958
rect 7932 31894 7984 31900
rect 8128 31414 8156 31962
rect 8116 31408 8168 31414
rect 8116 31350 8168 31356
rect 8220 31346 8248 32846
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 7748 31204 7800 31210
rect 7748 31146 7800 31152
rect 7760 30598 7788 31146
rect 7840 30864 7892 30870
rect 7840 30806 7892 30812
rect 7748 30592 7800 30598
rect 7748 30534 7800 30540
rect 7760 30394 7788 30534
rect 7748 30388 7800 30394
rect 7748 30330 7800 30336
rect 7852 29850 7880 30806
rect 8220 30734 8248 31282
rect 8300 30932 8352 30938
rect 8300 30874 8352 30880
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 8208 30728 8260 30734
rect 8208 30670 8260 30676
rect 8036 30394 8064 30670
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 8036 29850 8064 30330
rect 8312 30138 8340 30874
rect 8220 30110 8340 30138
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 7668 28966 7788 28994
rect 7564 26308 7616 26314
rect 7564 26250 7616 26256
rect 7288 25356 7340 25362
rect 7288 25298 7340 25304
rect 7300 24750 7328 25298
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 7300 23526 7328 24346
rect 7380 24132 7432 24138
rect 7380 24074 7432 24080
rect 7392 23798 7420 24074
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7288 23520 7340 23526
rect 7288 23462 7340 23468
rect 7484 23322 7512 23666
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 8090 7052 8978
rect 7208 8974 7236 17818
rect 7300 16794 7328 22714
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 7392 21146 7420 21422
rect 7484 21418 7512 21898
rect 7576 21434 7604 23598
rect 7472 21412 7524 21418
rect 7576 21406 7696 21434
rect 7472 21354 7524 21360
rect 7484 21146 7512 21354
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7484 21010 7512 21082
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 18834 7420 20334
rect 7576 19990 7604 21286
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7392 18358 7420 18566
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7484 18222 7512 18566
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7392 17338 7420 18090
rect 7576 17746 7604 18770
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7392 17134 7420 17274
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7392 16658 7420 17070
rect 7576 16998 7604 17682
rect 7668 17678 7696 21406
rect 7760 20058 7788 28966
rect 8024 28960 8076 28966
rect 8024 28902 8076 28908
rect 8036 27674 8064 28902
rect 8116 28620 8168 28626
rect 8116 28562 8168 28568
rect 8128 28082 8156 28562
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 8024 27668 8076 27674
rect 8024 27610 8076 27616
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 7944 27062 7972 27474
rect 7932 27056 7984 27062
rect 7932 26998 7984 27004
rect 7840 26784 7892 26790
rect 7840 26726 7892 26732
rect 7852 23186 7880 26726
rect 7944 23474 7972 26998
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 8036 25158 8064 26386
rect 8024 25152 8076 25158
rect 8024 25094 8076 25100
rect 8024 24404 8076 24410
rect 8024 24346 8076 24352
rect 8036 24313 8064 24346
rect 8022 24304 8078 24313
rect 8022 24239 8078 24248
rect 8220 23866 8248 30110
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8312 29238 8340 29990
rect 8300 29232 8352 29238
rect 8300 29174 8352 29180
rect 8312 29034 8340 29174
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8312 28218 8340 28970
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 8312 27878 8340 28154
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8404 26518 8432 39238
rect 8576 37120 8628 37126
rect 8576 37062 8628 37068
rect 8588 36718 8616 37062
rect 8576 36712 8628 36718
rect 8576 36654 8628 36660
rect 8588 36038 8616 36654
rect 8576 36032 8628 36038
rect 8576 35974 8628 35980
rect 8576 35148 8628 35154
rect 8576 35090 8628 35096
rect 8588 34746 8616 35090
rect 8576 34740 8628 34746
rect 8576 34682 8628 34688
rect 8588 33134 8616 34682
rect 8680 34490 8708 39630
rect 8850 39636 8906 40000
rect 9494 39658 9550 40000
rect 10138 39658 10194 40000
rect 10690 39658 10746 40000
rect 11334 39658 11390 40000
rect 11978 39658 12034 40000
rect 8850 39584 8852 39636
rect 8904 39584 8906 39636
rect 8850 39520 8906 39584
rect 9232 39630 9550 39658
rect 9232 39302 9260 39630
rect 9494 39520 9550 39630
rect 10060 39630 10194 39658
rect 9220 39296 9272 39302
rect 9220 39238 9272 39244
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 9680 36236 9732 36242
rect 9680 36178 9732 36184
rect 9496 36032 9548 36038
rect 9496 35974 9548 35980
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9508 35630 9536 35974
rect 9496 35624 9548 35630
rect 9496 35566 9548 35572
rect 8760 35488 8812 35494
rect 8760 35430 8812 35436
rect 8772 34610 8800 35430
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8760 34604 8812 34610
rect 8760 34546 8812 34552
rect 8680 34462 8800 34490
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8680 33386 8708 33798
rect 8668 33380 8720 33386
rect 8668 33322 8720 33328
rect 8588 33106 8708 33134
rect 8576 32836 8628 32842
rect 8576 32778 8628 32784
rect 8588 31890 8616 32778
rect 8576 31884 8628 31890
rect 8576 31826 8628 31832
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8496 28626 8524 31622
rect 8588 31142 8616 31826
rect 8576 31136 8628 31142
rect 8576 31078 8628 31084
rect 8576 30728 8628 30734
rect 8576 30670 8628 30676
rect 8588 30190 8616 30670
rect 8576 30184 8628 30190
rect 8576 30126 8628 30132
rect 8484 28620 8536 28626
rect 8484 28562 8536 28568
rect 8496 28218 8524 28562
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8484 28008 8536 28014
rect 8484 27950 8536 27956
rect 8496 27674 8524 27950
rect 8576 27940 8628 27946
rect 8576 27882 8628 27888
rect 8484 27668 8536 27674
rect 8484 27610 8536 27616
rect 8588 27538 8616 27882
rect 8576 27532 8628 27538
rect 8576 27474 8628 27480
rect 8588 26790 8616 27474
rect 8576 26784 8628 26790
rect 8576 26726 8628 26732
rect 8392 26512 8444 26518
rect 8392 26454 8444 26460
rect 8588 26450 8616 26726
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 7944 23446 8064 23474
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7852 22778 7880 23122
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7944 21146 7972 21422
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 8036 21010 8064 23446
rect 8312 23254 8340 23734
rect 8300 23248 8352 23254
rect 8300 23190 8352 23196
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8128 21146 8156 21966
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8024 21004 8076 21010
rect 8024 20946 8076 20952
rect 8036 20602 8064 20946
rect 8024 20596 8076 20602
rect 8076 20556 8156 20584
rect 8024 20538 8076 20544
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7760 19310 7788 19858
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7392 16250 7420 16594
rect 7668 16454 7696 17070
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7760 16266 7788 18294
rect 7852 17270 7880 19790
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 7944 17202 7972 17682
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7576 16238 7788 16266
rect 7392 15978 7420 16186
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7392 12714 7420 13874
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7300 11898 7328 12310
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7116 8498 7144 8910
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 6934 7052 7346
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6186 7052 6598
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6932 5914 6960 6122
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 5846 7052 6122
rect 7116 5846 7144 7822
rect 7208 6458 7236 8230
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 5960 4644 6040 4672
rect 5908 4626 5960 4632
rect 6012 4282 6040 4644
rect 6104 5120 6224 5148
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 4185 6132 5120
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6196 4486 6224 4694
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6090 4176 6146 4185
rect 5736 4126 5948 4154
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3670 5304 4014
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5368 2922 5396 3402
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5736 3058 5764 3334
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 4526 54 4844 82
rect 5080 128 5132 134
rect 5080 70 5132 76
rect 5354 96 5410 480
rect 3698 0 3754 54
rect 4526 0 4582 54
rect 5920 82 5948 4126
rect 6090 4111 6146 4120
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 6012 3534 6040 3946
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6012 2650 6040 3470
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6104 2310 6132 3878
rect 6196 3466 6224 4422
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6288 4146 6316 4218
rect 6840 4154 6868 5238
rect 7116 4554 7144 5782
rect 7300 5302 7328 11562
rect 7392 10062 7420 12650
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7484 9654 7512 10134
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7576 9586 7604 16238
rect 7840 16176 7892 16182
rect 7840 16118 7892 16124
rect 7852 16046 7880 16118
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15706 7880 15982
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7668 13814 7696 14826
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14550 7788 14758
rect 7852 14618 7880 15370
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7944 14482 7972 17138
rect 8036 16658 8064 17614
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8036 15706 8064 16594
rect 8128 16182 8156 20556
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8312 19446 8340 19994
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 8312 18970 8340 19382
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8220 15570 8248 18702
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8312 16726 8340 17274
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8312 16250 8340 16662
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8036 15162 8064 15506
rect 8220 15162 8248 15506
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8036 14958 8064 15098
rect 8312 15026 8340 15914
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7944 14074 7972 14418
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7668 13786 7972 13814
rect 7944 13462 7972 13786
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 7944 13190 7972 13398
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12986 7972 13126
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7944 12714 7972 12922
rect 8036 12850 8064 14554
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8128 13870 8156 14010
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8128 13258 8156 13806
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12442 7972 12650
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7944 11898 7972 12378
rect 8220 12374 8248 12582
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7760 11286 7788 11630
rect 7944 11626 7972 11834
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7944 11286 7972 11562
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7944 10810 7972 11222
rect 8128 11082 8156 12174
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7668 10062 7696 10610
rect 7944 10266 7972 10746
rect 8220 10266 8248 11086
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7944 9110 7972 10202
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7944 8566 7972 9046
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7932 8560 7984 8566
rect 7932 8502 7984 8508
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7576 7206 7604 7822
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6186 7604 7142
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6644 4140 6696 4146
rect 6840 4126 7052 4154
rect 7576 4146 7604 6122
rect 8036 5846 8064 8774
rect 8220 8430 8248 8910
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 7546 8156 7958
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8128 7002 8156 7210
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8128 6390 8156 6938
rect 8116 6384 8168 6390
rect 8168 6344 8248 6372
rect 8116 6326 8168 6332
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 8036 5370 8064 5782
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4554 7788 4966
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 6644 4082 6696 4088
rect 6288 4049 6316 4082
rect 6274 4040 6330 4049
rect 6274 3975 6330 3984
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6288 3194 6316 3606
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6564 3126 6592 3334
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6656 3058 6684 4082
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3126 6776 3878
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6748 2650 6776 3062
rect 6840 3058 6868 3538
rect 6932 3398 6960 3946
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 6274 82 6330 480
rect 5920 54 6330 82
rect 7024 82 7052 4126
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7760 2582 7788 4490
rect 7852 3738 7880 4762
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8128 4214 8156 4626
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8220 4146 8248 6344
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8220 3670 8248 4082
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8036 2650 8064 3538
rect 8220 3194 8248 3606
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8220 2922 8248 3130
rect 8312 3126 8340 14282
rect 8404 9602 8432 26250
rect 8588 25702 8616 26386
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 8496 24614 8524 24822
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8496 24342 8524 24550
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 8588 24138 8616 25638
rect 8576 24132 8628 24138
rect 8576 24074 8628 24080
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 8496 22438 8524 23122
rect 8484 22432 8536 22438
rect 8484 22374 8536 22380
rect 8496 21418 8524 22374
rect 8680 21536 8708 33106
rect 8772 30938 8800 34462
rect 9416 34202 9444 35022
rect 9404 34196 9456 34202
rect 9404 34138 9456 34144
rect 8852 33924 8904 33930
rect 8852 33866 8904 33872
rect 8864 33114 8892 33866
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8852 33108 8904 33114
rect 8852 33050 8904 33056
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 9310 31784 9366 31793
rect 9310 31719 9366 31728
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9036 31272 9088 31278
rect 9036 31214 9088 31220
rect 8760 30932 8812 30938
rect 8760 30874 8812 30880
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 8772 28694 8800 30670
rect 9048 30666 9076 31214
rect 9036 30660 9088 30666
rect 9036 30602 9088 30608
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 9324 30394 9352 31719
rect 9508 31686 9536 35566
rect 9692 35494 9720 36178
rect 9680 35488 9732 35494
rect 9680 35430 9732 35436
rect 9864 35216 9916 35222
rect 9864 35158 9916 35164
rect 9876 34406 9904 35158
rect 10060 34474 10088 39630
rect 10138 39520 10194 39630
rect 10428 39630 10746 39658
rect 10232 36644 10284 36650
rect 10232 36586 10284 36592
rect 10244 35630 10272 36586
rect 10428 36378 10456 39630
rect 10690 39520 10746 39630
rect 11072 39630 11390 39658
rect 10416 36372 10468 36378
rect 10416 36314 10468 36320
rect 11072 35834 11100 39630
rect 11334 39520 11390 39630
rect 11532 39630 12034 39658
rect 11532 36922 11560 39630
rect 11978 39520 12034 39630
rect 12530 39658 12586 40000
rect 13174 39658 13230 40000
rect 13818 39658 13874 40000
rect 14370 39658 14426 40000
rect 15014 39658 15070 40000
rect 12530 39630 12664 39658
rect 12530 39520 12586 39630
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 12070 37496 12126 37505
rect 12070 37431 12126 37440
rect 11520 36916 11572 36922
rect 11520 36858 11572 36864
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 11060 35828 11112 35834
rect 11060 35770 11112 35776
rect 10232 35624 10284 35630
rect 10232 35566 10284 35572
rect 10692 35488 10744 35494
rect 10744 35448 10824 35476
rect 10692 35430 10744 35436
rect 10508 35080 10560 35086
rect 10508 35022 10560 35028
rect 10048 34468 10100 34474
rect 10048 34410 10100 34416
rect 9864 34400 9916 34406
rect 9864 34342 9916 34348
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9680 32904 9732 32910
rect 9680 32846 9732 32852
rect 9692 32502 9720 32846
rect 9784 32774 9812 33934
rect 9772 32768 9824 32774
rect 9772 32710 9824 32716
rect 9876 32570 9904 34342
rect 10060 34202 10088 34410
rect 10324 34400 10376 34406
rect 10324 34342 10376 34348
rect 10048 34196 10100 34202
rect 10048 34138 10100 34144
rect 10060 33658 10088 34138
rect 10048 33652 10100 33658
rect 10048 33594 10100 33600
rect 10060 33386 10088 33594
rect 10336 33590 10364 34342
rect 10520 34134 10548 35022
rect 10508 34128 10560 34134
rect 10508 34070 10560 34076
rect 10692 33856 10744 33862
rect 10692 33798 10744 33804
rect 10324 33584 10376 33590
rect 10324 33526 10376 33532
rect 10704 33454 10732 33798
rect 10692 33448 10744 33454
rect 10692 33390 10744 33396
rect 10048 33380 10100 33386
rect 10048 33322 10100 33328
rect 10060 33257 10088 33322
rect 10324 33040 10376 33046
rect 10324 32982 10376 32988
rect 9956 32768 10008 32774
rect 9956 32710 10008 32716
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 9864 32564 9916 32570
rect 9864 32506 9916 32512
rect 9680 32496 9732 32502
rect 9680 32438 9732 32444
rect 9692 32026 9720 32438
rect 9876 32230 9904 32506
rect 9864 32224 9916 32230
rect 9864 32166 9916 32172
rect 9968 32026 9996 32710
rect 10060 32434 10088 32710
rect 10336 32570 10364 32982
rect 10324 32564 10376 32570
rect 10324 32506 10376 32512
rect 10048 32428 10100 32434
rect 10048 32370 10100 32376
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 9956 32020 10008 32026
rect 9956 31962 10008 31968
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9496 31680 9548 31686
rect 9496 31622 9548 31628
rect 9508 31278 9536 31622
rect 9692 31482 9720 31826
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9496 31272 9548 31278
rect 9496 31214 9548 31220
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9496 31136 9548 31142
rect 9496 31078 9548 31084
rect 9312 30388 9364 30394
rect 9312 30330 9364 30336
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8760 28688 8812 28694
rect 8760 28630 8812 28636
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8852 27940 8904 27946
rect 8852 27882 8904 27888
rect 8760 26376 8812 26382
rect 8760 26318 8812 26324
rect 8772 25498 8800 26318
rect 8864 26042 8892 27882
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8852 26036 8904 26042
rect 8852 25978 8904 25984
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8772 24818 8800 25434
rect 8864 24886 8892 25978
rect 9324 25838 9352 26182
rect 9312 25832 9364 25838
rect 9312 25774 9364 25780
rect 9404 25764 9456 25770
rect 9404 25706 9456 25712
rect 9416 25498 9444 25706
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8944 24676 8996 24682
rect 8944 24618 8996 24624
rect 9404 24676 9456 24682
rect 9404 24618 9456 24624
rect 8956 24206 8984 24618
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8772 23594 8800 24006
rect 8760 23588 8812 23594
rect 8760 23530 8812 23536
rect 8864 23322 8892 24142
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9324 23798 9352 24210
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9312 23520 9364 23526
rect 9312 23462 9364 23468
rect 8852 23316 8904 23322
rect 8852 23258 8904 23264
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8772 22642 8800 23054
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8772 22234 8800 22578
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8680 21508 8800 21536
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8496 21010 8524 21354
rect 8680 21146 8708 21354
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8496 19922 8524 20946
rect 8680 20466 8708 21082
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8680 19310 8708 19654
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8496 18222 8524 18770
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13326 8708 13670
rect 8772 13530 8800 21508
rect 9324 20942 9352 23462
rect 9416 22778 9444 24618
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9416 22438 9444 22714
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 22166 9444 22374
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9416 21690 9444 22102
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9416 21418 9444 21626
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 9416 20602 9444 21354
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9416 20330 9444 20538
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 8864 18426 8892 19110
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 9324 18154 9352 19110
rect 9416 18426 9444 20266
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9312 18148 9364 18154
rect 9312 18090 9364 18096
rect 9416 17882 9444 18158
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9140 16794 9168 17070
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8864 15162 8892 16186
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9140 15706 9168 16050
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8864 14890 8892 15098
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8956 14618 8984 14962
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8482 12880 8538 12889
rect 8482 12815 8538 12824
rect 8496 10146 8524 12815
rect 8588 12374 8616 13126
rect 8680 12986 8708 13262
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10266 8616 10610
rect 8680 10538 8708 11834
rect 8864 11558 8892 14418
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 9140 11354 9168 11698
rect 9324 11626 9352 16390
rect 9508 16114 9536 31078
rect 9784 30258 9812 31146
rect 10048 30932 10100 30938
rect 10048 30874 10100 30880
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 9784 29850 9812 30194
rect 10060 30122 10088 30874
rect 10048 30116 10100 30122
rect 10048 30058 10100 30064
rect 9772 29844 9824 29850
rect 9772 29786 9824 29792
rect 10048 29776 10100 29782
rect 10048 29718 10100 29724
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 9784 28762 9812 29582
rect 10060 28966 10088 29718
rect 10796 29594 10824 35448
rect 10876 34944 10928 34950
rect 10876 34886 10928 34892
rect 10888 34678 10916 34886
rect 10876 34672 10928 34678
rect 10876 34614 10928 34620
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 10980 33046 11008 34546
rect 10968 33040 11020 33046
rect 10968 32982 11020 32988
rect 10980 32434 11008 32982
rect 10968 32428 11020 32434
rect 10968 32370 11020 32376
rect 10876 31680 10928 31686
rect 10876 31622 10928 31628
rect 10888 31210 10916 31622
rect 10980 31346 11008 32370
rect 11164 31890 11192 36518
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11244 36236 11296 36242
rect 11244 36178 11296 36184
rect 11256 35494 11284 36178
rect 12084 35834 12112 37431
rect 12636 36378 12664 39630
rect 12820 39630 13230 39658
rect 12624 36372 12676 36378
rect 12624 36314 12676 36320
rect 12072 35828 12124 35834
rect 12072 35770 12124 35776
rect 12440 35624 12492 35630
rect 12440 35566 12492 35572
rect 11244 35488 11296 35494
rect 11244 35430 11296 35436
rect 12072 35488 12124 35494
rect 12072 35430 12124 35436
rect 11152 31884 11204 31890
rect 11152 31826 11204 31832
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10876 31204 10928 31210
rect 10876 31146 10928 31152
rect 10888 30938 10916 31146
rect 10980 30938 11008 31282
rect 10876 30932 10928 30938
rect 10876 30874 10928 30880
rect 10968 30932 11020 30938
rect 10968 30874 11020 30880
rect 10876 30728 10928 30734
rect 10876 30670 10928 30676
rect 10888 30394 10916 30670
rect 10876 30388 10928 30394
rect 10876 30330 10928 30336
rect 10796 29566 11008 29594
rect 10416 29504 10468 29510
rect 10416 29446 10468 29452
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10428 29034 10456 29446
rect 10416 29028 10468 29034
rect 10416 28970 10468 28976
rect 10048 28960 10100 28966
rect 10048 28902 10100 28908
rect 9772 28756 9824 28762
rect 9772 28698 9824 28704
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 9692 24274 9720 28018
rect 10060 28014 10088 28902
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10048 28008 10100 28014
rect 10048 27950 10100 27956
rect 10232 28008 10284 28014
rect 10232 27950 10284 27956
rect 9864 27940 9916 27946
rect 9864 27882 9916 27888
rect 9876 27849 9904 27882
rect 9862 27840 9918 27849
rect 9862 27775 9918 27784
rect 10060 27606 10088 27950
rect 10048 27600 10100 27606
rect 10048 27542 10100 27548
rect 10060 27130 10088 27542
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 10152 26586 10180 27406
rect 10244 27402 10272 27950
rect 10232 27396 10284 27402
rect 10232 27338 10284 27344
rect 10244 26994 10272 27338
rect 10336 27334 10364 28494
rect 10428 27674 10456 28970
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10704 28218 10732 28902
rect 10692 28212 10744 28218
rect 10692 28154 10744 28160
rect 10600 27940 10652 27946
rect 10600 27882 10652 27888
rect 10508 27872 10560 27878
rect 10612 27849 10640 27882
rect 10508 27814 10560 27820
rect 10598 27840 10654 27849
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 10324 26512 10376 26518
rect 10520 26500 10548 27814
rect 10598 27775 10654 27784
rect 10796 27470 10824 29446
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 10888 28626 10916 29106
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10888 27606 10916 28562
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 10888 26994 10916 27542
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10600 26852 10652 26858
rect 10600 26794 10652 26800
rect 10612 26586 10640 26794
rect 10980 26586 11008 29566
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 11164 28218 11192 28630
rect 11152 28212 11204 28218
rect 11152 28154 11204 28160
rect 11256 27062 11284 35430
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 11532 34474 11560 35090
rect 11520 34468 11572 34474
rect 11520 34410 11572 34416
rect 11980 34400 12032 34406
rect 11980 34342 12032 34348
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11520 34128 11572 34134
rect 11520 34070 11572 34076
rect 11704 34128 11756 34134
rect 11704 34070 11756 34076
rect 11428 33312 11480 33318
rect 11428 33254 11480 33260
rect 11440 33046 11468 33254
rect 11532 33114 11560 34070
rect 11716 33658 11744 34070
rect 11704 33652 11756 33658
rect 11704 33594 11756 33600
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11520 33108 11572 33114
rect 11520 33050 11572 33056
rect 11428 33040 11480 33046
rect 11428 32982 11480 32988
rect 11440 32570 11468 32982
rect 11992 32892 12020 34342
rect 12084 33930 12112 35430
rect 12164 34672 12216 34678
rect 12164 34614 12216 34620
rect 12072 33924 12124 33930
rect 12072 33866 12124 33872
rect 12084 33046 12112 33866
rect 12072 33040 12124 33046
rect 12072 32982 12124 32988
rect 12072 32904 12124 32910
rect 11992 32864 12072 32892
rect 12072 32846 12124 32852
rect 12084 32570 12112 32846
rect 12176 32570 12204 34614
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12268 34513 12296 34546
rect 12254 34504 12310 34513
rect 12254 34439 12310 34448
rect 12348 34468 12400 34474
rect 12348 34410 12400 34416
rect 12256 33040 12308 33046
rect 12256 32982 12308 32988
rect 11428 32564 11480 32570
rect 11428 32506 11480 32512
rect 12072 32564 12124 32570
rect 12072 32506 12124 32512
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 12162 32464 12218 32473
rect 12162 32399 12218 32408
rect 12176 32366 12204 32399
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11336 31884 11388 31890
rect 11336 31826 11388 31832
rect 11348 31142 11376 31826
rect 12268 31346 12296 32982
rect 12256 31340 12308 31346
rect 12256 31282 12308 31288
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11244 26852 11296 26858
rect 11244 26794 11296 26800
rect 10600 26580 10652 26586
rect 10600 26522 10652 26528
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 10376 26472 10548 26500
rect 10324 26454 10376 26460
rect 10612 26042 10640 26522
rect 10692 26512 10744 26518
rect 10692 26454 10744 26460
rect 10704 26042 10732 26454
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9784 24410 9812 25774
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10060 25498 10088 25638
rect 10704 25498 10732 25978
rect 10796 25702 10824 26318
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10796 25498 10824 25638
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10888 24818 10916 25298
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9692 23526 9720 24210
rect 9968 23866 9996 24346
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10152 24138 10180 24210
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 10152 23866 10180 24074
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10704 23594 10732 24006
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 10704 23254 10732 23530
rect 10980 23474 11008 26522
rect 11256 26518 11284 26794
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 11256 25838 11284 26454
rect 11244 25832 11296 25838
rect 11244 25774 11296 25780
rect 11256 25430 11284 25774
rect 11244 25424 11296 25430
rect 11244 25366 11296 25372
rect 11256 24818 11284 25366
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 11348 23474 11376 31078
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 12268 30870 12296 31282
rect 11612 30864 11664 30870
rect 11612 30806 11664 30812
rect 12256 30864 12308 30870
rect 12256 30806 12308 30812
rect 11520 30728 11572 30734
rect 11520 30670 11572 30676
rect 11532 30394 11560 30670
rect 11520 30388 11572 30394
rect 11520 30330 11572 30336
rect 11532 29850 11560 30330
rect 11624 30326 11652 30806
rect 11612 30320 11664 30326
rect 11612 30262 11664 30268
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11520 29844 11572 29850
rect 11520 29786 11572 29792
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 12268 29306 12296 29650
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12256 29096 12308 29102
rect 12256 29038 12308 29044
rect 11520 29028 11572 29034
rect 11520 28970 11572 28976
rect 11532 27588 11560 28970
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11704 27600 11756 27606
rect 11532 27560 11704 27588
rect 11704 27542 11756 27548
rect 11612 27464 11664 27470
rect 11532 27424 11612 27452
rect 11532 26586 11560 27424
rect 11612 27406 11664 27412
rect 11716 27130 11744 27542
rect 11978 27432 12034 27441
rect 11978 27367 12034 27376
rect 11796 27328 11848 27334
rect 11796 27270 11848 27276
rect 11808 27130 11836 27270
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11992 26042 12020 27367
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12084 26897 12112 26930
rect 12070 26888 12126 26897
rect 12070 26823 12126 26832
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12084 26042 12112 26386
rect 11980 26036 12032 26042
rect 11980 25978 12032 25984
rect 12072 26036 12124 26042
rect 12072 25978 12124 25984
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 12268 24954 12296 29038
rect 12360 28218 12388 34410
rect 12452 29782 12480 35566
rect 12820 35290 12848 39630
rect 13174 39520 13230 39630
rect 13740 39630 13874 39658
rect 13740 35834 13768 39630
rect 13818 39520 13874 39630
rect 14108 39630 14426 39658
rect 13728 35828 13780 35834
rect 13728 35770 13780 35776
rect 14108 35290 14136 39630
rect 14370 39520 14426 39630
rect 14752 39630 15070 39658
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 12808 35284 12860 35290
rect 12808 35226 12860 35232
rect 14096 35284 14148 35290
rect 14096 35226 14148 35232
rect 12716 35148 12768 35154
rect 12716 35090 12768 35096
rect 12728 34610 12756 35090
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 13912 34536 13964 34542
rect 13912 34478 13964 34484
rect 13544 34060 13596 34066
rect 13544 34002 13596 34008
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 12544 33522 12572 33798
rect 12532 33516 12584 33522
rect 12532 33458 12584 33464
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 12544 32026 12572 33458
rect 12820 33046 12848 33458
rect 13556 33318 13584 34002
rect 13544 33312 13596 33318
rect 13544 33254 13596 33260
rect 12808 33040 12860 33046
rect 12808 32982 12860 32988
rect 13556 32978 13584 33254
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13556 32230 13584 32914
rect 13544 32224 13596 32230
rect 13544 32166 13596 32172
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 12440 29776 12492 29782
rect 12440 29718 12492 29724
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 12452 28694 12480 29582
rect 13360 28960 13412 28966
rect 13360 28902 13412 28908
rect 13372 28762 13400 28902
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 12440 28688 12492 28694
rect 12440 28630 12492 28636
rect 12348 28212 12400 28218
rect 12348 28154 12400 28160
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12360 24562 12388 28154
rect 12452 27538 12480 28630
rect 13268 28620 13320 28626
rect 13268 28562 13320 28568
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12636 27674 12664 28358
rect 13280 28218 13308 28562
rect 13268 28212 13320 28218
rect 13268 28154 13320 28160
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 12452 25362 12480 27474
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12360 24534 12572 24562
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23730 11468 24006
rect 11532 23866 11560 24210
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 12072 23792 12124 23798
rect 12072 23734 12124 23740
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 10796 23446 11008 23474
rect 11256 23446 11376 23474
rect 10416 23248 10468 23254
rect 10336 23208 10416 23236
rect 10336 22438 10364 23208
rect 10416 23190 10468 23196
rect 10692 23248 10744 23254
rect 10692 23190 10744 23196
rect 10796 23032 10824 23446
rect 10520 23004 10824 23032
rect 11152 23044 11204 23050
rect 10520 22681 10548 23004
rect 11152 22986 11204 22992
rect 10968 22704 11020 22710
rect 10506 22672 10562 22681
rect 10968 22646 11020 22652
rect 10506 22607 10562 22616
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10336 22098 10364 22374
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9692 21486 9720 21966
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9600 20806 9628 21422
rect 9692 21078 9720 21422
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 10060 21146 10088 21354
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9692 20398 9720 20878
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9692 20058 9720 20334
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9876 19174 9904 19246
rect 10060 19174 10088 20742
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10244 19310 10272 19858
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10428 18970 10456 19926
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9600 17746 9628 18702
rect 9692 18290 9720 18770
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9784 18086 9812 18362
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17882 9812 18022
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9600 16794 9628 17682
rect 9784 17338 9812 17818
rect 9876 17814 9904 18294
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 17882 10364 18022
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9692 15570 9720 16526
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 14618 9720 15506
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9784 12850 9812 16050
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9968 15706 9996 15914
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9968 15162 9996 15642
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 14550 9904 14758
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 10520 14346 10548 22607
rect 10980 22506 11008 22646
rect 11164 22642 11192 22986
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 10968 22500 11020 22506
rect 10968 22442 11020 22448
rect 10980 22234 11008 22442
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10796 21078 10824 21830
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 11164 20942 11192 22578
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10980 20466 11008 20742
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10876 19984 10928 19990
rect 10980 19972 11008 20266
rect 11072 19990 11100 20742
rect 11164 20534 11192 20878
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 10928 19944 11008 19972
rect 10876 19926 10928 19932
rect 10980 19514 11008 19944
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11256 19334 11284 23446
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11348 22642 11376 23054
rect 11440 22710 11468 23666
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11428 22704 11480 22710
rect 11428 22646 11480 22652
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11428 22432 11480 22438
rect 11428 22374 11480 22380
rect 11348 21894 11376 22374
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11164 19306 11284 19334
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10704 18834 10732 19178
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10704 18426 10732 18770
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10796 16726 10824 17070
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10612 16250 10640 16526
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10600 15904 10652 15910
rect 10704 15892 10732 16662
rect 10652 15864 10732 15892
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10612 15162 10640 15302
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10612 14822 10640 15098
rect 10888 15094 10916 17070
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10980 15026 11008 15302
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 11072 14890 11100 16526
rect 11164 15094 11192 19306
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 15638 11284 16934
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10612 14074 10640 14758
rect 11072 14482 11100 14826
rect 11256 14618 11284 15574
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10612 13802 10640 14010
rect 10888 13938 10916 14282
rect 11164 14074 11192 14486
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 11348 13814 11376 21286
rect 11440 18329 11468 22374
rect 11532 20806 11560 23530
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 12084 23322 12112 23734
rect 12452 23594 12480 24142
rect 12440 23588 12492 23594
rect 12440 23530 12492 23536
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12072 23316 12124 23322
rect 12268 23304 12296 23462
rect 12452 23322 12480 23530
rect 12440 23316 12492 23322
rect 12268 23276 12388 23304
rect 12072 23258 12124 23264
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11980 23180 12032 23186
rect 11980 23122 12032 23128
rect 11900 22420 11928 23122
rect 11992 22778 12020 23122
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 12084 22438 12112 22918
rect 12360 22545 12388 23276
rect 12440 23258 12492 23264
rect 12544 23202 12572 24534
rect 12728 24313 12756 27814
rect 13082 27568 13138 27577
rect 13082 27503 13084 27512
rect 13136 27503 13138 27512
rect 13084 27474 13136 27480
rect 13096 27130 13124 27474
rect 13084 27124 13136 27130
rect 13084 27066 13136 27072
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12714 24304 12770 24313
rect 12714 24239 12770 24248
rect 12452 23174 12572 23202
rect 12728 23186 12756 24239
rect 12716 23180 12768 23186
rect 12346 22536 12402 22545
rect 12256 22500 12308 22506
rect 12346 22471 12402 22480
rect 12256 22442 12308 22448
rect 12072 22432 12124 22438
rect 11900 22392 12020 22420
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11992 22166 12020 22392
rect 12072 22374 12124 22380
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11624 21690 11652 22102
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11704 21072 11756 21078
rect 11704 21014 11756 21020
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11716 20602 11744 21014
rect 11992 20602 12020 21830
rect 12084 21554 12112 21898
rect 12176 21690 12204 21966
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12084 20874 12112 21490
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 12176 20058 12204 21626
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11426 18320 11482 18329
rect 11426 18255 11482 18264
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11440 16794 11468 17818
rect 11532 17814 11560 18702
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11532 17338 11560 17750
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17338 12204 17478
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11716 15162 11744 15574
rect 12084 15434 12112 17002
rect 12176 16998 12204 17274
rect 12268 17134 12296 22442
rect 12452 21350 12480 23174
rect 12716 23122 12768 23128
rect 12820 22778 12848 26998
rect 13096 23474 13124 27066
rect 12912 23446 13124 23474
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12820 22506 12848 22714
rect 12912 22574 12940 23446
rect 12900 22568 12952 22574
rect 12900 22510 12952 22516
rect 13174 22536 13230 22545
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12544 21418 12572 21898
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12624 21412 12676 21418
rect 12624 21354 12676 21360
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12544 20806 12572 21354
rect 12636 21146 12664 21354
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12912 21026 12940 22510
rect 13174 22471 13230 22480
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21622 13124 21966
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 12636 20998 12940 21026
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12346 20496 12402 20505
rect 12346 20431 12402 20440
rect 12360 20398 12388 20431
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12544 17066 12572 17478
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12176 16250 12204 16662
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11624 14074 11652 14350
rect 11992 14074 12020 14758
rect 12084 14346 12112 15370
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12636 13814 12664 20998
rect 13188 20942 13216 22471
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13464 21690 13492 22102
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13280 21010 13308 21490
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13280 20602 13308 20946
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 17610 12756 20334
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12820 17202 12848 17614
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16726 12848 17138
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 12820 16046 12848 16662
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12912 16182 12940 16526
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12728 14414 12756 15302
rect 13004 15094 13032 15506
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12728 14074 12756 14350
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 11256 13786 11376 13814
rect 12544 13786 12664 13814
rect 10244 13530 10272 13738
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9876 12918 9904 13398
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9692 12714 9720 12786
rect 9784 12753 9812 12786
rect 9770 12744 9826 12753
rect 9680 12708 9732 12714
rect 9770 12679 9826 12688
rect 10232 12708 10284 12714
rect 9680 12650 9732 12656
rect 10232 12650 10284 12656
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 12102 9536 12582
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10810 8800 10950
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8864 10674 8892 11290
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8496 10118 8708 10146
rect 8404 9574 8524 9602
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8404 9110 8432 9454
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8496 9042 8524 9574
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8404 4078 8432 5034
rect 8588 4690 8616 5102
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8588 4282 8616 4626
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8574 4176 8630 4185
rect 8574 4111 8630 4120
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8404 3738 8432 4014
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8312 2854 8340 3062
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 8588 2514 8616 4111
rect 8680 3097 8708 10118
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8864 8498 8892 9454
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7342 8800 7822
rect 8864 7410 8892 8298
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 8760 7336 8812 7342
rect 8812 7284 8892 7290
rect 8760 7278 8892 7284
rect 8772 7262 8892 7278
rect 8772 7213 8800 7262
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6186 8800 6598
rect 8864 6304 8892 7262
rect 9232 7002 9260 7346
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8944 6316 8996 6322
rect 8864 6276 8944 6304
rect 8944 6258 8996 6264
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 5914 8800 6122
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8956 5846 8984 6258
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 5370 9352 8434
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8864 4146 8892 5170
rect 9416 5166 9444 11494
rect 9508 9178 9536 12038
rect 9600 11830 9628 12310
rect 9692 11898 9720 12650
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9784 11354 9812 12174
rect 10244 12170 10272 12650
rect 10520 12170 10548 13194
rect 10888 12986 10916 13262
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9876 10810 9904 11222
rect 10244 11150 10272 12106
rect 10520 11762 10548 12106
rect 10888 11762 10916 12922
rect 11150 11792 11206 11801
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10876 11756 10928 11762
rect 11150 11727 11206 11736
rect 10876 11698 10928 11704
rect 11164 11694 11192 11727
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10428 11286 10456 11562
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10428 10674 10456 11222
rect 10796 10742 10824 11494
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10152 10198 10180 10474
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10266 10640 10406
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9586 9720 9998
rect 9784 9722 9812 10134
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9600 7954 9628 9386
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8634 9720 8978
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9600 7546 9628 7890
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 9324 3602 9352 4966
rect 9416 4826 9444 5102
rect 9692 4826 9720 8570
rect 9784 8022 9812 9658
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 8974 10456 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10244 8430 10272 8842
rect 10796 8634 10824 8978
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9784 7478 9812 7958
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9784 7274 9812 7414
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9784 6934 9812 7210
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9784 6458 9812 6870
rect 9876 6866 9904 8230
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 6934 10180 7142
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9876 5914 9904 6802
rect 10336 6322 10364 7822
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10428 6186 10456 6870
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10612 5846 10640 7686
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5370 10180 5646
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9416 3738 9444 4558
rect 9784 4214 9812 4694
rect 10152 4622 10180 5306
rect 10612 5234 10640 5782
rect 10980 5778 11008 6122
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 10152 4154 10180 4558
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10416 4208 10468 4214
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8666 3088 8722 3097
rect 9416 3058 9444 3674
rect 8666 3023 8722 3032
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9600 2650 9628 3878
rect 9784 3398 9812 4150
rect 10152 4126 10364 4154
rect 10416 4150 10468 4156
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9876 3194 9904 3606
rect 10336 3466 10364 4126
rect 10428 3534 10456 4150
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 3194 10180 3334
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10152 2854 10180 3130
rect 10428 3058 10456 3470
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10416 2916 10468 2922
rect 10520 2904 10548 3674
rect 10704 3602 10732 3878
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10796 3058 10824 4490
rect 11072 4214 11100 6054
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10468 2876 10548 2904
rect 10416 2858 10468 2864
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7102 82 7158 480
rect 7024 54 7158 82
rect 7576 82 7604 2314
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 7930 82 7986 480
rect 7576 54 7986 82
rect 8680 82 8708 2246
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8758 82 8814 480
rect 8680 54 8814 82
rect 5354 0 5410 40
rect 6274 0 6330 54
rect 7102 0 7158 54
rect 7930 0 7986 54
rect 8758 0 8814 54
rect 9586 82 9642 480
rect 9876 82 9904 2246
rect 9586 54 9904 82
rect 10336 82 10364 2586
rect 10888 2417 10916 4014
rect 11164 3398 11192 4966
rect 11256 4078 11284 13786
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11518 12880 11574 12889
rect 11518 12815 11574 12824
rect 11532 12782 11560 12815
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11992 12646 12020 13330
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11348 12374 11376 12582
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 12070 12472 12126 12481
rect 12070 12407 12126 12416
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11348 11898 11376 12310
rect 11992 11898 12020 12310
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 12084 11354 12112 12407
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10810 11468 11086
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11440 6458 11468 6938
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11532 6118 11560 6734
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11992 5778 12020 6734
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 5370 12020 5714
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11348 4690 11376 5102
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11348 4282 11376 4626
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11532 3738 11560 5034
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 12176 4154 12204 11630
rect 12348 7472 12400 7478
rect 12438 7440 12494 7449
rect 12400 7420 12438 7426
rect 12348 7414 12438 7420
rect 12360 7398 12438 7414
rect 12438 7375 12494 7384
rect 12544 5370 12572 13786
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 11218 12664 12582
rect 12912 12345 12940 14894
rect 12898 12336 12954 12345
rect 12898 12271 12954 12280
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10470 12664 11154
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12084 4126 12204 4154
rect 11704 4072 11756 4078
rect 11624 4049 11704 4060
rect 11610 4040 11704 4049
rect 11666 4032 11704 4040
rect 11704 4014 11756 4020
rect 11610 3975 11666 3984
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 2514 11192 3334
rect 11256 2582 11284 3402
rect 11440 3194 11468 3606
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11808 3194 11836 3470
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11520 3120 11572 3126
rect 11334 3088 11390 3097
rect 11520 3062 11572 3068
rect 11334 3023 11390 3032
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11348 2514 11376 3023
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 10874 2408 10930 2417
rect 10874 2343 10930 2352
rect 10414 82 10470 480
rect 10336 54 10470 82
rect 9586 0 9642 54
rect 10414 0 10470 54
rect 11334 82 11390 480
rect 11532 82 11560 3062
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 12084 2009 12112 4126
rect 12070 2000 12126 2009
rect 12070 1935 12126 1944
rect 11334 54 11560 82
rect 12162 82 12218 480
rect 12268 82 12296 4422
rect 12360 4282 12388 4626
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12636 2514 12664 10406
rect 12912 4154 12940 12271
rect 13004 11898 13032 15030
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13280 11937 13308 12242
rect 13266 11928 13322 11937
rect 12992 11892 13044 11898
rect 13266 11863 13322 11872
rect 12992 11834 13044 11840
rect 13004 11694 13032 11834
rect 13280 11830 13308 11863
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 12992 11688 13044 11694
rect 13372 11665 13400 14894
rect 13556 14822 13584 32166
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 13740 28665 13768 29038
rect 13726 28656 13782 28665
rect 13726 28591 13782 28600
rect 13924 20602 13952 34478
rect 14752 34202 14780 39630
rect 15014 39520 15070 39630
rect 15658 39658 15714 40000
rect 15658 39630 15792 39658
rect 15658 39520 15714 39630
rect 15764 34746 15792 39630
rect 15752 34740 15804 34746
rect 15752 34682 15804 34688
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13924 20398 13952 20538
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14738 17504 14794 17513
rect 14289 17436 14585 17456
rect 14738 17439 14794 17448
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14752 16250 14780 17439
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 12992 11630 13044 11636
rect 13358 11656 13414 11665
rect 13358 11591 13414 11600
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 12912 4126 13032 4154
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12162 54 12296 82
rect 12728 82 12756 3878
rect 13004 3194 13032 4126
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13096 3534 13124 3878
rect 13372 3602 13400 4966
rect 13464 4690 13492 12786
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13464 4282 13492 4626
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13372 3194 13400 3538
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13004 2990 13032 3130
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 13648 2553 13676 5510
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 13912 4548 13964 4554
rect 13912 4490 13964 4496
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13634 2544 13690 2553
rect 13634 2479 13690 2488
rect 13832 2417 13860 4014
rect 13818 2408 13874 2417
rect 13818 2343 13874 2352
rect 12990 82 13046 480
rect 12728 54 13046 82
rect 11334 0 11390 54
rect 12162 0 12218 54
rect 12990 0 13046 54
rect 13818 82 13874 480
rect 13924 82 13952 4490
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13818 54 13952 82
rect 14200 82 14228 4422
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14646 82 14702 480
rect 14200 54 14702 82
rect 13818 0 13874 54
rect 14646 0 14702 54
rect 15474 82 15530 480
rect 15580 82 15608 3334
rect 15474 54 15608 82
rect 15474 0 15530 54
<< via2 >>
rect 570 33088 626 33144
rect 1490 27512 1546 27568
rect 2870 22516 2872 22536
rect 2872 22516 2924 22536
rect 2924 22516 2926 22536
rect 2870 22480 2926 22516
rect 110 20032 166 20088
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3422 28600 3478 28656
rect 3238 23704 3294 23760
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3238 11736 3294 11792
rect 110 6704 166 6760
rect 3422 12280 3478 12336
rect 3422 11736 3478 11792
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3974 18264 4030 18320
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3974 2352 4030 2408
rect 4802 29144 4858 29200
rect 4526 22616 4582 22672
rect 4802 23432 4858 23488
rect 4986 23432 5042 23488
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6182 34448 6238 34504
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 5262 20440 5318 20496
rect 4710 12824 4766 12880
rect 4710 12724 4712 12744
rect 4712 12724 4764 12744
rect 4764 12724 4766 12744
rect 4710 12688 4766 12724
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 7562 32444 7564 32464
rect 7564 32444 7616 32464
rect 7616 32444 7618 32464
rect 7562 32408 7618 32444
rect 6918 23740 6920 23760
rect 6920 23740 6972 23760
rect 6972 23740 6974 23760
rect 6918 23704 6974 23740
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 5998 18536 6054 18592
rect 4618 4156 4620 4176
rect 4620 4156 4672 4176
rect 4672 4156 4674 4176
rect 4618 4120 4674 4156
rect 4618 3032 4674 3088
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 2318 1944 2374 2000
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6274 11600 6330 11656
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 8022 24248 8078 24304
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 5354 40 5410 96
rect 6090 4120 6146 4176
rect 6274 3984 6330 4040
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 9310 31728 9366 31784
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 12070 37440 12126 37496
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8482 12824 8538 12880
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 9862 27784 9918 27840
rect 10598 27784 10654 27840
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 12254 34448 12310 34504
rect 12162 32408 12218 32464
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11978 27376 12034 27432
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 12070 26832 12126 26888
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 10506 22616 10562 22672
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 13082 27532 13138 27568
rect 13082 27512 13084 27532
rect 13084 27512 13136 27532
rect 13136 27512 13138 27532
rect 12714 24248 12770 24304
rect 12346 22480 12402 22536
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11426 18264 11482 18320
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 13174 22480 13230 22536
rect 12346 20440 12402 20496
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 9770 12688 9826 12744
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8574 4120 8630 4176
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 11150 11736 11206 11792
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8666 3032 8722 3088
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11518 12824 11574 12880
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 12070 12416 12126 12472
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 12438 7384 12494 7440
rect 12898 12280 12954 12336
rect 11610 3984 11666 4040
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11334 3032 11390 3088
rect 10874 2352 10930 2408
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12070 1944 12126 2000
rect 13266 11872 13322 11928
rect 13726 28600 13782 28656
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14738 17448 14794 17504
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 13358 11600 13414 11656
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 13634 2488 13690 2544
rect 13818 2352 13874 2408
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 12065 37498 12131 37501
rect 15520 37498 16000 37528
rect 12065 37496 16000 37498
rect 12065 37440 12070 37496
rect 12126 37440 16000 37496
rect 12065 37438 16000 37440
rect 12065 37435 12131 37438
rect 15520 37408 16000 37438
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 6177 34506 6243 34509
rect 9438 34506 9444 34508
rect 6177 34504 9444 34506
rect 6177 34448 6182 34504
rect 6238 34448 9444 34504
rect 6177 34446 9444 34448
rect 6177 34443 6243 34446
rect 9438 34444 9444 34446
rect 9508 34506 9514 34508
rect 12249 34506 12315 34509
rect 9508 34504 12315 34506
rect 9508 34448 12254 34504
rect 12310 34448 12315 34504
rect 9508 34446 12315 34448
rect 9508 34444 9514 34446
rect 12249 34443 12315 34446
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 0 33328 480 33448
rect 62 33146 122 33328
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 565 33146 631 33149
rect 62 33144 631 33146
rect 62 33088 570 33144
rect 626 33088 631 33144
rect 62 33086 631 33088
rect 565 33083 631 33086
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 7557 32466 7623 32469
rect 12157 32466 12223 32469
rect 15520 32466 16000 32496
rect 7557 32464 12223 32466
rect 7557 32408 7562 32464
rect 7618 32408 12162 32464
rect 12218 32408 12223 32464
rect 7557 32406 12223 32408
rect 7557 32403 7623 32406
rect 12157 32403 12223 32406
rect 15518 32376 16000 32466
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 9305 31786 9371 31789
rect 15518 31786 15578 32376
rect 9305 31784 15578 31786
rect 9305 31728 9310 31784
rect 9366 31728 15578 31784
rect 9305 31726 15578 31728
rect 9305 31723 9371 31726
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 4797 29202 4863 29205
rect 6126 29202 6132 29204
rect 4797 29200 6132 29202
rect 4797 29144 4802 29200
rect 4858 29144 6132 29200
rect 4797 29142 6132 29144
rect 4797 29139 4863 29142
rect 6126 29140 6132 29142
rect 6196 29140 6202 29204
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 3417 28658 3483 28661
rect 13721 28658 13787 28661
rect 3417 28656 13787 28658
rect 3417 28600 3422 28656
rect 3478 28600 13726 28656
rect 13782 28600 13787 28656
rect 3417 28598 13787 28600
rect 3417 28595 3483 28598
rect 13721 28595 13787 28598
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 9857 27842 9923 27845
rect 10593 27842 10659 27845
rect 9857 27840 10659 27842
rect 9857 27784 9862 27840
rect 9918 27784 10598 27840
rect 10654 27784 10659 27840
rect 9857 27782 10659 27784
rect 9857 27779 9923 27782
rect 10593 27779 10659 27782
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 1485 27570 1551 27573
rect 13077 27570 13143 27573
rect 1485 27568 13143 27570
rect 1485 27512 1490 27568
rect 1546 27512 13082 27568
rect 13138 27512 13143 27568
rect 1485 27510 13143 27512
rect 1485 27507 1551 27510
rect 13077 27507 13143 27510
rect 11973 27434 12039 27437
rect 15520 27434 16000 27464
rect 11973 27432 16000 27434
rect 11973 27376 11978 27432
rect 12034 27376 16000 27432
rect 11973 27374 16000 27376
rect 11973 27371 12039 27374
rect 15520 27344 16000 27374
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 6126 26828 6132 26892
rect 6196 26890 6202 26892
rect 12065 26890 12131 26893
rect 6196 26888 12131 26890
rect 6196 26832 12070 26888
rect 12126 26832 12131 26888
rect 6196 26830 12131 26832
rect 6196 26828 6202 26830
rect 12065 26827 12131 26830
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 8017 24306 8083 24309
rect 12709 24306 12775 24309
rect 8017 24304 12775 24306
rect 8017 24248 8022 24304
rect 8078 24248 12714 24304
rect 12770 24248 12775 24304
rect 8017 24246 12775 24248
rect 8017 24243 8083 24246
rect 12709 24243 12775 24246
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 3233 23762 3299 23765
rect 6913 23762 6979 23765
rect 3233 23760 6979 23762
rect 3233 23704 3238 23760
rect 3294 23704 6918 23760
rect 6974 23704 6979 23760
rect 3233 23702 6979 23704
rect 3233 23699 3299 23702
rect 6913 23699 6979 23702
rect 4797 23490 4863 23493
rect 4981 23490 5047 23493
rect 4797 23488 5047 23490
rect 4797 23432 4802 23488
rect 4858 23432 4986 23488
rect 5042 23432 5047 23488
rect 4797 23430 5047 23432
rect 4797 23427 4863 23430
rect 4981 23427 5047 23430
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 4521 22674 4587 22677
rect 10501 22674 10567 22677
rect 4521 22672 10567 22674
rect 4521 22616 4526 22672
rect 4582 22616 10506 22672
rect 10562 22616 10567 22672
rect 4521 22614 10567 22616
rect 4521 22611 4587 22614
rect 10501 22611 10567 22614
rect 2865 22538 2931 22541
rect 12341 22538 12407 22541
rect 2865 22536 12407 22538
rect 2865 22480 2870 22536
rect 2926 22480 12346 22536
rect 12402 22480 12407 22536
rect 2865 22478 12407 22480
rect 2865 22475 2931 22478
rect 12341 22475 12407 22478
rect 13169 22538 13235 22541
rect 15520 22538 16000 22568
rect 13169 22536 16000 22538
rect 13169 22480 13174 22536
rect 13230 22480 16000 22536
rect 13169 22478 16000 22480
rect 13169 22475 13235 22478
rect 15520 22448 16000 22478
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 5257 20498 5323 20501
rect 12341 20498 12407 20501
rect 5257 20496 12407 20498
rect 5257 20440 5262 20496
rect 5318 20440 12346 20496
rect 12402 20440 12407 20496
rect 5257 20438 12407 20440
rect 5257 20435 5323 20438
rect 12341 20435 12407 20438
rect 6277 20160 6597 20161
rect 0 20088 480 20120
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 0 20032 110 20088
rect 166 20032 480 20088
rect 0 20000 480 20032
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 5993 18594 6059 18597
rect 6126 18594 6132 18596
rect 5993 18592 6132 18594
rect 5993 18536 5998 18592
rect 6054 18536 6132 18592
rect 5993 18534 6132 18536
rect 5993 18531 6059 18534
rect 6126 18532 6132 18534
rect 6196 18532 6202 18596
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 3969 18322 4035 18325
rect 11421 18322 11487 18325
rect 3969 18320 11487 18322
rect 3969 18264 3974 18320
rect 4030 18264 11426 18320
rect 11482 18264 11487 18320
rect 3969 18262 11487 18264
rect 3969 18259 4035 18262
rect 11421 18259 11487 18262
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 14733 17506 14799 17509
rect 15520 17506 16000 17536
rect 14733 17504 16000 17506
rect 14733 17448 14738 17504
rect 14794 17448 16000 17504
rect 14733 17446 16000 17448
rect 14733 17443 14799 17446
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 15520 17416 16000 17446
rect 14277 17375 14597 17376
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 4705 12882 4771 12885
rect 8477 12882 8543 12885
rect 11513 12882 11579 12885
rect 4705 12880 11579 12882
rect 4705 12824 4710 12880
rect 4766 12824 8482 12880
rect 8538 12824 11518 12880
rect 11574 12824 11579 12880
rect 4705 12822 11579 12824
rect 4705 12819 4771 12822
rect 8477 12819 8543 12822
rect 11513 12819 11579 12822
rect 4705 12746 4771 12749
rect 9765 12746 9831 12749
rect 4705 12744 9831 12746
rect 4705 12688 4710 12744
rect 4766 12688 9770 12744
rect 9826 12688 9831 12744
rect 4705 12686 9831 12688
rect 4705 12683 4771 12686
rect 9765 12683 9831 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 12065 12474 12131 12477
rect 15520 12474 16000 12504
rect 12065 12472 16000 12474
rect 12065 12416 12070 12472
rect 12126 12416 16000 12472
rect 12065 12414 16000 12416
rect 12065 12411 12131 12414
rect 15520 12384 16000 12414
rect 3417 12338 3483 12341
rect 12893 12338 12959 12341
rect 3417 12336 12959 12338
rect 3417 12280 3422 12336
rect 3478 12280 12898 12336
rect 12954 12280 12959 12336
rect 3417 12278 12959 12280
rect 3417 12275 3483 12278
rect 12893 12275 12959 12278
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 9438 11868 9444 11932
rect 9508 11930 9514 11932
rect 13261 11930 13327 11933
rect 9508 11928 13327 11930
rect 9508 11872 13266 11928
rect 13322 11872 13327 11928
rect 9508 11870 13327 11872
rect 9508 11868 9514 11870
rect 13261 11867 13327 11870
rect 3233 11794 3299 11797
rect 3417 11794 3483 11797
rect 11145 11794 11211 11797
rect 3233 11792 11211 11794
rect 3233 11736 3238 11792
rect 3294 11736 3422 11792
rect 3478 11736 11150 11792
rect 11206 11736 11211 11792
rect 3233 11734 11211 11736
rect 3233 11731 3299 11734
rect 3417 11731 3483 11734
rect 11145 11731 11211 11734
rect 6269 11658 6335 11661
rect 13353 11658 13419 11661
rect 6269 11656 13419 11658
rect 6269 11600 6274 11656
rect 6330 11600 13358 11656
rect 13414 11600 13419 11656
rect 6269 11598 13419 11600
rect 6269 11595 6335 11598
rect 13353 11595 13419 11598
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 12433 7442 12499 7445
rect 15520 7442 16000 7472
rect 12433 7440 16000 7442
rect 12433 7384 12438 7440
rect 12494 7384 16000 7440
rect 12433 7382 16000 7384
rect 12433 7379 12499 7382
rect 15520 7352 16000 7382
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 0 6760 480 6792
rect 0 6704 110 6760
rect 166 6704 480 6760
rect 0 6672 480 6704
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 4613 4178 4679 4181
rect 6085 4178 6151 4181
rect 8569 4178 8635 4181
rect 4613 4176 8635 4178
rect 4613 4120 4618 4176
rect 4674 4120 6090 4176
rect 6146 4120 8574 4176
rect 8630 4120 8635 4176
rect 4613 4118 8635 4120
rect 4613 4115 4679 4118
rect 6085 4115 6151 4118
rect 8569 4115 8635 4118
rect 6269 4042 6335 4045
rect 11605 4042 11671 4045
rect 6269 4040 11671 4042
rect 6269 3984 6274 4040
rect 6330 3984 11610 4040
rect 11666 3984 11671 4040
rect 6269 3982 11671 3984
rect 6269 3979 6335 3982
rect 11605 3979 11671 3982
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 4613 3090 4679 3093
rect 8661 3090 8727 3093
rect 11329 3090 11395 3093
rect 4613 3088 11395 3090
rect 4613 3032 4618 3088
rect 4674 3032 8666 3088
rect 8722 3032 11334 3088
rect 11390 3032 11395 3088
rect 4613 3030 11395 3032
rect 4613 3027 4679 3030
rect 8661 3027 8727 3030
rect 11329 3027 11395 3030
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 13629 2546 13695 2549
rect 15520 2546 16000 2576
rect 13629 2544 16000 2546
rect 13629 2488 13634 2544
rect 13690 2488 16000 2544
rect 13629 2486 16000 2488
rect 13629 2483 13695 2486
rect 15520 2456 16000 2486
rect 3969 2410 4035 2413
rect 10869 2410 10935 2413
rect 13813 2410 13879 2413
rect 3969 2408 13879 2410
rect 3969 2352 3974 2408
rect 4030 2352 10874 2408
rect 10930 2352 13818 2408
rect 13874 2352 13879 2408
rect 3969 2350 13879 2352
rect 3969 2347 4035 2350
rect 10869 2347 10935 2350
rect 13813 2347 13879 2350
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 2313 2002 2379 2005
rect 12065 2002 12131 2005
rect 2313 2000 12131 2002
rect 2313 1944 2318 2000
rect 2374 1944 12070 2000
rect 12126 1944 12131 2000
rect 2313 1942 12131 1944
rect 2313 1939 2379 1942
rect 12065 1939 12131 1942
rect 5349 98 5415 101
rect 9438 98 9444 100
rect 5349 96 9444 98
rect 5349 40 5354 96
rect 5410 40 9444 96
rect 5349 38 9444 40
rect 5349 35 5415 38
rect 9438 36 9444 38
rect 9508 36 9514 100
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 9444 34444 9508 34508
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6132 29140 6196 29204
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6132 26828 6196 26892
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 6132 18532 6196 18596
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 9444 11868 9508 11932
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
rect 9444 36 9508 100
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6131 29204 6197 29205
rect 6131 29140 6132 29204
rect 6196 29140 6197 29204
rect 6131 29139 6197 29140
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 6134 26893 6194 29139
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6131 26892 6197 26893
rect 6131 26828 6132 26892
rect 6196 26828 6197 26892
rect 6131 26827 6197 26828
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 6134 18597 6194 26827
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6131 18596 6197 18597
rect 6131 18532 6132 18596
rect 6196 18532 6197 18596
rect 6131 18531 6197 18532
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 9443 34508 9509 34509
rect 9443 34444 9444 34508
rect 9508 34444 9509 34508
rect 9443 34443 9509 34444
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 9446 11933 9506 34443
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 9443 11932 9509 11933
rect 9443 11868 9444 11932
rect 9508 11868 9509 11932
rect 9443 11867 9509 11868
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 9446 101 9506 11867
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
rect 9443 100 9509 101
rect 9443 36 9444 100
rect 9508 36 9509 100
rect 9443 35 9509 36
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_21 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_25 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_73
timestamp 1586364061
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_77
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _200_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_109
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _178_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_48
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_138 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_73
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_126
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_70
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_47
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _181_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 774 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_41
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_106
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_145
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_38
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_48
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_136
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_42
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_46
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_87
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_69
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_42
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_68
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_113
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_33
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_37
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_76
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_107
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_111
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_115
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_139
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_49
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_109
timestamp 1586364061
transform 1 0 11132 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_38
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_38
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_24_55
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_72
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 774 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_31
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_42
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_48
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_52
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_102
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_115
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_111
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_decap_12  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_140
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_144
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_38
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_58
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_62
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_66
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_buf_1  _081_
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_41
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_or3_4  _069_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_48
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_52
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_4  FILLER_30_96
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 406 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_118
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_26
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 130 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_or3_4  _098_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_or3_4  _080_
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__C
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_8  _067_
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_43
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 406 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_60
timestamp 1586364061
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_81
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_85
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_32_98
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 774 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_120
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_132
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_144
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 3312 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_8  _159_
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_44
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_57
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_67
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_71
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_104
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_108
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_113
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_121
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_130
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_126
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_137
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_132
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_141
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_145
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_144
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_30
timestamp 1586364061
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_66
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_70
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_83
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_103
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_35_140
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_18
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_38
timestamp 1586364061
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_36_53
timestamp 1586364061
transform 1 0 5980 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_1  _093_
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_58
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_65
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_69
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_104
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 2300 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_20
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_33
timestamp 1586364061
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_37
timestamp 1586364061
transform 1 0 4508 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 6072 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_52
timestamp 1586364061
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_56
timestamp 1586364061
transform 1 0 6256 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_60
timestamp 1586364061
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_77
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_81
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_97
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_102
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_137
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_141
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_145
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_or2_4  _171_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 -1 23392
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 4784 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_35
timestamp 1586364061
transform 1 0 4324 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_39
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 130 592
use scs8hd_nor3_4  _155_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 23392
box -38 -48 1234 592
use scs8hd_decap_3  FILLER_38_42
timestamp 1586364061
transform 1 0 4968 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_58
timestamp 1586364061
transform 1 0 6440 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_63
timestamp 1586364061
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_67
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_97
timestamp 1586364061
transform 1 0 10028 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_109
timestamp 1586364061
transform 1 0 11132 0 -1 23392
box -38 -48 774 592
use scs8hd_or2_4  _077_
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 682 592
use scs8hd_fill_2  FILLER_38_124
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _120_
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 866 592
use scs8hd_nor3_4  _156_
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 1234 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 4140 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__C
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_32
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_1  _076_
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 6164 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_42
timestamp 1586364061
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_53
timestamp 1586364061
transform 1 0 5980 0 -1 24480
box -38 -48 222 592
use scs8hd_or3_4  _119_
timestamp 1586364061
transform 1 0 6716 0 -1 24480
box -38 -48 866 592
use scs8hd_or4_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 6532 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_57
timestamp 1586364061
transform 1 0 6348 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_74
timestamp 1586364061
transform 1 0 7912 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_70
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 7728 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_81
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_78
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 314 592
use scs8hd_or4_4  _147_
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__D
timestamp 1586364061
transform 1 0 9108 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_91
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_95
timestamp 1586364061
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_85
timestamp 1586364061
transform 1 0 8924 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_89
timestamp 1586364061
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 11224 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_99
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_119
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_144
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_36
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_or4_4  _095_
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_or4_4  _137_
timestamp 1586364061
transform 1 0 6992 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_73
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_77
timestamp 1586364061
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_81
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_97
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_101
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 774 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__D
timestamp 1586364061
transform 1 0 4692 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 4324 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_37
timestamp 1586364061
transform 1 0 4508 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_41
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 222 592
use scs8hd_nor3_4  _157_
timestamp 1586364061
transform 1 0 5244 0 -1 25568
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 5060 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 7176 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_58
timestamp 1586364061
transform 1 0 6440 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_62
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 8188 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_79
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_88
timestamp 1586364061
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_104
timestamp 1586364061
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_108
timestamp 1586364061
transform 1 0 11040 0 -1 25568
box -38 -48 406 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_115
timestamp 1586364061
transform 1 0 11684 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_119
timestamp 1586364061
transform 1 0 12052 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_131
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_42_143
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4784 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 4416 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_35
timestamp 1586364061
transform 1 0 4324 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_38
timestamp 1586364061
transform 1 0 4600 0 1 25568
box -38 -48 222 592
use scs8hd_or2_4  _129_
timestamp 1586364061
transform 1 0 5336 0 1 25568
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 5152 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_42
timestamp 1586364061
transform 1 0 4968 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_53
timestamp 1586364061
transform 1 0 5980 0 1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 774 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 7728 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 7544 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 8740 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_81
timestamp 1586364061
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_85
timestamp 1586364061
transform 1 0 8924 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_100
timestamp 1586364061
transform 1 0 10304 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_104
timestamp 1586364061
transform 1 0 10672 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_108
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_114
timestamp 1586364061
transform 1 0 11592 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_118
timestamp 1586364061
transform 1 0 11960 0 1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_43_121
timestamp 1586364061
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 4784 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 5796 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_49
timestamp 1586364061
transform 1 0 5612 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_53
timestamp 1586364061
transform 1 0 5980 0 -1 26656
box -38 -48 406 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 6348 0 -1 26656
box -38 -48 866 592
use scs8hd_decap_6  FILLER_44_66
timestamp 1586364061
transform 1 0 7176 0 -1 26656
box -38 -48 590 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 8004 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7728 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_74
timestamp 1586364061
transform 1 0 7912 0 -1 26656
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_84
timestamp 1586364061
transform 1 0 8832 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_88
timestamp 1586364061
transform 1 0 9200 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_44_91
timestamp 1586364061
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_98
timestamp 1586364061
transform 1 0 10120 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_111
timestamp 1586364061
transform 1 0 11316 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_115
timestamp 1586364061
transform 1 0 11684 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_122
timestamp 1586364061
transform 1 0 12328 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_134
timestamp 1586364061
transform 1 0 13432 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 4784 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 4140 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_35
timestamp 1586364061
transform 1 0 4324 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_53
timestamp 1586364061
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 7360 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_65
timestamp 1586364061
transform 1 0 7084 0 1 26656
box -38 -48 314 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 7728 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_70
timestamp 1586364061
transform 1 0 7544 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_83
timestamp 1586364061
transform 1 0 8740 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 8924 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 9292 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_87
timestamp 1586364061
transform 1 0 9108 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_91
timestamp 1586364061
transform 1 0 9476 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_95
timestamp 1586364061
transform 1 0 9844 0 1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 26656
box -38 -48 866 592
use scs8hd_decap_3  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_115
timestamp 1586364061
transform 1 0 11684 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_119
timestamp 1586364061
transform 1 0 12052 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_126
timestamp 1586364061
transform 1 0 12696 0 1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_45_132
timestamp 1586364061
transform 1 0 13248 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_144
timestamp 1586364061
transform 1 0 14352 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_nand2_4  _109_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 3220 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 3404 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_23
timestamp 1586364061
transform 1 0 3220 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_8  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_34
timestamp 1586364061
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 130 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 4140 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_38
timestamp 1586364061
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_36
timestamp 1586364061
transform 1 0 4416 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_40
timestamp 1586364061
transform 1 0 4784 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use scs8hd_nor3_4  _158_
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_53
timestamp 1586364061
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_57
timestamp 1586364061
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_61
timestamp 1586364061
transform 1 0 6716 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_57
timestamp 1586364061
transform 1 0 6348 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 6532 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 6900 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_65
timestamp 1586364061
transform 1 0 7084 0 -1 27744
box -38 -48 774 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 6900 0 1 27744
box -38 -48 866 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 7912 0 -1 27744
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_73
timestamp 1586364061
transform 1 0 7820 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_46_83
timestamp 1586364061
transform 1 0 8740 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_72
timestamp 1586364061
transform 1 0 7728 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_76
timestamp 1586364061
transform 1 0 8096 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 9660 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_87
timestamp 1586364061
transform 1 0 9108 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_91
timestamp 1586364061
transform 1 0 9476 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_95
timestamp 1586364061
transform 1 0 9844 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10212 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_109
timestamp 1586364061
transform 1 0 11132 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_114
timestamp 1586364061
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_118
timestamp 1586364061
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_122
timestamp 1586364061
transform 1 0 12328 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 27744
box -38 -48 866 592
use scs8hd_or2_4  _072_
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 682 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 13248 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_126
timestamp 1586364061
transform 1 0 12696 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_133
timestamp 1586364061
transform 1 0 13340 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_130
timestamp 1586364061
transform 1 0 13064 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_134
timestamp 1586364061
transform 1 0 13432 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_47_138
timestamp 1586364061
transform 1 0 13800 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_8  _162_
timestamp 1586364061
transform 1 0 4692 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_36
timestamp 1586364061
transform 1 0 4416 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_48
timestamp 1586364061
transform 1 0 5520 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_52
timestamp 1586364061
transform 1 0 5888 0 -1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 7268 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_65
timestamp 1586364061
transform 1 0 7084 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_48_69
timestamp 1586364061
transform 1 0 7452 0 -1 28832
box -38 -48 590 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 8004 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_84
timestamp 1586364061
transform 1 0 8832 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 28832
box -38 -48 866 592
use scs8hd_fill_1  FILLER_48_97
timestamp 1586364061
transform 1 0 10028 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_107
timestamp 1586364061
transform 1 0 10948 0 -1 28832
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 28832
box -38 -48 866 592
use scs8hd_decap_8  FILLER_48_124
timestamp 1586364061
transform 1 0 12512 0 -1 28832
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_135
timestamp 1586364061
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_143
timestamp 1586364061
transform 1 0 14260 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_19
timestamp 1586364061
transform 1 0 2852 0 1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_49_22
timestamp 1586364061
transform 1 0 3128 0 1 28832
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_33
timestamp 1586364061
transform 1 0 4140 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_37
timestamp 1586364061
transform 1 0 4508 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_50
timestamp 1586364061
transform 1 0 5704 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_54
timestamp 1586364061
transform 1 0 6072 0 1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8556 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_71
timestamp 1586364061
transform 1 0 7636 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_77
timestamp 1586364061
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_92
timestamp 1586364061
transform 1 0 9568 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_96
timestamp 1586364061
transform 1 0 9936 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_109
timestamp 1586364061
transform 1 0 11132 0 1 28832
box -38 -48 1142 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_fill_1  FILLER_49_121
timestamp 1586364061
transform 1 0 12236 0 1 28832
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 13248 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_126
timestamp 1586364061
transform 1 0 12696 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_130
timestamp 1586364061
transform 1 0 13064 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_137
timestamp 1586364061
transform 1 0 13708 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_141
timestamp 1586364061
transform 1 0 14076 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_145
timestamp 1586364061
transform 1 0 14444 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_19
timestamp 1586364061
transform 1 0 2852 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_23
timestamp 1586364061
transform 1 0 3220 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_36
timestamp 1586364061
transform 1 0 4416 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_48
timestamp 1586364061
transform 1 0 5520 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_52
timestamp 1586364061
transform 1 0 5888 0 -1 29920
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_58
timestamp 1586364061
transform 1 0 6440 0 -1 29920
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 8372 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_71
timestamp 1586364061
transform 1 0 7636 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_75
timestamp 1586364061
transform 1 0 8004 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_8  FILLER_50_82
timestamp 1586364061
transform 1 0 8648 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 29920
box -38 -48 222 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 11224 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_102
timestamp 1586364061
transform 1 0 10488 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_106
timestamp 1586364061
transform 1 0 10856 0 -1 29920
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_8  FILLER_50_113
timestamp 1586364061
transform 1 0 11500 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_12  FILLER_50_124
timestamp 1586364061
transform 1 0 12512 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_136
timestamp 1586364061
transform 1 0 13616 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_144
timestamp 1586364061
transform 1 0 14352 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 222 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 3956 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_34
timestamp 1586364061
transform 1 0 4232 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_40
timestamp 1586364061
transform 1 0 4784 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 29920
box -38 -48 866 592
use scs8hd_decap_4  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_55
timestamp 1586364061
transform 1 0 6164 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 6256 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_58
timestamp 1586364061
transform 1 0 6440 0 1 29920
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_73
timestamp 1586364061
transform 1 0 7820 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_77
timestamp 1586364061
transform 1 0 8188 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_81
timestamp 1586364061
transform 1 0 8556 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_85
timestamp 1586364061
transform 1 0 8924 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_89
timestamp 1586364061
transform 1 0 9292 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_104
timestamp 1586364061
transform 1 0 10672 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_108
timestamp 1586364061
transform 1 0 11040 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_114
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_118
timestamp 1586364061
transform 1 0 11960 0 1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 406 592
use scs8hd_inv_8  _161_
timestamp 1586364061
transform 1 0 4600 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 4416 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_53_31
timestamp 1586364061
transform 1 0 3956 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_34
timestamp 1586364061
transform 1 0 4232 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 5612 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_47
timestamp 1586364061
transform 1 0 5428 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_51
timestamp 1586364061
transform 1 0 5796 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_55
timestamp 1586364061
transform 1 0 6164 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_47
timestamp 1586364061
transform 1 0 5428 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_55
timestamp 1586364061
transform 1 0 6164 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_66
timestamp 1586364061
transform 1 0 7176 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_52_67
timestamp 1586364061
transform 1 0 7268 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_63
timestamp 1586364061
transform 1 0 6900 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7084 0 -1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 31008
box -38 -48 866 592
use scs8hd_or2_4  _145_
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 682 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_78
timestamp 1586364061
transform 1 0 8280 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_53_83
timestamp 1586364061
transform 1 0 8740 0 1 31008
box -38 -48 314 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 9016 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_84
timestamp 1586364061
transform 1 0 8832 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_88
timestamp 1586364061
transform 1 0 9200 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_95
timestamp 1586364061
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_104
timestamp 1586364061
transform 1 0 10672 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_108
timestamp 1586364061
transform 1 0 11040 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_99
timestamp 1586364061
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_103
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_121
timestamp 1586364061
transform 1 0 12236 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_113
timestamp 1586364061
transform 1 0 11500 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_117
timestamp 1586364061
transform 1 0 11868 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_121
timestamp 1586364061
transform 1 0 12236 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_133
timestamp 1586364061
transform 1 0 13340 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_35
timestamp 1586364061
transform 1 0 4324 0 -1 32096
box -38 -48 774 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 5244 0 -1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_54_43
timestamp 1586364061
transform 1 0 5060 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_54
timestamp 1586364061
transform 1 0 6072 0 -1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_58
timestamp 1586364061
transform 1 0 6440 0 -1 32096
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_71
timestamp 1586364061
transform 1 0 7636 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_75
timestamp 1586364061
transform 1 0 8004 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_79
timestamp 1586364061
transform 1 0 8372 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 9016 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_84
timestamp 1586364061
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_88
timestamp 1586364061
transform 1 0 9200 0 -1 32096
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_106
timestamp 1586364061
transform 1 0 10856 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_113
timestamp 1586364061
transform 1 0 11500 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_125
timestamp 1586364061
transform 1 0 12604 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_54_137
timestamp 1586364061
transform 1 0 13708 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_36
timestamp 1586364061
transform 1 0 4416 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_40
timestamp 1586364061
transform 1 0 4784 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7360 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_79
timestamp 1586364061
transform 1 0 8372 0 1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_55_83
timestamp 1586364061
transform 1 0 8740 0 1 32096
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_89
timestamp 1586364061
transform 1 0 9292 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_92
timestamp 1586364061
transform 1 0 9568 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_105
timestamp 1586364061
transform 1 0 10764 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_109
timestamp 1586364061
transform 1 0 11132 0 1 32096
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_113
timestamp 1586364061
transform 1 0 11500 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_117
timestamp 1586364061
transform 1 0 11868 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_121
timestamp 1586364061
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_126
timestamp 1586364061
transform 1 0 12696 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_130
timestamp 1586364061
transform 1 0 13064 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_134
timestamp 1586364061
transform 1 0 13432 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_56_29
timestamp 1586364061
transform 1 0 3772 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_56_38
timestamp 1586364061
transform 1 0 4600 0 -1 33184
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 5520 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_42
timestamp 1586364061
transform 1 0 4968 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_46
timestamp 1586364061
transform 1 0 5336 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_61
timestamp 1586364061
transform 1 0 6716 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_65
timestamp 1586364061
transform 1 0 7084 0 -1 33184
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_3  FILLER_56_70
timestamp 1586364061
transform 1 0 7544 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_82
timestamp 1586364061
transform 1 0 8648 0 -1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_86
timestamp 1586364061
transform 1 0 9016 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_2  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 33184
box -38 -48 866 592
use scs8hd_fill_1  FILLER_56_97
timestamp 1586364061
transform 1 0 10028 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_107
timestamp 1586364061
transform 1 0 10948 0 -1 33184
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_111
timestamp 1586364061
transform 1 0 11316 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_114
timestamp 1586364061
transform 1 0 11592 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_124
timestamp 1586364061
transform 1 0 12512 0 -1 33184
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_135
timestamp 1586364061
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_143
timestamp 1586364061
transform 1 0 14260 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 3404 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_23
timestamp 1586364061
transform 1 0 3220 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_36
timestamp 1586364061
transform 1 0 4416 0 1 33184
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 5152 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_42
timestamp 1586364061
transform 1 0 4968 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_53
timestamp 1586364061
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8740 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_71
timestamp 1586364061
transform 1 0 7636 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_75
timestamp 1586364061
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_79
timestamp 1586364061
transform 1 0 8372 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_94
timestamp 1586364061
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_113
timestamp 1586364061
transform 1 0 11500 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_117
timestamp 1586364061
transform 1 0 11868 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_132
timestamp 1586364061
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_136
timestamp 1586364061
transform 1 0 13616 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_144
timestamp 1586364061
transform 1 0 14352 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 5244 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_43
timestamp 1586364061
transform 1 0 5060 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_47
timestamp 1586364061
transform 1 0 5428 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_62
timestamp 1586364061
transform 1 0 6808 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_66
timestamp 1586364061
transform 1 0 7176 0 -1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8648 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_79
timestamp 1586364061
transform 1 0 8372 0 -1 34272
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_84
timestamp 1586364061
transform 1 0 8832 0 -1 34272
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_104
timestamp 1586364061
transform 1 0 10672 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_108
timestamp 1586364061
transform 1 0 11040 0 -1 34272
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_121
timestamp 1586364061
transform 1 0 12236 0 -1 34272
box -38 -48 222 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 13340 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_58_125
timestamp 1586364061
transform 1 0 12604 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_8  FILLER_58_137
timestamp 1586364061
transform 1 0 13708 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 590 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_36
timestamp 1586364061
transform 1 0 4416 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_40
timestamp 1586364061
transform 1 0 4784 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 5152 0 1 34272
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 4968 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_53
timestamp 1586364061
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_46
timestamp 1586364061
transform 1 0 5336 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_50
timestamp 1586364061
transform 1 0 5704 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_6  FILLER_60_54
timestamp 1586364061
transform 1 0 6072 0 -1 35360
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_57
timestamp 1586364061
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8648 0 1 34272
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_73
timestamp 1586364061
transform 1 0 7820 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_78
timestamp 1586364061
transform 1 0 8280 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_71
timestamp 1586364061
transform 1 0 7636 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_60_75
timestamp 1586364061
transform 1 0 8004 0 -1 35360
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_93
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_84
timestamp 1586364061
transform 1 0 8832 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_1  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_97
timestamp 1586364061
transform 1 0 10028 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_110
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_103
timestamp 1586364061
transform 1 0 10580 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_60_107
timestamp 1586364061
transform 1 0 10948 0 -1 35360
box -38 -48 590 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 11500 0 -1 35360
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 11500 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_59_115
timestamp 1586364061
transform 1 0 11684 0 1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_59_121
timestamp 1586364061
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 13432 0 1 34272
box -38 -48 406 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 12696 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 13248 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_126
timestamp 1586364061
transform 1 0 12696 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_130
timestamp 1586364061
transform 1 0 13064 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_138
timestamp 1586364061
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_125
timestamp 1586364061
transform 1 0 12604 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_130
timestamp 1586364061
transform 1 0 13064 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_142
timestamp 1586364061
transform 1 0 14168 0 1 34272
box -38 -48 406 592
use scs8hd_decap_4  FILLER_60_142
timestamp 1586364061
transform 1 0 14168 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_57
timestamp 1586364061
transform 1 0 6348 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 8648 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 8464 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_78
timestamp 1586364061
transform 1 0 8280 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_91
timestamp 1586364061
transform 1 0 9476 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_95
timestamp 1586364061
transform 1 0 9844 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 10764 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_103
timestamp 1586364061
transform 1 0 10580 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_107
timestamp 1586364061
transform 1 0 10948 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 35360
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 11776 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_114
timestamp 1586364061
transform 1 0 11592 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_118
timestamp 1586364061
transform 1 0 11960 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 12972 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_127
timestamp 1586364061
transform 1 0 12788 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_131
timestamp 1586364061
transform 1 0 13156 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 36448
box -38 -48 866 592
use scs8hd_decap_8  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_62_64
timestamp 1586364061
transform 1 0 6992 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 8648 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_74
timestamp 1586364061
transform 1 0 7912 0 -1 36448
box -38 -48 774 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_84
timestamp 1586364061
transform 1 0 8832 0 -1 36448
box -38 -48 774 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 11224 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_97
timestamp 1586364061
transform 1 0 10028 0 -1 36448
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_62_109
timestamp 1586364061
transform 1 0 11132 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_114
timestamp 1586364061
transform 1 0 11592 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_126
timestamp 1586364061
transform 1 0 12696 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_62_138
timestamp 1586364061
transform 1 0 13800 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_66
timestamp 1586364061
transform 1 0 7176 0 1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 8004 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 7820 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_70
timestamp 1586364061
transform 1 0 7544 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_84
timestamp 1586364061
transform 1 0 8832 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_96
timestamp 1586364061
transform 1 0 9936 0 1 36448
box -38 -48 774 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 10764 0 1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_63_104
timestamp 1586364061
transform 1 0 10672 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_109
timestamp 1586364061
transform 1 0 11132 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 11316 0 1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_63_113
timestamp 1586364061
transform 1 0 11500 0 1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_63_121
timestamp 1586364061
transform 1 0 12236 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_64_77
timestamp 1586364061
transform 1 0 8188 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_89
timestamp 1586364061
transform 1 0 9292 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal2 s 5814 39520 5870 40000 6 address[0]
port 0 nsew default input
rlabel metal2 s 6366 39520 6422 40000 6 address[1]
port 1 nsew default input
rlabel metal2 s 7010 39520 7066 40000 6 address[2]
port 2 nsew default input
rlabel metal2 s 7654 39520 7710 40000 6 address[3]
port 3 nsew default input
rlabel metal2 s 8298 39520 8354 40000 6 address[4]
port 4 nsew default input
rlabel metal2 s 8850 39520 8906 40000 6 address[5]
port 5 nsew default input
rlabel metal2 s 9494 39520 9550 40000 6 address[6]
port 6 nsew default input
rlabel metal2 s 386 0 442 480 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 1214 0 1270 480 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 2042 0 2098 480 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 6274 0 6330 480 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal2 s 294 39520 350 40000 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 846 39520 902 40000 6 chany_top_in[1]
port 26 nsew default input
rlabel metal2 s 1490 39520 1546 40000 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_in[3]
port 28 nsew default input
rlabel metal2 s 2686 39520 2742 40000 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_in[5]
port 30 nsew default input
rlabel metal2 s 3974 39520 4030 40000 6 chany_top_in[6]
port 31 nsew default input
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_in[7]
port 32 nsew default input
rlabel metal2 s 5170 39520 5226 40000 6 chany_top_in[8]
port 33 nsew default input
rlabel metal2 s 10690 39520 10746 40000 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal2 s 11978 39520 12034 40000 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal2 s 13174 39520 13230 40000 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 13818 39520 13874 40000 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 14370 39520 14426 40000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal2 s 15014 39520 15070 40000 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal2 s 15658 39520 15714 40000 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal2 s 10138 39520 10194 40000 6 data_in
port 43 nsew default input
rlabel metal2 s 7930 0 7986 480 6 enable
port 44 nsew default input
rlabel metal3 s 0 6672 480 6792 6 left_grid_pin_1_
port 45 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 left_grid_pin_5_
port 46 nsew default tristate
rlabel metal3 s 0 33328 480 33448 6 left_grid_pin_9_
port 47 nsew default tristate
rlabel metal3 s 15520 2456 16000 2576 6 right_grid_pin_0_
port 48 nsew default tristate
rlabel metal3 s 15520 27344 16000 27464 6 right_grid_pin_10_
port 49 nsew default tristate
rlabel metal3 s 15520 32376 16000 32496 6 right_grid_pin_12_
port 50 nsew default tristate
rlabel metal3 s 15520 37408 16000 37528 6 right_grid_pin_14_
port 51 nsew default tristate
rlabel metal3 s 15520 7352 16000 7472 6 right_grid_pin_2_
port 52 nsew default tristate
rlabel metal3 s 15520 12384 16000 12504 6 right_grid_pin_4_
port 53 nsew default tristate
rlabel metal3 s 15520 17416 16000 17536 6 right_grid_pin_6_
port 54 nsew default tristate
rlabel metal3 s 15520 22448 16000 22568 6 right_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 56 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 57 nsew default input
<< end >>
