magic
tech sky130A
magscale 1 2
timestamp 1606931228
<< locali >>
rect 12391 19261 12483 19295
rect 12449 19227 12483 19261
rect 12541 15895 12575 16201
rect 12173 14807 12207 14909
rect 5825 13311 5859 13413
rect 11989 11543 12023 11849
rect 15669 11611 15703 11781
rect 4905 8279 4939 8381
rect 8217 7871 8251 8041
<< viali >>
rect 1961 20009 1995 20043
rect 4537 20009 4571 20043
rect 5181 20009 5215 20043
rect 5641 20009 5675 20043
rect 9137 20009 9171 20043
rect 14013 20009 14047 20043
rect 14565 20009 14599 20043
rect 16221 20009 16255 20043
rect 16773 20009 16807 20043
rect 17325 20009 17359 20043
rect 18521 20009 18555 20043
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 3525 19873 3559 19907
rect 4445 19873 4479 19907
rect 5549 19873 5583 19907
rect 9045 19873 9079 19907
rect 10149 19873 10183 19907
rect 13093 19873 13127 19907
rect 13829 19873 13863 19907
rect 14381 19873 14415 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 16589 19873 16623 19907
rect 17141 19873 17175 19907
rect 17693 19873 17727 19907
rect 18337 19873 18371 19907
rect 4721 19805 4755 19839
rect 5825 19805 5859 19839
rect 9321 19805 9355 19839
rect 10241 19805 10275 19839
rect 10425 19805 10459 19839
rect 13369 19805 13403 19839
rect 2513 19737 2547 19771
rect 8677 19737 8711 19771
rect 15669 19737 15703 19771
rect 17877 19737 17911 19771
rect 4077 19669 4111 19703
rect 9781 19669 9815 19703
rect 2421 19329 2455 19363
rect 20361 19329 20395 19363
rect 1685 19261 1719 19295
rect 2237 19261 2271 19295
rect 3249 19261 3283 19295
rect 5089 19261 5123 19295
rect 7665 19261 7699 19295
rect 9413 19261 9447 19295
rect 9873 19261 9907 19295
rect 11805 19261 11839 19295
rect 12357 19261 12391 19295
rect 12633 19261 12667 19295
rect 13369 19261 13403 19295
rect 13645 19261 13679 19295
rect 14105 19261 14139 19295
rect 14657 19261 14691 19295
rect 15577 19261 15611 19295
rect 16313 19261 16347 19295
rect 17233 19261 17267 19295
rect 18061 19261 18095 19295
rect 18337 19261 18371 19295
rect 18797 19261 18831 19295
rect 19349 19261 19383 19295
rect 20177 19261 20211 19295
rect 3516 19193 3550 19227
rect 5356 19193 5390 19227
rect 7932 19193 7966 19227
rect 10140 19193 10174 19227
rect 12449 19193 12483 19227
rect 12909 19193 12943 19227
rect 14933 19193 14967 19227
rect 15853 19193 15887 19227
rect 17509 19193 17543 19227
rect 1869 19125 1903 19159
rect 4629 19125 4663 19159
rect 6469 19125 6503 19159
rect 9045 19125 9079 19159
rect 11253 19125 11287 19159
rect 11989 19125 12023 19159
rect 14289 19125 14323 19159
rect 16497 19125 16531 19159
rect 18981 19125 19015 19159
rect 19533 19125 19567 19159
rect 1593 18921 1627 18955
rect 4077 18921 4111 18955
rect 4537 18921 4571 18955
rect 6837 18921 6871 18955
rect 13001 18921 13035 18955
rect 15853 18921 15887 18955
rect 2237 18853 2271 18887
rect 5724 18853 5758 18887
rect 12173 18853 12207 18887
rect 13461 18853 13495 18887
rect 14289 18853 14323 18887
rect 16681 18853 16715 18887
rect 17785 18853 17819 18887
rect 18521 18853 18555 18887
rect 1409 18785 1443 18819
rect 1961 18785 1995 18819
rect 3341 18785 3375 18819
rect 3433 18785 3467 18819
rect 4445 18785 4479 18819
rect 7205 18785 7239 18819
rect 8033 18785 8067 18819
rect 8677 18785 8711 18819
rect 10324 18785 10358 18819
rect 11897 18785 11931 18819
rect 13369 18785 13403 18819
rect 14013 18785 14047 18819
rect 15761 18785 15795 18819
rect 16405 18785 16439 18819
rect 17509 18785 17543 18819
rect 18245 18785 18279 18819
rect 3525 18717 3559 18751
rect 4629 18717 4663 18751
rect 5457 18717 5491 18751
rect 8125 18717 8159 18751
rect 8217 18717 8251 18751
rect 8861 18717 8895 18751
rect 10057 18717 10091 18751
rect 13645 18717 13679 18751
rect 15945 18717 15979 18751
rect 2973 18581 3007 18615
rect 7665 18581 7699 18615
rect 11437 18581 11471 18615
rect 15393 18581 15427 18615
rect 5273 18377 5307 18411
rect 8217 18377 8251 18411
rect 11253 18377 11287 18411
rect 14289 18377 14323 18411
rect 16681 18377 16715 18411
rect 17601 18377 17635 18411
rect 5917 18241 5951 18275
rect 7297 18241 7331 18275
rect 8769 18241 8803 18275
rect 12449 18241 12483 18275
rect 14933 18241 14967 18275
rect 18337 18241 18371 18275
rect 1593 18173 1627 18207
rect 2145 18173 2179 18207
rect 2973 18173 3007 18207
rect 7113 18173 7147 18207
rect 8677 18173 8711 18207
rect 9873 18173 9907 18207
rect 12716 18173 12750 18207
rect 14657 18173 14691 18207
rect 15301 18173 15335 18207
rect 17417 18173 17451 18207
rect 18061 18173 18095 18207
rect 2421 18105 2455 18139
rect 3240 18105 3274 18139
rect 5641 18105 5675 18139
rect 6285 18105 6319 18139
rect 8585 18105 8619 18139
rect 10140 18105 10174 18139
rect 15568 18105 15602 18139
rect 1777 18037 1811 18071
rect 4353 18037 4387 18071
rect 5733 18037 5767 18071
rect 13829 18037 13863 18071
rect 14749 18037 14783 18071
rect 1593 17833 1627 17867
rect 3341 17833 3375 17867
rect 6745 17833 6779 17867
rect 10149 17833 10183 17867
rect 12081 17833 12115 17867
rect 15301 17833 15335 17867
rect 15669 17833 15703 17867
rect 17417 17833 17451 17867
rect 13360 17765 13394 17799
rect 1409 17697 1443 17731
rect 1961 17697 1995 17731
rect 2685 17697 2719 17731
rect 5365 17697 5399 17731
rect 5632 17697 5666 17731
rect 7021 17697 7055 17731
rect 10057 17697 10091 17731
rect 12449 17697 12483 17731
rect 15761 17697 15795 17731
rect 17785 17697 17819 17731
rect 18429 17697 18463 17731
rect 2145 17629 2179 17663
rect 7205 17629 7239 17663
rect 10333 17629 10367 17663
rect 12541 17629 12575 17663
rect 12725 17629 12759 17663
rect 13093 17629 13127 17663
rect 15945 17629 15979 17663
rect 17877 17629 17911 17663
rect 18061 17629 18095 17663
rect 2881 17493 2915 17527
rect 9689 17493 9723 17527
rect 14473 17493 14507 17527
rect 1593 17289 1627 17323
rect 5641 17289 5675 17323
rect 12449 17289 12483 17323
rect 16957 17289 16991 17323
rect 2145 17153 2179 17187
rect 2973 17153 3007 17187
rect 6101 17153 6135 17187
rect 6193 17153 6227 17187
rect 13001 17153 13035 17187
rect 13461 17153 13495 17187
rect 17417 17153 17451 17187
rect 17601 17153 17635 17187
rect 1409 17085 1443 17119
rect 1961 17085 1995 17119
rect 3240 17085 3274 17119
rect 6009 17085 6043 17119
rect 7481 17085 7515 17119
rect 7748 17085 7782 17119
rect 9689 17085 9723 17119
rect 17325 17085 17359 17119
rect 18061 17085 18095 17119
rect 18317 17085 18351 17119
rect 9956 17017 9990 17051
rect 4353 16949 4387 16983
rect 8861 16949 8895 16983
rect 9229 16949 9263 16983
rect 11069 16949 11103 16983
rect 12817 16949 12851 16983
rect 12909 16949 12943 16983
rect 19441 16949 19475 16983
rect 1685 16745 1719 16779
rect 2881 16745 2915 16779
rect 6377 16745 6411 16779
rect 9689 16745 9723 16779
rect 10057 16745 10091 16779
rect 10149 16745 10183 16779
rect 12541 16745 12575 16779
rect 13553 16745 13587 16779
rect 16681 16745 16715 16779
rect 11152 16677 11186 16711
rect 18144 16677 18178 16711
rect 1501 16609 1535 16643
rect 2063 16609 2097 16643
rect 3249 16609 3283 16643
rect 3341 16609 3375 16643
rect 5264 16609 5298 16643
rect 6653 16609 6687 16643
rect 7380 16609 7414 16643
rect 8953 16609 8987 16643
rect 12909 16609 12943 16643
rect 13921 16609 13955 16643
rect 15557 16609 15591 16643
rect 17877 16609 17911 16643
rect 2237 16541 2271 16575
rect 3525 16541 3559 16575
rect 4997 16541 5031 16575
rect 7113 16541 7147 16575
rect 10241 16541 10275 16575
rect 10885 16541 10919 16575
rect 13001 16541 13035 16575
rect 13185 16541 13219 16575
rect 14013 16541 14047 16575
rect 14197 16541 14231 16575
rect 15301 16541 15335 16575
rect 8493 16405 8527 16439
rect 8769 16405 8803 16439
rect 12265 16405 12299 16439
rect 19257 16405 19291 16439
rect 1961 16201 1995 16235
rect 4261 16201 4295 16235
rect 10425 16201 10459 16235
rect 12541 16201 12575 16235
rect 12633 16201 12667 16235
rect 15025 16201 15059 16235
rect 16037 16201 16071 16235
rect 17693 16201 17727 16235
rect 18061 16201 18095 16235
rect 5273 16133 5307 16167
rect 2605 16065 2639 16099
rect 4721 16065 4755 16099
rect 4813 16065 4847 16099
rect 5825 16065 5859 16099
rect 7941 16065 7975 16099
rect 8125 16065 8159 16099
rect 1777 15997 1811 16031
rect 2872 15997 2906 16031
rect 7849 15997 7883 16031
rect 9045 15997 9079 16031
rect 5641 15929 5675 15963
rect 6285 15929 6319 15963
rect 9312 15929 9346 15963
rect 14749 16133 14783 16167
rect 12909 16065 12943 16099
rect 13369 16065 13403 16099
rect 15577 16065 15611 16099
rect 16313 16065 16347 16099
rect 18705 16065 18739 16099
rect 12817 15997 12851 16031
rect 13636 15997 13670 16031
rect 16221 15997 16255 16031
rect 16580 15929 16614 15963
rect 18521 15929 18555 15963
rect 3985 15861 4019 15895
rect 4629 15861 4663 15895
rect 5733 15861 5767 15895
rect 7481 15861 7515 15895
rect 12541 15861 12575 15895
rect 15393 15861 15427 15895
rect 15485 15861 15519 15895
rect 18429 15861 18463 15895
rect 1593 15657 1627 15691
rect 3249 15657 3283 15691
rect 6193 15657 6227 15691
rect 6469 15657 6503 15691
rect 6837 15657 6871 15691
rect 7297 15657 7331 15691
rect 7849 15657 7883 15691
rect 9045 15657 9079 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 13001 15657 13035 15691
rect 14013 15657 14047 15691
rect 14473 15657 14507 15691
rect 15485 15657 15519 15691
rect 17141 15657 17175 15691
rect 17969 15657 18003 15691
rect 18981 15657 19015 15691
rect 2237 15589 2271 15623
rect 7205 15589 7239 15623
rect 11244 15589 11278 15623
rect 14381 15589 14415 15623
rect 16028 15589 16062 15623
rect 1409 15521 1443 15555
rect 1971 15521 2005 15555
rect 5080 15521 5114 15555
rect 6653 15521 6687 15555
rect 8033 15521 8067 15555
rect 8953 15521 8987 15555
rect 10057 15521 10091 15555
rect 10977 15521 11011 15555
rect 13369 15521 13403 15555
rect 15669 15521 15703 15555
rect 18337 15521 18371 15555
rect 4813 15453 4847 15487
rect 7481 15453 7515 15487
rect 9229 15453 9263 15487
rect 10241 15453 10275 15487
rect 13461 15453 13495 15487
rect 13645 15453 13679 15487
rect 14565 15453 14599 15487
rect 15761 15453 15795 15487
rect 17417 15453 17451 15487
rect 18429 15453 18463 15487
rect 18613 15453 18647 15487
rect 8585 15385 8619 15419
rect 12357 15317 12391 15351
rect 1593 15113 1627 15147
rect 5641 15113 5675 15147
rect 10149 15113 10183 15147
rect 13369 15113 13403 15147
rect 16589 15113 16623 15147
rect 19717 15113 19751 15147
rect 2145 14977 2179 15011
rect 2789 14977 2823 15011
rect 6193 14977 6227 15011
rect 8769 14977 8803 15011
rect 11897 14977 11931 15011
rect 14013 14977 14047 15011
rect 14933 14977 14967 15011
rect 16221 14977 16255 15011
rect 17141 14977 17175 15011
rect 18337 14977 18371 15011
rect 1409 14909 1443 14943
rect 1971 14909 2005 14943
rect 3056 14909 3090 14943
rect 6101 14909 6135 14943
rect 6837 14909 6871 14943
rect 7104 14909 7138 14943
rect 9036 14909 9070 14943
rect 11805 14909 11839 14943
rect 12173 14909 12207 14943
rect 13737 14909 13771 14943
rect 16037 14909 16071 14943
rect 16957 14909 16991 14943
rect 18604 14909 18638 14943
rect 11713 14841 11747 14875
rect 14841 14841 14875 14875
rect 17049 14841 17083 14875
rect 4169 14773 4203 14807
rect 6009 14773 6043 14807
rect 8217 14773 8251 14807
rect 11345 14773 11379 14807
rect 12173 14773 12207 14807
rect 13829 14773 13863 14807
rect 14381 14773 14415 14807
rect 14749 14773 14783 14807
rect 15577 14773 15611 14807
rect 15945 14773 15979 14807
rect 1777 14569 1811 14603
rect 2973 14569 3007 14603
rect 5457 14569 5491 14603
rect 8769 14569 8803 14603
rect 9689 14569 9723 14603
rect 12633 14569 12667 14603
rect 14841 14569 14875 14603
rect 15853 14569 15887 14603
rect 17325 14569 17359 14603
rect 2421 14501 2455 14535
rect 4322 14501 4356 14535
rect 6193 14501 6227 14535
rect 8677 14501 8711 14535
rect 10876 14501 10910 14535
rect 16221 14501 16255 14535
rect 18696 14501 18730 14535
rect 1593 14433 1627 14467
rect 2145 14433 2179 14467
rect 3341 14433 3375 14467
rect 6920 14433 6954 14467
rect 10609 14433 10643 14467
rect 12725 14433 12759 14467
rect 13728 14433 13762 14467
rect 16313 14433 16347 14467
rect 17233 14433 17267 14467
rect 17877 14433 17911 14467
rect 18429 14433 18463 14467
rect 3433 14365 3467 14399
rect 3617 14365 3651 14399
rect 4077 14365 4111 14399
rect 6653 14365 6687 14399
rect 8861 14365 8895 14399
rect 12817 14365 12851 14399
rect 13461 14365 13495 14399
rect 16497 14365 16531 14399
rect 17417 14365 17451 14399
rect 16865 14297 16899 14331
rect 8033 14229 8067 14263
rect 8309 14229 8343 14263
rect 11989 14229 12023 14263
rect 12265 14229 12299 14263
rect 19809 14229 19843 14263
rect 1593 14025 1627 14059
rect 3617 14025 3651 14059
rect 6377 14025 6411 14059
rect 6837 14025 6871 14059
rect 9781 14025 9815 14059
rect 13553 14025 13587 14059
rect 17417 14025 17451 14059
rect 11161 13957 11195 13991
rect 2145 13889 2179 13923
rect 3157 13889 3191 13923
rect 4169 13889 4203 13923
rect 4997 13889 5031 13923
rect 7297 13889 7331 13923
rect 7389 13889 7423 13923
rect 8401 13889 8435 13923
rect 11805 13889 11839 13923
rect 13093 13889 13127 13923
rect 14565 13889 14599 13923
rect 16037 13889 16071 13923
rect 1409 13821 1443 13855
rect 1961 13821 1995 13855
rect 11529 13821 11563 13855
rect 13001 13821 13035 13855
rect 13737 13821 13771 13855
rect 14289 13821 14323 13855
rect 14381 13821 14415 13855
rect 16304 13821 16338 13855
rect 3985 13753 4019 13787
rect 5264 13753 5298 13787
rect 7205 13753 7239 13787
rect 8668 13753 8702 13787
rect 12909 13753 12943 13787
rect 4077 13685 4111 13719
rect 11621 13685 11655 13719
rect 12541 13685 12575 13719
rect 13921 13685 13955 13719
rect 5457 13481 5491 13515
rect 6009 13481 6043 13515
rect 6469 13481 6503 13515
rect 8217 13481 8251 13515
rect 12081 13481 12115 13515
rect 12633 13481 12667 13515
rect 13093 13481 13127 13515
rect 13829 13481 13863 13515
rect 14289 13481 14323 13515
rect 15301 13481 15335 13515
rect 2329 13413 2363 13447
rect 5825 13413 5859 13447
rect 10149 13413 10183 13447
rect 13001 13413 13035 13447
rect 14197 13413 14231 13447
rect 17132 13413 17166 13447
rect 2063 13345 2097 13379
rect 5365 13345 5399 13379
rect 6377 13345 6411 13379
rect 7757 13345 7791 13379
rect 8585 13345 8619 13379
rect 9413 13345 9447 13379
rect 10241 13345 10275 13379
rect 10793 13345 10827 13379
rect 15669 13345 15703 13379
rect 16865 13345 16899 13379
rect 5549 13277 5583 13311
rect 5825 13277 5859 13311
rect 6561 13277 6595 13311
rect 8677 13277 8711 13311
rect 8861 13277 8895 13311
rect 10425 13277 10459 13311
rect 13185 13277 13219 13311
rect 14381 13277 14415 13311
rect 15761 13277 15795 13311
rect 15853 13277 15887 13311
rect 4997 13209 5031 13243
rect 9229 13141 9263 13175
rect 9781 13141 9815 13175
rect 18245 13141 18279 13175
rect 1961 12937 1995 12971
rect 2513 12937 2547 12971
rect 3065 12937 3099 12971
rect 6101 12937 6135 12971
rect 9505 12937 9539 12971
rect 14565 12937 14599 12971
rect 16957 12937 16991 12971
rect 3617 12869 3651 12903
rect 18061 12869 18095 12903
rect 4169 12801 4203 12835
rect 6837 12801 6871 12835
rect 12449 12801 12483 12835
rect 14841 12801 14875 12835
rect 18613 12801 18647 12835
rect 1777 12733 1811 12767
rect 2329 12733 2363 12767
rect 2881 12733 2915 12767
rect 4721 12733 4755 12767
rect 7481 12733 7515 12767
rect 8125 12733 8159 12767
rect 10609 12733 10643 12767
rect 13185 12733 13219 12767
rect 13452 12733 13486 12767
rect 15577 12733 15611 12767
rect 18429 12733 18463 12767
rect 3985 12665 4019 12699
rect 4988 12665 5022 12699
rect 8392 12665 8426 12699
rect 10876 12665 10910 12699
rect 15844 12665 15878 12699
rect 18521 12665 18555 12699
rect 4077 12597 4111 12631
rect 7297 12597 7331 12631
rect 11989 12597 12023 12631
rect 5457 12393 5491 12427
rect 7481 12393 7515 12427
rect 8585 12393 8619 12427
rect 9045 12393 9079 12427
rect 14197 12393 14231 12427
rect 15485 12393 15519 12427
rect 16957 12393 16991 12427
rect 18981 12393 19015 12427
rect 19441 12393 19475 12427
rect 2329 12325 2363 12359
rect 3065 12325 3099 12359
rect 4322 12325 4356 12359
rect 6000 12325 6034 12359
rect 11704 12325 11738 12359
rect 2053 12257 2087 12291
rect 2789 12257 2823 12291
rect 5733 12257 5767 12291
rect 7849 12257 7883 12291
rect 7941 12257 7975 12291
rect 8953 12257 8987 12291
rect 10517 12257 10551 12291
rect 14105 12257 14139 12291
rect 14933 12257 14967 12291
rect 15853 12257 15887 12291
rect 16497 12257 16531 12291
rect 17141 12257 17175 12291
rect 17325 12257 17359 12291
rect 17592 12257 17626 12291
rect 19349 12257 19383 12291
rect 4077 12189 4111 12223
rect 8125 12189 8159 12223
rect 9137 12189 9171 12223
rect 10609 12189 10643 12223
rect 10793 12189 10827 12223
rect 11437 12189 11471 12223
rect 14381 12189 14415 12223
rect 15945 12189 15979 12223
rect 16129 12189 16163 12223
rect 19533 12189 19567 12223
rect 12817 12121 12851 12155
rect 13737 12121 13771 12155
rect 7113 12053 7147 12087
rect 10149 12053 10183 12087
rect 14749 12053 14783 12087
rect 18705 12053 18739 12087
rect 4169 11849 4203 11883
rect 4445 11849 4479 11883
rect 6837 11849 6871 11883
rect 9321 11849 9355 11883
rect 11989 11849 12023 11883
rect 17233 11849 17267 11883
rect 18061 11849 18095 11883
rect 1961 11713 1995 11747
rect 2789 11713 2823 11747
rect 4905 11713 4939 11747
rect 4997 11713 5031 11747
rect 7389 11713 7423 11747
rect 7941 11713 7975 11747
rect 9689 11713 9723 11747
rect 1777 11645 1811 11679
rect 3056 11645 3090 11679
rect 7297 11645 7331 11679
rect 10149 11645 10183 11679
rect 10416 11645 10450 11679
rect 8208 11577 8242 11611
rect 15577 11781 15611 11815
rect 15669 11781 15703 11815
rect 12909 11713 12943 11747
rect 13001 11713 13035 11747
rect 13737 11713 13771 11747
rect 12265 11645 12299 11679
rect 13461 11645 13495 11679
rect 14197 11645 14231 11679
rect 18613 11713 18647 11747
rect 19717 11713 19751 11747
rect 15853 11645 15887 11679
rect 12817 11577 12851 11611
rect 14464 11577 14498 11611
rect 15669 11577 15703 11611
rect 16098 11577 16132 11611
rect 17509 11577 17543 11611
rect 18429 11577 18463 11611
rect 19984 11577 20018 11611
rect 4813 11509 4847 11543
rect 7205 11509 7239 11543
rect 11529 11509 11563 11543
rect 11989 11509 12023 11543
rect 12081 11509 12115 11543
rect 12449 11509 12483 11543
rect 18521 11509 18555 11543
rect 18889 11509 18923 11543
rect 21097 11509 21131 11543
rect 1593 11305 1627 11339
rect 4537 11305 4571 11339
rect 8861 11305 8895 11339
rect 11161 11305 11195 11339
rect 11897 11305 11931 11339
rect 13277 11305 13311 11339
rect 13737 11305 13771 11339
rect 15301 11305 15335 11339
rect 6837 11237 6871 11271
rect 9137 11237 9171 11271
rect 12265 11237 12299 11271
rect 15761 11237 15795 11271
rect 1409 11169 1443 11203
rect 1961 11169 1995 11203
rect 3249 11169 3283 11203
rect 3341 11169 3375 11203
rect 7748 11169 7782 11203
rect 11253 11169 11287 11203
rect 13645 11169 13679 11203
rect 15669 11169 15703 11203
rect 2145 11101 2179 11135
rect 3525 11101 3559 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 7481 11101 7515 11135
rect 11437 11101 11471 11135
rect 12357 11101 12391 11135
rect 12449 11101 12483 11135
rect 13829 11101 13863 11135
rect 15945 11101 15979 11135
rect 6469 11033 6503 11067
rect 10793 11033 10827 11067
rect 2881 10965 2915 10999
rect 2053 10761 2087 10795
rect 14565 10761 14599 10795
rect 3065 10693 3099 10727
rect 8217 10693 8251 10727
rect 8493 10693 8527 10727
rect 11437 10693 11471 10727
rect 2697 10625 2731 10659
rect 3709 10625 3743 10659
rect 4721 10625 4755 10659
rect 6837 10625 6871 10659
rect 9045 10625 9079 10659
rect 10057 10625 10091 10659
rect 12449 10625 12483 10659
rect 18061 10625 18095 10659
rect 2421 10557 2455 10591
rect 2513 10557 2547 10591
rect 4537 10557 4571 10591
rect 6009 10557 6043 10591
rect 9689 10557 9723 10591
rect 10324 10557 10358 10591
rect 13185 10557 13219 10591
rect 15761 10557 15795 10591
rect 18328 10557 18362 10591
rect 7104 10489 7138 10523
rect 8861 10489 8895 10523
rect 8953 10489 8987 10523
rect 13452 10489 13486 10523
rect 16028 10489 16062 10523
rect 3433 10421 3467 10455
rect 3525 10421 3559 10455
rect 4077 10421 4111 10455
rect 4445 10421 4479 10455
rect 5825 10421 5859 10455
rect 9505 10421 9539 10455
rect 14841 10421 14875 10455
rect 17141 10421 17175 10455
rect 17417 10421 17451 10455
rect 19441 10421 19475 10455
rect 3433 10217 3467 10251
rect 5457 10217 5491 10251
rect 12357 10217 12391 10251
rect 14013 10217 14047 10251
rect 15393 10217 15427 10251
rect 8401 10149 8435 10183
rect 11244 10149 11278 10183
rect 12878 10149 12912 10183
rect 15853 10149 15887 10183
rect 16672 10149 16706 10183
rect 2044 10081 2078 10115
rect 4077 10081 4111 10115
rect 4344 10081 4378 10115
rect 5733 10081 5767 10115
rect 6000 10081 6034 10115
rect 8493 10081 8527 10115
rect 10977 10081 11011 10115
rect 15761 10081 15795 10115
rect 16405 10081 16439 10115
rect 1777 10013 1811 10047
rect 8677 10013 8711 10047
rect 12633 10013 12667 10047
rect 16037 10013 16071 10047
rect 3157 9877 3191 9911
rect 7113 9877 7147 9911
rect 8033 9877 8067 9911
rect 17785 9877 17819 9911
rect 3065 9673 3099 9707
rect 4077 9605 4111 9639
rect 5733 9605 5767 9639
rect 10149 9605 10183 9639
rect 10425 9605 10459 9639
rect 14013 9605 14047 9639
rect 16589 9605 16623 9639
rect 3709 9537 3743 9571
rect 4721 9537 4755 9571
rect 6377 9537 6411 9571
rect 7481 9537 7515 9571
rect 10977 9537 11011 9571
rect 14565 9537 14599 9571
rect 17141 9537 17175 9571
rect 3525 9469 3559 9503
rect 6193 9469 6227 9503
rect 8769 9469 8803 9503
rect 9036 9469 9070 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 17049 9469 17083 9503
rect 4445 9401 4479 9435
rect 6101 9401 6135 9435
rect 10885 9401 10919 9435
rect 16957 9401 16991 9435
rect 3433 9333 3467 9367
rect 4537 9333 4571 9367
rect 6837 9333 6871 9367
rect 7205 9333 7239 9367
rect 7297 9333 7331 9367
rect 10793 9333 10827 9367
rect 1961 9129 1995 9163
rect 2513 9129 2547 9163
rect 4629 9129 4663 9163
rect 5181 9129 5215 9163
rect 6377 9129 6411 9163
rect 9689 9129 9723 9163
rect 10149 9061 10183 9095
rect 1777 8993 1811 9027
rect 2329 8993 2363 9027
rect 5089 8993 5123 9027
rect 7941 8993 7975 9027
rect 8208 8993 8242 9027
rect 10057 8993 10091 9027
rect 5273 8925 5307 8959
rect 10241 8925 10275 8959
rect 9321 8857 9355 8891
rect 4721 8789 4755 8823
rect 4077 8517 4111 8551
rect 8493 8517 8527 8551
rect 1685 8449 1719 8483
rect 4629 8449 4663 8483
rect 5641 8449 5675 8483
rect 7113 8449 7147 8483
rect 9321 8449 9355 8483
rect 1409 8381 1443 8415
rect 2145 8381 2179 8415
rect 2412 8381 2446 8415
rect 4537 8381 4571 8415
rect 4905 8381 4939 8415
rect 5549 8381 5583 8415
rect 9137 8381 9171 8415
rect 9229 8381 9263 8415
rect 4445 8313 4479 8347
rect 7380 8313 7414 8347
rect 3525 8245 3559 8279
rect 4905 8245 4939 8279
rect 5089 8245 5123 8279
rect 5457 8245 5491 8279
rect 8769 8245 8803 8279
rect 4537 8041 4571 8075
rect 8125 8041 8159 8075
rect 8217 8041 8251 8075
rect 8861 8041 8895 8075
rect 18613 8041 18647 8075
rect 2329 7973 2363 8007
rect 2042 7905 2076 7939
rect 4445 7905 4479 7939
rect 5356 7905 5390 7939
rect 7012 7905 7046 7939
rect 8769 7905 8803 7939
rect 18435 7905 18469 7939
rect 4721 7837 4755 7871
rect 5089 7837 5123 7871
rect 6745 7837 6779 7871
rect 8217 7837 8251 7871
rect 8953 7837 8987 7871
rect 6469 7769 6503 7803
rect 4077 7701 4111 7735
rect 8401 7701 8435 7735
rect 4353 7497 4387 7531
rect 6009 7497 6043 7531
rect 19165 7497 19199 7531
rect 2973 7361 3007 7395
rect 7849 7361 7883 7395
rect 8769 7361 8803 7395
rect 8953 7361 8987 7395
rect 3240 7293 3274 7327
rect 4629 7293 4663 7327
rect 4885 7293 4919 7327
rect 8677 7293 8711 7327
rect 18981 7293 19015 7327
rect 6837 7225 6871 7259
rect 7665 7225 7699 7259
rect 7297 7157 7331 7191
rect 7757 7157 7791 7191
rect 8309 7157 8343 7191
rect 8585 6953 8619 6987
rect 8677 6885 8711 6919
rect 4445 6817 4479 6851
rect 5089 6817 5123 6851
rect 7481 6817 7515 6851
rect 7573 6817 7607 6851
rect 19441 6817 19475 6851
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 7757 6749 7791 6783
rect 8861 6749 8895 6783
rect 4077 6681 4111 6715
rect 8217 6681 8251 6715
rect 19625 6681 19659 6715
rect 7113 6613 7147 6647
rect 20085 6409 20119 6443
rect 19901 6205 19935 6239
rect 20453 5865 20487 5899
rect 20269 5729 20303 5763
rect 20729 5321 20763 5355
rect 20545 5117 20579 5151
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2866 20040 2872 20052
rect 1995 20012 2872 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 5169 20043 5227 20049
rect 5169 20040 5181 20043
rect 4571 20012 5181 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 5169 20009 5181 20012
rect 5215 20009 5227 20043
rect 5626 20040 5632 20052
rect 5587 20012 5632 20040
rect 5169 20003 5227 20009
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9306 20040 9312 20052
rect 9171 20012 9312 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9306 20000 9312 20012
rect 9364 20000 9370 20052
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 14001 20043 14059 20049
rect 14001 20040 14013 20043
rect 12952 20012 14013 20040
rect 12952 20000 12958 20012
rect 14001 20009 14013 20012
rect 14047 20009 14059 20043
rect 14001 20003 14059 20009
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 14332 20012 14565 20040
rect 14332 20000 14338 20012
rect 14553 20009 14565 20012
rect 14599 20009 14611 20043
rect 14553 20003 14611 20009
rect 15654 20000 15660 20052
rect 15712 20040 15718 20052
rect 16209 20043 16267 20049
rect 16209 20040 16221 20043
rect 15712 20012 16221 20040
rect 15712 20000 15718 20012
rect 16209 20009 16221 20012
rect 16255 20009 16267 20043
rect 16209 20003 16267 20009
rect 16298 20000 16304 20052
rect 16356 20040 16362 20052
rect 16761 20043 16819 20049
rect 16761 20040 16773 20043
rect 16356 20012 16773 20040
rect 16356 20000 16362 20012
rect 16761 20009 16773 20012
rect 16807 20009 16819 20043
rect 16761 20003 16819 20009
rect 16850 20000 16856 20052
rect 16908 20040 16914 20052
rect 17313 20043 17371 20049
rect 17313 20040 17325 20043
rect 16908 20012 17325 20040
rect 16908 20000 16914 20012
rect 17313 20009 17325 20012
rect 17359 20009 17371 20043
rect 17313 20003 17371 20009
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18472 20012 18521 20040
rect 18472 20000 18478 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18509 20003 18567 20009
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 3513 19907 3571 19913
rect 3513 19873 3525 19907
rect 3559 19904 3571 19907
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3559 19876 4445 19904
rect 3559 19873 3571 19876
rect 3513 19867 3571 19873
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 5537 19907 5595 19913
rect 5537 19873 5549 19907
rect 5583 19904 5595 19907
rect 5994 19904 6000 19916
rect 5583 19876 6000 19904
rect 5583 19873 5595 19876
rect 5537 19867 5595 19873
rect 5994 19864 6000 19876
rect 6052 19904 6058 19916
rect 9033 19907 9091 19913
rect 9033 19904 9045 19907
rect 6052 19876 9045 19904
rect 6052 19864 6058 19876
rect 9033 19873 9045 19876
rect 9079 19873 9091 19907
rect 9033 19867 9091 19873
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9732 19876 10149 19904
rect 9732 19864 9738 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 13078 19904 13084 19916
rect 13039 19876 13084 19904
rect 10137 19867 10195 19873
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 13814 19904 13820 19916
rect 13775 19876 13820 19904
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 14369 19907 14427 19913
rect 14369 19873 14381 19907
rect 14415 19873 14427 19907
rect 14369 19867 14427 19873
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4890 19836 4896 19848
rect 4755 19808 4896 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 5810 19836 5816 19848
rect 5771 19808 5816 19836
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 10042 19836 10048 19848
rect 9355 19808 10048 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 10042 19796 10048 19808
rect 10100 19796 10106 19848
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 10413 19839 10471 19845
rect 10413 19805 10425 19839
rect 10459 19836 10471 19839
rect 10962 19836 10968 19848
rect 10459 19808 10968 19836
rect 10459 19805 10471 19808
rect 10413 19799 10471 19805
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19768 2559 19771
rect 2774 19768 2780 19780
rect 2547 19740 2780 19768
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 2774 19728 2780 19740
rect 2832 19728 2838 19780
rect 8665 19771 8723 19777
rect 8665 19737 8677 19771
rect 8711 19768 8723 19771
rect 10244 19768 10272 19799
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 14090 19836 14096 19848
rect 13403 19808 14096 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 8711 19740 10272 19768
rect 8711 19737 8723 19740
rect 8665 19731 8723 19737
rect 13262 19728 13268 19780
rect 13320 19768 13326 19780
rect 14384 19768 14412 19867
rect 15378 19864 15384 19916
rect 15436 19904 15442 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 15436 19876 15485 19904
rect 15436 19864 15442 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 16025 19907 16083 19913
rect 16025 19904 16037 19907
rect 15712 19876 16037 19904
rect 15712 19864 15718 19876
rect 16025 19873 16037 19876
rect 16071 19873 16083 19907
rect 16574 19904 16580 19916
rect 16535 19876 16580 19904
rect 16025 19867 16083 19873
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 16666 19864 16672 19916
rect 16724 19904 16730 19916
rect 17129 19907 17187 19913
rect 17129 19904 17141 19907
rect 16724 19876 17141 19904
rect 16724 19864 16730 19876
rect 17129 19873 17141 19876
rect 17175 19873 17187 19907
rect 17129 19867 17187 19873
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18506 19904 18512 19916
rect 18371 19876 18512 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 17696 19836 17724 19867
rect 18506 19864 18512 19876
rect 18564 19864 18570 19916
rect 18598 19836 18604 19848
rect 17696 19808 18604 19836
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 13320 19740 14412 19768
rect 13320 19728 13326 19740
rect 15194 19728 15200 19780
rect 15252 19768 15258 19780
rect 15657 19771 15715 19777
rect 15657 19768 15669 19771
rect 15252 19740 15669 19768
rect 15252 19728 15258 19740
rect 15657 19737 15669 19740
rect 15703 19737 15715 19771
rect 15657 19731 15715 19737
rect 17034 19728 17040 19780
rect 17092 19768 17098 19780
rect 17865 19771 17923 19777
rect 17865 19768 17877 19771
rect 17092 19740 17877 19768
rect 17092 19728 17098 19740
rect 17865 19737 17877 19740
rect 17911 19737 17923 19771
rect 17865 19731 17923 19737
rect 2222 19660 2228 19712
rect 2280 19700 2286 19712
rect 4065 19703 4123 19709
rect 4065 19700 4077 19703
rect 2280 19672 4077 19700
rect 2280 19660 2286 19672
rect 4065 19669 4077 19672
rect 4111 19669 4123 19703
rect 9766 19700 9772 19712
rect 9727 19672 9772 19700
rect 4065 19663 4123 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 3108 19468 4844 19496
rect 3108 19456 3114 19468
rect 1762 19320 1768 19372
rect 1820 19360 1826 19372
rect 2409 19363 2467 19369
rect 2409 19360 2421 19363
rect 1820 19332 2421 19360
rect 1820 19320 1826 19332
rect 2409 19329 2421 19332
rect 2455 19329 2467 19363
rect 4816 19360 4844 19468
rect 20346 19360 20352 19372
rect 4816 19332 5212 19360
rect 20307 19332 20352 19360
rect 2409 19323 2467 19329
rect 1670 19292 1676 19304
rect 1631 19264 1676 19292
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19261 3295 19295
rect 3237 19255 3295 19261
rect 198 19184 204 19236
rect 256 19224 262 19236
rect 3050 19224 3056 19236
rect 256 19196 3056 19224
rect 256 19184 262 19196
rect 3050 19184 3056 19196
rect 3108 19184 3114 19236
rect 1857 19159 1915 19165
rect 1857 19125 1869 19159
rect 1903 19156 1915 19159
rect 2958 19156 2964 19168
rect 1903 19128 2964 19156
rect 1903 19125 1915 19128
rect 1857 19119 1915 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3252 19156 3280 19255
rect 4982 19252 4988 19304
rect 5040 19292 5046 19304
rect 5077 19295 5135 19301
rect 5077 19292 5089 19295
rect 5040 19264 5089 19292
rect 5040 19252 5046 19264
rect 5077 19261 5089 19264
rect 5123 19261 5135 19295
rect 5184 19292 5212 19332
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 7650 19292 7656 19304
rect 5184 19264 7512 19292
rect 7611 19264 7656 19292
rect 5077 19255 5135 19261
rect 3504 19227 3562 19233
rect 3504 19193 3516 19227
rect 3550 19224 3562 19227
rect 5344 19227 5402 19233
rect 3550 19196 4936 19224
rect 3550 19193 3562 19196
rect 3504 19187 3562 19193
rect 4908 19168 4936 19196
rect 5344 19193 5356 19227
rect 5390 19224 5402 19227
rect 5810 19224 5816 19236
rect 5390 19196 5816 19224
rect 5390 19193 5402 19196
rect 5344 19187 5402 19193
rect 5810 19184 5816 19196
rect 5868 19224 5874 19236
rect 6822 19224 6828 19236
rect 5868 19196 6828 19224
rect 5868 19184 5874 19196
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 7484 19224 7512 19264
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 9401 19295 9459 19301
rect 7852 19264 9352 19292
rect 7852 19224 7880 19264
rect 7484 19196 7880 19224
rect 7920 19227 7978 19233
rect 7920 19193 7932 19227
rect 7966 19224 7978 19227
rect 8754 19224 8760 19236
rect 7966 19196 8760 19224
rect 7966 19193 7978 19196
rect 7920 19187 7978 19193
rect 8754 19184 8760 19196
rect 8812 19184 8818 19236
rect 3418 19156 3424 19168
rect 3252 19128 3424 19156
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 3602 19116 3608 19168
rect 3660 19156 3666 19168
rect 4062 19156 4068 19168
rect 3660 19128 4068 19156
rect 3660 19116 3666 19128
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4617 19159 4675 19165
rect 4617 19156 4629 19159
rect 4212 19128 4629 19156
rect 4212 19116 4218 19128
rect 4617 19125 4629 19128
rect 4663 19125 4675 19159
rect 4617 19119 4675 19125
rect 4890 19116 4896 19168
rect 4948 19156 4954 19168
rect 6457 19159 6515 19165
rect 6457 19156 6469 19159
rect 4948 19128 6469 19156
rect 4948 19116 4954 19128
rect 6457 19125 6469 19128
rect 6503 19125 6515 19159
rect 6457 19119 6515 19125
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 9033 19159 9091 19165
rect 9033 19156 9045 19159
rect 8260 19128 9045 19156
rect 8260 19116 8266 19128
rect 9033 19125 9045 19128
rect 9079 19125 9091 19159
rect 9324 19156 9352 19264
rect 9401 19261 9413 19295
rect 9447 19292 9459 19295
rect 9674 19292 9680 19304
rect 9447 19264 9680 19292
rect 9447 19261 9459 19264
rect 9401 19255 9459 19261
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19292 9919 19295
rect 9950 19292 9956 19304
rect 9907 19264 9956 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 9950 19252 9956 19264
rect 10008 19252 10014 19304
rect 11793 19295 11851 19301
rect 11793 19261 11805 19295
rect 11839 19292 11851 19295
rect 12345 19295 12403 19301
rect 12345 19292 12357 19295
rect 11839 19264 12357 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 12345 19261 12357 19264
rect 12391 19261 12403 19295
rect 12618 19292 12624 19304
rect 12579 19264 12624 19292
rect 12345 19255 12403 19261
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 13354 19292 13360 19304
rect 13315 19264 13360 19292
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 13814 19292 13820 19304
rect 13679 19264 13820 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 14090 19292 14096 19304
rect 14051 19264 14096 19292
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14366 19252 14372 19304
rect 14424 19292 14430 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 14424 19264 14657 19292
rect 14424 19252 14430 19264
rect 14645 19261 14657 19264
rect 14691 19261 14703 19295
rect 15562 19292 15568 19304
rect 15523 19264 15568 19292
rect 14645 19255 14703 19261
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 16298 19292 16304 19304
rect 16259 19264 16304 19292
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 16850 19252 16856 19304
rect 16908 19292 16914 19304
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 16908 19264 17233 19292
rect 16908 19252 16914 19264
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 18012 19264 18061 19292
rect 18012 19252 18018 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19292 18383 19295
rect 18785 19295 18843 19301
rect 18785 19292 18797 19295
rect 18371 19264 18797 19292
rect 18371 19261 18383 19264
rect 18325 19255 18383 19261
rect 18785 19261 18797 19264
rect 18831 19261 18843 19295
rect 18785 19255 18843 19261
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19024 19264 19349 19292
rect 19024 19252 19030 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19337 19255 19395 19261
rect 20165 19295 20223 19301
rect 20165 19261 20177 19295
rect 20211 19292 20223 19295
rect 22094 19292 22100 19304
rect 20211 19264 22100 19292
rect 20211 19261 20223 19264
rect 20165 19255 20223 19261
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 10134 19233 10140 19236
rect 10128 19224 10140 19233
rect 10095 19196 10140 19224
rect 10128 19187 10140 19196
rect 10134 19184 10140 19187
rect 10192 19184 10198 19236
rect 12066 19224 12072 19236
rect 10244 19196 12072 19224
rect 10244 19156 10272 19196
rect 12066 19184 12072 19196
rect 12124 19184 12130 19236
rect 12437 19227 12495 19233
rect 12437 19193 12449 19227
rect 12483 19224 12495 19227
rect 12897 19227 12955 19233
rect 12897 19224 12909 19227
rect 12483 19196 12909 19224
rect 12483 19193 12495 19196
rect 12437 19187 12495 19193
rect 12897 19193 12909 19196
rect 12943 19193 12955 19227
rect 13906 19224 13912 19236
rect 12897 19187 12955 19193
rect 13096 19196 13912 19224
rect 9324 19128 10272 19156
rect 9033 19119 9091 19125
rect 10318 19116 10324 19168
rect 10376 19156 10382 19168
rect 10962 19156 10968 19168
rect 10376 19128 10968 19156
rect 10376 19116 10382 19128
rect 10962 19116 10968 19128
rect 11020 19156 11026 19168
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11020 19128 11253 19156
rect 11020 19116 11026 19128
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 11977 19159 12035 19165
rect 11977 19125 11989 19159
rect 12023 19156 12035 19159
rect 13096 19156 13124 19196
rect 13906 19184 13912 19196
rect 13964 19184 13970 19236
rect 14921 19227 14979 19233
rect 14921 19193 14933 19227
rect 14967 19224 14979 19227
rect 15654 19224 15660 19236
rect 14967 19196 15660 19224
rect 14967 19193 14979 19196
rect 14921 19187 14979 19193
rect 15654 19184 15660 19196
rect 15712 19184 15718 19236
rect 15841 19227 15899 19233
rect 15841 19193 15853 19227
rect 15887 19224 15899 19227
rect 16574 19224 16580 19236
rect 15887 19196 16580 19224
rect 15887 19193 15899 19196
rect 15841 19187 15899 19193
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 17402 19184 17408 19236
rect 17460 19224 17466 19236
rect 17497 19227 17555 19233
rect 17497 19224 17509 19227
rect 17460 19196 17509 19224
rect 17460 19184 17466 19196
rect 17497 19193 17509 19196
rect 17543 19193 17555 19227
rect 17497 19187 17555 19193
rect 18874 19184 18880 19236
rect 18932 19224 18938 19236
rect 18932 19196 19564 19224
rect 18932 19184 18938 19196
rect 12023 19128 13124 19156
rect 12023 19125 12035 19128
rect 11977 19119 12035 19125
rect 13446 19116 13452 19168
rect 13504 19156 13510 19168
rect 14277 19159 14335 19165
rect 14277 19156 14289 19159
rect 13504 19128 14289 19156
rect 13504 19116 13510 19128
rect 14277 19125 14289 19128
rect 14323 19125 14335 19159
rect 14277 19119 14335 19125
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 16485 19159 16543 19165
rect 16485 19156 16497 19159
rect 15344 19128 16497 19156
rect 15344 19116 15350 19128
rect 16485 19125 16497 19128
rect 16531 19125 16543 19159
rect 16485 19119 16543 19125
rect 17586 19116 17592 19168
rect 17644 19156 17650 19168
rect 19536 19165 19564 19196
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 17644 19128 18981 19156
rect 17644 19116 17650 19128
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 18969 19119 19027 19125
rect 19521 19159 19579 19165
rect 19521 19125 19533 19159
rect 19567 19125 19579 19159
rect 19521 19119 19579 19125
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 4065 18955 4123 18961
rect 4065 18952 4077 18955
rect 3804 18924 4077 18952
rect 2225 18887 2283 18893
rect 2225 18853 2237 18887
rect 2271 18884 2283 18887
rect 2314 18884 2320 18896
rect 2271 18856 2320 18884
rect 2271 18853 2283 18856
rect 2225 18847 2283 18853
rect 2314 18844 2320 18856
rect 2372 18844 2378 18896
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1486 18816 1492 18828
rect 1443 18788 1492 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1486 18776 1492 18788
rect 1544 18776 1550 18828
rect 1946 18816 1952 18828
rect 1907 18788 1952 18816
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 3234 18776 3240 18828
rect 3292 18816 3298 18828
rect 3329 18819 3387 18825
rect 3329 18816 3341 18819
rect 3292 18788 3341 18816
rect 3292 18776 3298 18788
rect 3329 18785 3341 18788
rect 3375 18785 3387 18819
rect 3329 18779 3387 18785
rect 3421 18819 3479 18825
rect 3421 18785 3433 18819
rect 3467 18816 3479 18819
rect 3804 18816 3832 18924
rect 4065 18921 4077 18924
rect 4111 18921 4123 18955
rect 4065 18915 4123 18921
rect 4525 18955 4583 18961
rect 4525 18921 4537 18955
rect 4571 18952 4583 18955
rect 5166 18952 5172 18964
rect 4571 18924 5172 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 6822 18952 6828 18964
rect 6783 18924 6828 18952
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 6914 18912 6920 18964
rect 6972 18952 6978 18964
rect 11054 18952 11060 18964
rect 6972 18924 11060 18952
rect 6972 18912 6978 18924
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 11698 18912 11704 18964
rect 11756 18952 11762 18964
rect 12434 18952 12440 18964
rect 11756 18924 12440 18952
rect 11756 18912 11762 18924
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12989 18955 13047 18961
rect 12989 18921 13001 18955
rect 13035 18952 13047 18955
rect 13078 18952 13084 18964
rect 13035 18924 13084 18952
rect 13035 18921 13047 18924
rect 12989 18915 13047 18921
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 15841 18955 15899 18961
rect 15841 18952 15853 18955
rect 14516 18924 15853 18952
rect 14516 18912 14522 18924
rect 15841 18921 15853 18924
rect 15887 18952 15899 18955
rect 16022 18952 16028 18964
rect 15887 18924 16028 18952
rect 15887 18921 15899 18924
rect 15841 18915 15899 18921
rect 16022 18912 16028 18924
rect 16080 18912 16086 18964
rect 18966 18952 18972 18964
rect 17788 18924 18972 18952
rect 5712 18887 5770 18893
rect 5712 18853 5724 18887
rect 5758 18884 5770 18887
rect 5902 18884 5908 18896
rect 5758 18856 5908 18884
rect 5758 18853 5770 18856
rect 5712 18847 5770 18853
rect 5902 18844 5908 18856
rect 5960 18844 5966 18896
rect 7098 18844 7104 18896
rect 7156 18884 7162 18896
rect 10042 18884 10048 18896
rect 7156 18856 10048 18884
rect 7156 18844 7162 18856
rect 10042 18844 10048 18856
rect 10100 18844 10106 18896
rect 12161 18887 12219 18893
rect 12161 18853 12173 18887
rect 12207 18884 12219 18887
rect 13262 18884 13268 18896
rect 12207 18856 13268 18884
rect 12207 18853 12219 18856
rect 12161 18847 12219 18853
rect 13262 18844 13268 18856
rect 13320 18844 13326 18896
rect 13446 18884 13452 18896
rect 13407 18856 13452 18884
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 14277 18887 14335 18893
rect 14277 18853 14289 18887
rect 14323 18884 14335 18887
rect 16298 18884 16304 18896
rect 14323 18856 16304 18884
rect 14323 18853 14335 18856
rect 14277 18847 14335 18853
rect 16298 18844 16304 18856
rect 16356 18844 16362 18896
rect 16666 18884 16672 18896
rect 16627 18856 16672 18884
rect 16666 18844 16672 18856
rect 16724 18844 16730 18896
rect 17788 18893 17816 18924
rect 18966 18912 18972 18924
rect 19024 18912 19030 18964
rect 17773 18887 17831 18893
rect 17773 18853 17785 18887
rect 17819 18853 17831 18887
rect 17773 18847 17831 18853
rect 18509 18887 18567 18893
rect 18509 18853 18521 18887
rect 18555 18884 18567 18887
rect 18598 18884 18604 18896
rect 18555 18856 18604 18884
rect 18555 18853 18567 18856
rect 18509 18847 18567 18853
rect 18598 18844 18604 18856
rect 18656 18844 18662 18896
rect 3467 18788 3832 18816
rect 4433 18819 4491 18825
rect 3467 18785 3479 18788
rect 3421 18779 3479 18785
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 7193 18819 7251 18825
rect 4479 18788 7144 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 3568 18720 3613 18748
rect 3568 18708 3574 18720
rect 4154 18708 4160 18760
rect 4212 18748 4218 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 4212 18720 4629 18748
rect 4212 18708 4218 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 5040 18720 5457 18748
rect 5040 18708 5046 18720
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 7116 18748 7144 18788
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7239 18788 8033 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8665 18819 8723 18825
rect 8665 18785 8677 18819
rect 8711 18816 8723 18819
rect 9766 18816 9772 18828
rect 8711 18788 9772 18816
rect 8711 18785 8723 18788
rect 8665 18779 8723 18785
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 10318 18825 10324 18828
rect 10312 18779 10324 18825
rect 10376 18816 10382 18828
rect 11885 18819 11943 18825
rect 10376 18788 10412 18816
rect 10318 18776 10324 18779
rect 10376 18776 10382 18788
rect 11885 18785 11897 18819
rect 11931 18816 11943 18819
rect 12434 18816 12440 18828
rect 11931 18788 12440 18816
rect 11931 18785 11943 18788
rect 11885 18779 11943 18785
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 13357 18819 13415 18825
rect 13357 18816 13369 18819
rect 12952 18788 13369 18816
rect 12952 18776 12958 18788
rect 13357 18785 13369 18788
rect 13403 18785 13415 18819
rect 13357 18779 13415 18785
rect 14001 18819 14059 18825
rect 14001 18785 14013 18819
rect 14047 18816 14059 18819
rect 14090 18816 14096 18828
rect 14047 18788 14096 18816
rect 14047 18785 14059 18788
rect 14001 18779 14059 18785
rect 14090 18776 14096 18788
rect 14148 18776 14154 18828
rect 15746 18816 15752 18828
rect 15707 18788 15752 18816
rect 15746 18776 15752 18788
rect 15804 18776 15810 18828
rect 16393 18819 16451 18825
rect 16393 18785 16405 18819
rect 16439 18816 16451 18819
rect 16574 18816 16580 18828
rect 16439 18788 16580 18816
rect 16439 18785 16451 18788
rect 16393 18779 16451 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 16816 18788 17509 18816
rect 16816 18776 16822 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17497 18779 17555 18785
rect 18233 18819 18291 18825
rect 18233 18785 18245 18819
rect 18279 18816 18291 18819
rect 18279 18788 18644 18816
rect 18279 18785 18291 18788
rect 18233 18779 18291 18785
rect 18616 18760 18644 18788
rect 7742 18748 7748 18760
rect 7116 18720 7748 18748
rect 5445 18711 5503 18717
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 8110 18748 8116 18760
rect 8071 18720 8116 18748
rect 8110 18708 8116 18720
rect 8168 18708 8174 18760
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8260 18720 8305 18748
rect 8260 18708 8266 18720
rect 8478 18708 8484 18760
rect 8536 18748 8542 18760
rect 8849 18751 8907 18757
rect 8849 18748 8861 18751
rect 8536 18720 8861 18748
rect 8536 18708 8542 18720
rect 8849 18717 8861 18720
rect 8895 18717 8907 18751
rect 8849 18711 8907 18717
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10045 18751 10103 18757
rect 10045 18748 10057 18751
rect 10008 18720 10057 18748
rect 10008 18708 10014 18720
rect 10045 18717 10057 18720
rect 10091 18717 10103 18751
rect 10045 18711 10103 18717
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18748 13691 18751
rect 13722 18748 13728 18760
rect 13679 18720 13728 18748
rect 13679 18717 13691 18720
rect 13633 18711 13691 18717
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 15930 18708 15936 18760
rect 15988 18748 15994 18760
rect 15988 18720 16033 18748
rect 15988 18708 15994 18720
rect 18598 18708 18604 18760
rect 18656 18708 18662 18760
rect 566 18640 572 18692
rect 624 18680 630 18692
rect 9674 18680 9680 18692
rect 624 18652 4108 18680
rect 624 18640 630 18652
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 2961 18615 3019 18621
rect 2961 18612 2973 18615
rect 2188 18584 2973 18612
rect 2188 18572 2194 18584
rect 2961 18581 2973 18584
rect 3007 18581 3019 18615
rect 4080 18612 4108 18652
rect 6380 18652 9680 18680
rect 6380 18612 6408 18652
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 12802 18640 12808 18692
rect 12860 18680 12866 18692
rect 20346 18680 20352 18692
rect 12860 18652 20352 18680
rect 12860 18640 12866 18652
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 4080 18584 6408 18612
rect 2961 18575 3019 18581
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7653 18615 7711 18621
rect 7653 18612 7665 18615
rect 7156 18584 7665 18612
rect 7156 18572 7162 18584
rect 7653 18581 7665 18584
rect 7699 18581 7711 18615
rect 7653 18575 7711 18581
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 8812 18584 11437 18612
rect 8812 18572 8818 18584
rect 11425 18581 11437 18584
rect 11471 18581 11483 18615
rect 11425 18575 11483 18581
rect 14642 18572 14648 18624
rect 14700 18612 14706 18624
rect 15381 18615 15439 18621
rect 15381 18612 15393 18615
rect 14700 18584 15393 18612
rect 14700 18572 14706 18584
rect 15381 18581 15393 18584
rect 15427 18581 15439 18615
rect 15381 18575 15439 18581
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 5261 18411 5319 18417
rect 5261 18408 5273 18411
rect 2004 18380 5273 18408
rect 2004 18368 2010 18380
rect 5261 18377 5273 18380
rect 5307 18377 5319 18411
rect 5261 18371 5319 18377
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 8168 18380 8217 18408
rect 8168 18368 8174 18380
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 8205 18371 8263 18377
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 11241 18411 11299 18417
rect 11241 18408 11253 18411
rect 10192 18380 11253 18408
rect 10192 18368 10198 18380
rect 11241 18377 11253 18380
rect 11287 18377 11299 18411
rect 11241 18371 11299 18377
rect 13446 18368 13452 18420
rect 13504 18408 13510 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13504 18380 14289 18408
rect 13504 18368 13510 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 14277 18371 14335 18377
rect 15028 18380 16681 18408
rect 1596 18244 3096 18272
rect 1596 18213 1624 18244
rect 1581 18207 1639 18213
rect 1581 18173 1593 18207
rect 1627 18173 1639 18207
rect 2130 18204 2136 18216
rect 2091 18176 2136 18204
rect 1581 18167 1639 18173
rect 2130 18164 2136 18176
rect 2188 18164 2194 18216
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18173 3019 18207
rect 3068 18204 3096 18244
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 5718 18272 5724 18284
rect 4120 18244 5724 18272
rect 4120 18232 4126 18244
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 5902 18272 5908 18284
rect 5863 18244 5908 18272
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 6003 18244 7297 18272
rect 6003 18204 6031 18244
rect 7285 18241 7297 18244
rect 7331 18241 7343 18275
rect 8754 18272 8760 18284
rect 8715 18244 8760 18272
rect 7285 18235 7343 18241
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 12437 18275 12495 18281
rect 8996 18244 9996 18272
rect 8996 18232 9002 18244
rect 7098 18204 7104 18216
rect 3068 18176 6031 18204
rect 7059 18176 7104 18204
rect 2961 18167 3019 18173
rect 1670 18096 1676 18148
rect 1728 18136 1734 18148
rect 2409 18139 2467 18145
rect 2409 18136 2421 18139
rect 1728 18108 2421 18136
rect 1728 18096 1734 18108
rect 2409 18105 2421 18108
rect 2455 18105 2467 18139
rect 2409 18099 2467 18105
rect 2976 18080 3004 18167
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 8665 18207 8723 18213
rect 7800 18176 8616 18204
rect 7800 18164 7806 18176
rect 3228 18139 3286 18145
rect 3228 18105 3240 18139
rect 3274 18136 3286 18139
rect 4154 18136 4160 18148
rect 3274 18108 4160 18136
rect 3274 18105 3286 18108
rect 3228 18099 3286 18105
rect 4154 18096 4160 18108
rect 4212 18096 4218 18148
rect 8588 18145 8616 18176
rect 8665 18173 8677 18207
rect 8711 18204 8723 18207
rect 8846 18204 8852 18216
rect 8711 18176 8852 18204
rect 8711 18173 8723 18176
rect 8665 18167 8723 18173
rect 8846 18164 8852 18176
rect 8904 18164 8910 18216
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9824 18176 9873 18204
rect 9824 18164 9830 18176
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 9968 18204 9996 18244
rect 12437 18241 12449 18275
rect 12483 18272 12495 18275
rect 12483 18244 12572 18272
rect 12483 18241 12495 18244
rect 12437 18235 12495 18241
rect 11882 18204 11888 18216
rect 9968 18176 11888 18204
rect 9861 18167 9919 18173
rect 5629 18139 5687 18145
rect 5629 18105 5641 18139
rect 5675 18136 5687 18139
rect 6273 18139 6331 18145
rect 6273 18136 6285 18139
rect 5675 18108 6285 18136
rect 5675 18105 5687 18108
rect 5629 18099 5687 18105
rect 6273 18105 6285 18108
rect 6319 18105 6331 18139
rect 8573 18139 8631 18145
rect 6273 18099 6331 18105
rect 7668 18108 8524 18136
rect 1762 18068 1768 18080
rect 1723 18040 1768 18068
rect 1762 18028 1768 18040
rect 1820 18028 1826 18080
rect 2958 18068 2964 18080
rect 2871 18040 2964 18068
rect 2958 18028 2964 18040
rect 3016 18068 3022 18080
rect 3418 18068 3424 18080
rect 3016 18040 3424 18068
rect 3016 18028 3022 18040
rect 3418 18028 3424 18040
rect 3476 18028 3482 18080
rect 3510 18028 3516 18080
rect 3568 18068 3574 18080
rect 4062 18068 4068 18080
rect 3568 18040 4068 18068
rect 3568 18028 3574 18040
rect 4062 18028 4068 18040
rect 4120 18068 4126 18080
rect 4341 18071 4399 18077
rect 4341 18068 4353 18071
rect 4120 18040 4353 18068
rect 4120 18028 4126 18040
rect 4341 18037 4353 18040
rect 4387 18037 4399 18071
rect 5718 18068 5724 18080
rect 5679 18040 5724 18068
rect 4341 18031 4399 18037
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 7668 18068 7696 18108
rect 5868 18040 7696 18068
rect 5868 18028 5874 18040
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 8386 18068 8392 18080
rect 7800 18040 8392 18068
rect 7800 18028 7806 18040
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 8496 18068 8524 18108
rect 8573 18105 8585 18139
rect 8619 18136 8631 18139
rect 9398 18136 9404 18148
rect 8619 18108 9404 18136
rect 8619 18105 8631 18108
rect 8573 18099 8631 18105
rect 9398 18096 9404 18108
rect 9456 18096 9462 18148
rect 9876 18136 9904 18167
rect 11882 18164 11888 18176
rect 11940 18164 11946 18216
rect 9950 18136 9956 18148
rect 9876 18108 9956 18136
rect 9950 18096 9956 18108
rect 10008 18096 10014 18148
rect 10128 18139 10186 18145
rect 10128 18105 10140 18139
rect 10174 18136 10186 18139
rect 10226 18136 10232 18148
rect 10174 18108 10232 18136
rect 10174 18105 10186 18108
rect 10128 18099 10186 18105
rect 10226 18096 10232 18108
rect 10284 18096 10290 18148
rect 10410 18096 10416 18148
rect 10468 18136 10474 18148
rect 12158 18136 12164 18148
rect 10468 18108 12164 18136
rect 10468 18096 10474 18108
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 12544 18136 12572 18244
rect 13446 18232 13452 18284
rect 13504 18272 13510 18284
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 13504 18244 14933 18272
rect 13504 18232 13510 18244
rect 14921 18241 14933 18244
rect 14967 18272 14979 18275
rect 15028 18272 15056 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 16669 18371 16727 18377
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 17862 18408 17868 18420
rect 17635 18380 17868 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 14967 18244 15056 18272
rect 18325 18275 18383 18281
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 18506 18272 18512 18284
rect 18371 18244 18512 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 12704 18207 12762 18213
rect 12704 18173 12716 18207
rect 12750 18204 12762 18207
rect 13464 18204 13492 18232
rect 14642 18204 14648 18216
rect 12750 18176 13492 18204
rect 14603 18176 14648 18204
rect 12750 18173 12762 18176
rect 12704 18167 12762 18173
rect 14642 18164 14648 18176
rect 14700 18164 14706 18216
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18204 15347 18207
rect 17402 18204 17408 18216
rect 15335 18176 15516 18204
rect 17363 18176 17408 18204
rect 15335 18173 15347 18176
rect 15289 18167 15347 18173
rect 13078 18136 13084 18148
rect 12544 18108 13084 18136
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 15488 18080 15516 18176
rect 17402 18164 17408 18176
rect 17460 18164 17466 18216
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18966 18204 18972 18216
rect 18095 18176 18972 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18966 18164 18972 18176
rect 19024 18164 19030 18216
rect 15556 18139 15614 18145
rect 15556 18105 15568 18139
rect 15602 18136 15614 18139
rect 15930 18136 15936 18148
rect 15602 18108 15936 18136
rect 15602 18105 15614 18108
rect 15556 18099 15614 18105
rect 15930 18096 15936 18108
rect 15988 18096 15994 18148
rect 19702 18096 19708 18148
rect 19760 18136 19766 18148
rect 22554 18136 22560 18148
rect 19760 18108 22560 18136
rect 19760 18096 19766 18108
rect 22554 18096 22560 18108
rect 22612 18096 22618 18148
rect 8938 18068 8944 18080
rect 8496 18040 8944 18068
rect 8938 18028 8944 18040
rect 8996 18028 9002 18080
rect 9030 18028 9036 18080
rect 9088 18068 9094 18080
rect 10686 18068 10692 18080
rect 9088 18040 10692 18068
rect 9088 18028 9094 18040
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 10962 18028 10968 18080
rect 11020 18068 11026 18080
rect 11606 18068 11612 18080
rect 11020 18040 11612 18068
rect 11020 18028 11026 18040
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 13722 18028 13728 18080
rect 13780 18068 13786 18080
rect 13817 18071 13875 18077
rect 13817 18068 13829 18071
rect 13780 18040 13829 18068
rect 13780 18028 13786 18040
rect 13817 18037 13829 18040
rect 13863 18037 13875 18071
rect 13817 18031 13875 18037
rect 14737 18071 14795 18077
rect 14737 18037 14749 18071
rect 14783 18068 14795 18071
rect 15286 18068 15292 18080
rect 14783 18040 15292 18068
rect 14783 18037 14795 18040
rect 14737 18031 14795 18037
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 15470 18028 15476 18080
rect 15528 18028 15534 18080
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 20254 18068 20260 18080
rect 19668 18040 20260 18068
rect 19668 18028 19674 18040
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 21634 18068 21640 18080
rect 20956 18040 21640 18068
rect 20956 18028 20962 18040
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 3234 17824 3240 17876
rect 3292 17864 3298 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 3292 17836 3341 17864
rect 3292 17824 3298 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 3329 17827 3387 17833
rect 5902 17824 5908 17876
rect 5960 17864 5966 17876
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 5960 17836 6745 17864
rect 5960 17824 5966 17836
rect 6733 17833 6745 17836
rect 6779 17833 6791 17867
rect 6733 17827 6791 17833
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 9916 17836 10149 17864
rect 9916 17824 9922 17836
rect 10137 17833 10149 17836
rect 10183 17833 10195 17867
rect 10137 17827 10195 17833
rect 12069 17867 12127 17873
rect 12069 17833 12081 17867
rect 12115 17864 12127 17867
rect 12894 17864 12900 17876
rect 12115 17836 12900 17864
rect 12115 17833 12127 17836
rect 12069 17827 12127 17833
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15654 17864 15660 17876
rect 15615 17836 15660 17864
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 17405 17867 17463 17873
rect 17405 17833 17417 17867
rect 17451 17864 17463 17867
rect 18598 17864 18604 17876
rect 17451 17836 18604 17864
rect 17451 17833 17463 17836
rect 17405 17827 17463 17833
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 9674 17756 9680 17808
rect 9732 17796 9738 17808
rect 12710 17796 12716 17808
rect 9732 17768 12716 17796
rect 9732 17756 9738 17768
rect 12710 17756 12716 17768
rect 12768 17796 12774 17808
rect 13348 17799 13406 17805
rect 12768 17768 13308 17796
rect 12768 17756 12774 17768
rect 2682 17737 2688 17740
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1397 17691 1455 17697
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2673 17731 2688 17737
rect 1995 17700 2360 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 1412 17592 1440 17691
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 2133 17663 2191 17669
rect 2133 17660 2145 17663
rect 1636 17632 2145 17660
rect 1636 17620 1642 17632
rect 2133 17629 2145 17632
rect 2179 17629 2191 17663
rect 2332 17660 2360 17700
rect 2673 17697 2685 17731
rect 2673 17691 2688 17697
rect 2682 17688 2688 17691
rect 2740 17688 2746 17740
rect 4982 17688 4988 17740
rect 5040 17728 5046 17740
rect 5353 17731 5411 17737
rect 5353 17728 5365 17731
rect 5040 17700 5365 17728
rect 5040 17688 5046 17700
rect 5353 17697 5365 17700
rect 5399 17697 5411 17731
rect 5353 17691 5411 17697
rect 5620 17731 5678 17737
rect 5620 17697 5632 17731
rect 5666 17728 5678 17731
rect 6178 17728 6184 17740
rect 5666 17700 6184 17728
rect 5666 17697 5678 17700
rect 5620 17691 5678 17697
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 7006 17728 7012 17740
rect 6967 17700 7012 17728
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 7116 17700 10057 17728
rect 5166 17660 5172 17672
rect 2332 17632 5172 17660
rect 2133 17623 2191 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6362 17620 6368 17672
rect 6420 17660 6426 17672
rect 7116 17660 7144 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 12437 17731 12495 17737
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 13170 17728 13176 17740
rect 12483 17700 13176 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 13280 17728 13308 17768
rect 13348 17765 13360 17799
rect 13394 17796 13406 17799
rect 13722 17796 13728 17808
rect 13394 17768 13728 17796
rect 13394 17765 13406 17768
rect 13348 17759 13406 17765
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 15749 17731 15807 17737
rect 15749 17728 15761 17731
rect 13280 17700 15761 17728
rect 15749 17697 15761 17700
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 18417 17731 18475 17737
rect 18417 17728 18429 17731
rect 17819 17700 18429 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 18417 17697 18429 17700
rect 18463 17697 18475 17731
rect 18417 17691 18475 17697
rect 6420 17632 7144 17660
rect 7193 17663 7251 17669
rect 6420 17620 6426 17632
rect 7193 17629 7205 17663
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10410 17660 10416 17672
rect 10367 17632 10416 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 7208 17592 7236 17623
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 12526 17660 12532 17672
rect 12487 17632 12532 17660
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 13078 17660 13084 17672
rect 12759 17632 12940 17660
rect 13039 17632 13084 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 1412 17564 5028 17592
rect 2866 17524 2872 17536
rect 2827 17496 2872 17524
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 5000 17524 5028 17564
rect 6288 17564 7236 17592
rect 6288 17524 6316 17564
rect 5000 17496 6316 17524
rect 9677 17527 9735 17533
rect 9677 17493 9689 17527
rect 9723 17524 9735 17527
rect 10134 17524 10140 17536
rect 9723 17496 10140 17524
rect 9723 17493 9735 17496
rect 9677 17487 9735 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 12912 17524 12940 17632
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 15930 17660 15936 17672
rect 15891 17632 15936 17660
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 17865 17663 17923 17669
rect 17865 17660 17877 17663
rect 17000 17632 17877 17660
rect 17000 17620 17006 17632
rect 17865 17629 17877 17632
rect 17911 17629 17923 17663
rect 17865 17623 17923 17629
rect 18049 17663 18107 17669
rect 18049 17629 18061 17663
rect 18095 17660 18107 17663
rect 19426 17660 19432 17672
rect 18095 17632 19432 17660
rect 18095 17629 18107 17632
rect 18049 17623 18107 17629
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 13446 17524 13452 17536
rect 12912 17496 13452 17524
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 14461 17527 14519 17533
rect 14461 17493 14473 17527
rect 14507 17524 14519 17527
rect 14550 17524 14556 17536
rect 14507 17496 14556 17524
rect 14507 17493 14519 17496
rect 14461 17487 14519 17493
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 3142 17320 3148 17332
rect 1627 17292 3148 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 3234 17280 3240 17332
rect 3292 17320 3298 17332
rect 5629 17323 5687 17329
rect 3292 17292 3924 17320
rect 3292 17280 3298 17292
rect 3896 17252 3924 17292
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 5718 17320 5724 17332
rect 5675 17292 5724 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 12437 17323 12495 17329
rect 5828 17292 11008 17320
rect 5828 17252 5856 17292
rect 3896 17224 5856 17252
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 2133 17187 2191 17193
rect 2133 17184 2145 17187
rect 1544 17156 2145 17184
rect 1544 17144 1550 17156
rect 2133 17153 2145 17156
rect 2179 17153 2191 17187
rect 2958 17184 2964 17196
rect 2919 17156 2964 17184
rect 2133 17147 2191 17153
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 6086 17184 6092 17196
rect 6047 17156 6092 17184
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6178 17144 6184 17196
rect 6236 17184 6242 17196
rect 6236 17156 6281 17184
rect 6236 17144 6242 17156
rect 1394 17116 1400 17128
rect 1355 17088 1400 17116
rect 1394 17076 1400 17088
rect 1452 17076 1458 17128
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17085 2007 17119
rect 1949 17079 2007 17085
rect 3228 17119 3286 17125
rect 3228 17085 3240 17119
rect 3274 17116 3286 17119
rect 4062 17116 4068 17128
rect 3274 17088 4068 17116
rect 3274 17085 3286 17088
rect 3228 17079 3286 17085
rect 1964 16980 1992 17079
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17116 6055 17119
rect 6362 17116 6368 17128
rect 6043 17088 6368 17116
rect 6043 17085 6055 17088
rect 5997 17079 6055 17085
rect 6362 17076 6368 17088
rect 6420 17076 6426 17128
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17085 7527 17119
rect 7469 17079 7527 17085
rect 7736 17119 7794 17125
rect 7736 17085 7748 17119
rect 7782 17116 7794 17119
rect 8202 17116 8208 17128
rect 7782 17088 8208 17116
rect 7782 17085 7794 17088
rect 7736 17079 7794 17085
rect 7098 17008 7104 17060
rect 7156 17048 7162 17060
rect 7484 17048 7512 17079
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 8754 17076 8760 17128
rect 8812 17116 8818 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 8812 17088 9689 17116
rect 8812 17076 8818 17088
rect 9677 17085 9689 17088
rect 9723 17116 9735 17119
rect 9766 17116 9772 17128
rect 9723 17088 9772 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 10980 17116 11008 17292
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12618 17320 12624 17332
rect 12483 17292 12624 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 16942 17320 16948 17332
rect 16903 17292 16948 17320
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 11054 17212 11060 17264
rect 11112 17252 11118 17264
rect 14458 17252 14464 17264
rect 11112 17224 14464 17252
rect 11112 17212 11118 17224
rect 14458 17212 14464 17224
rect 14516 17212 14522 17264
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12308 17156 13001 17184
rect 12308 17144 12314 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 13228 17156 13461 17184
rect 13228 17144 13234 17156
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 16022 17144 16028 17196
rect 16080 17184 16086 17196
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 16080 17156 17417 17184
rect 16080 17144 16086 17156
rect 17405 17153 17417 17156
rect 17451 17153 17463 17187
rect 17586 17184 17592 17196
rect 17547 17156 17592 17184
rect 17405 17147 17463 17153
rect 17586 17144 17592 17156
rect 17644 17184 17650 17196
rect 17644 17156 18184 17184
rect 17644 17144 17650 17156
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 10980 17088 17325 17116
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17920 17088 18061 17116
rect 17920 17076 17926 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18156 17116 18184 17156
rect 18305 17119 18363 17125
rect 18305 17116 18317 17119
rect 18156 17088 18317 17116
rect 18049 17079 18107 17085
rect 18305 17085 18317 17088
rect 18351 17085 18363 17119
rect 18305 17079 18363 17085
rect 7650 17048 7656 17060
rect 7156 17020 7656 17048
rect 7156 17008 7162 17020
rect 7650 17008 7656 17020
rect 7708 17048 7714 17060
rect 8772 17048 8800 17076
rect 7708 17020 8800 17048
rect 9944 17051 10002 17057
rect 7708 17008 7714 17020
rect 9944 17017 9956 17051
rect 9990 17048 10002 17051
rect 10410 17048 10416 17060
rect 9990 17020 10416 17048
rect 9990 17017 10002 17020
rect 9944 17011 10002 17017
rect 10410 17008 10416 17020
rect 10468 17008 10474 17060
rect 4062 16980 4068 16992
rect 1964 16952 4068 16980
rect 4062 16940 4068 16952
rect 4120 16940 4126 16992
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4341 16983 4399 16989
rect 4341 16980 4353 16983
rect 4212 16952 4353 16980
rect 4212 16940 4218 16952
rect 4341 16949 4353 16952
rect 4387 16949 4399 16983
rect 4341 16943 4399 16949
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 8849 16983 8907 16989
rect 8849 16980 8861 16983
rect 8260 16952 8861 16980
rect 8260 16940 8266 16952
rect 8849 16949 8861 16952
rect 8895 16949 8907 16983
rect 8849 16943 8907 16949
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16980 9275 16983
rect 10042 16980 10048 16992
rect 9263 16952 10048 16980
rect 9263 16949 9275 16952
rect 9217 16943 9275 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 10284 16952 11069 16980
rect 10284 16940 10290 16952
rect 11057 16949 11069 16952
rect 11103 16949 11115 16983
rect 11057 16943 11115 16949
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12584 16952 12817 16980
rect 12584 16940 12590 16952
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 12805 16943 12863 16949
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 19426 16980 19432 16992
rect 12952 16952 12997 16980
rect 19387 16952 19432 16980
rect 12952 16940 12958 16952
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2056 16748 2881 16776
rect 1489 16643 1547 16649
rect 1489 16609 1501 16643
rect 1535 16640 1547 16643
rect 1578 16640 1584 16652
rect 1535 16612 1584 16640
rect 1535 16609 1547 16612
rect 1489 16603 1547 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 2056 16649 2084 16748
rect 2869 16745 2881 16748
rect 2915 16745 2927 16779
rect 2869 16739 2927 16745
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 4246 16776 4252 16788
rect 3936 16748 4252 16776
rect 3936 16736 3942 16748
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 6236 16748 6377 16776
rect 6236 16736 6242 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 6365 16739 6423 16745
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16745 9735 16779
rect 10042 16776 10048 16788
rect 10003 16748 10048 16776
rect 9677 16739 9735 16745
rect 5166 16668 5172 16720
rect 5224 16708 5230 16720
rect 9692 16708 9720 16739
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 12526 16776 12532 16788
rect 10192 16748 10237 16776
rect 12487 16748 12532 16776
rect 10192 16736 10198 16748
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 12952 16748 13553 16776
rect 12952 16736 12958 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 13541 16739 13599 16745
rect 15930 16736 15936 16788
rect 15988 16776 15994 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 15988 16748 16681 16776
rect 15988 16736 15994 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 5224 16680 9720 16708
rect 11140 16711 11198 16717
rect 5224 16668 5230 16680
rect 11140 16677 11152 16711
rect 11186 16708 11198 16711
rect 18132 16711 18190 16717
rect 11186 16680 13216 16708
rect 11186 16677 11198 16680
rect 11140 16671 11198 16677
rect 2051 16643 2109 16649
rect 2051 16609 2063 16643
rect 2097 16609 2109 16643
rect 3234 16640 3240 16652
rect 3195 16612 3240 16640
rect 2051 16603 2109 16609
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16640 3387 16643
rect 4246 16640 4252 16652
rect 3375 16612 4252 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 5252 16643 5310 16649
rect 5252 16609 5264 16643
rect 5298 16640 5310 16643
rect 5810 16640 5816 16652
rect 5298 16612 5816 16640
rect 5298 16609 5310 16612
rect 5252 16603 5310 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 7190 16640 7196 16652
rect 6687 16612 7196 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7368 16643 7426 16649
rect 7368 16609 7380 16643
rect 7414 16640 7426 16643
rect 8202 16640 8208 16652
rect 7414 16612 8208 16640
rect 7414 16609 7426 16612
rect 7368 16603 7426 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8312 16612 8953 16640
rect 1394 16532 1400 16584
rect 1452 16572 1458 16584
rect 2225 16575 2283 16581
rect 2225 16572 2237 16575
rect 1452 16544 2237 16572
rect 1452 16532 1458 16544
rect 2225 16541 2237 16544
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 3513 16575 3571 16581
rect 3513 16541 3525 16575
rect 3559 16572 3571 16575
rect 3970 16572 3976 16584
rect 3559 16544 3976 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4982 16572 4988 16584
rect 4943 16544 4988 16572
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 7098 16572 7104 16584
rect 7059 16544 7104 16572
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8312 16572 8340 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 12894 16640 12900 16652
rect 12855 16612 12900 16640
rect 8941 16603 8999 16609
rect 12894 16600 12900 16612
rect 12952 16600 12958 16652
rect 10226 16572 10232 16584
rect 8168 16544 8340 16572
rect 10187 16544 10232 16572
rect 8168 16532 8174 16544
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 10870 16572 10876 16584
rect 10831 16544 10876 16572
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 12986 16572 12992 16584
rect 12947 16544 12992 16572
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 13188 16581 13216 16680
rect 18132 16677 18144 16711
rect 18178 16708 18190 16711
rect 19426 16708 19432 16720
rect 18178 16680 19432 16708
rect 18178 16677 18190 16680
rect 18132 16671 18190 16677
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 13906 16640 13912 16652
rect 13867 16612 13912 16640
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15545 16643 15603 16649
rect 15545 16640 15557 16643
rect 15252 16612 15557 16640
rect 15252 16600 15258 16612
rect 15545 16609 15557 16612
rect 15591 16609 15603 16643
rect 15545 16603 15603 16609
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 17862 16640 17868 16652
rect 16356 16612 17868 16640
rect 16356 16600 16362 16612
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16541 13231 16575
rect 13998 16572 14004 16584
rect 13959 16544 14004 16572
rect 13173 16535 13231 16541
rect 13188 16504 13216 16535
rect 13998 16532 14004 16544
rect 14056 16532 14062 16584
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16572 14243 16575
rect 14734 16572 14740 16584
rect 14231 16544 14740 16572
rect 14231 16541 14243 16544
rect 14185 16535 14243 16541
rect 14200 16504 14228 16535
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 13188 16476 14228 16504
rect 8478 16436 8484 16448
rect 8439 16408 8484 16436
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 8754 16436 8760 16448
rect 8715 16408 8760 16436
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 12250 16436 12256 16448
rect 12211 16408 12256 16436
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 15304 16436 15332 16535
rect 15470 16436 15476 16448
rect 15304 16408 15476 16436
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 19242 16436 19248 16448
rect 19203 16408 19248 16436
rect 19242 16396 19248 16408
rect 19300 16396 19306 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2958 16232 2964 16244
rect 2608 16204 2964 16232
rect 2608 16105 2636 16204
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 4246 16232 4252 16244
rect 4207 16204 4252 16232
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 10410 16232 10416 16244
rect 10371 16204 10416 16232
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 12529 16235 12587 16241
rect 12529 16201 12541 16235
rect 12575 16232 12587 16235
rect 12621 16235 12679 16241
rect 12621 16232 12633 16235
rect 12575 16204 12633 16232
rect 12575 16201 12587 16204
rect 12529 16195 12587 16201
rect 12621 16201 12633 16204
rect 12667 16232 12679 16235
rect 13078 16232 13084 16244
rect 12667 16204 13084 16232
rect 12667 16201 12679 16204
rect 12621 16195 12679 16201
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13998 16192 14004 16244
rect 14056 16232 14062 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14056 16204 15025 16232
rect 14056 16192 14062 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 16025 16235 16083 16241
rect 16025 16232 16037 16235
rect 15528 16204 16037 16232
rect 15528 16192 15534 16204
rect 16025 16201 16037 16204
rect 16071 16201 16083 16235
rect 16025 16195 16083 16201
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 5261 16167 5319 16173
rect 5261 16164 5273 16167
rect 4120 16136 5273 16164
rect 4120 16124 4126 16136
rect 5261 16133 5273 16136
rect 5307 16133 5319 16167
rect 5261 16127 5319 16133
rect 10778 16124 10784 16176
rect 10836 16164 10842 16176
rect 12802 16164 12808 16176
rect 10836 16136 12808 16164
rect 10836 16124 10842 16136
rect 12802 16124 12808 16136
rect 12860 16124 12866 16176
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16065 2651 16099
rect 4706 16096 4712 16108
rect 4667 16068 4712 16096
rect 2593 16059 2651 16065
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16065 4859 16099
rect 5810 16096 5816 16108
rect 5771 16068 5816 16096
rect 4801 16059 4859 16065
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 2860 16031 2918 16037
rect 2860 15997 2872 16031
rect 2906 16028 2918 16031
rect 4154 16028 4160 16040
rect 2906 16000 4160 16028
rect 2906 15997 2918 16000
rect 2860 15991 2918 15997
rect 4154 15988 4160 16000
rect 4212 16028 4218 16040
rect 4816 16028 4844 16059
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7800 16068 7941 16096
rect 7800 16056 7806 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 8113 16099 8171 16105
rect 8113 16065 8125 16099
rect 8159 16096 8171 16099
rect 8202 16096 8208 16108
rect 8159 16068 8208 16096
rect 8159 16065 8171 16068
rect 8113 16059 8171 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 12894 16096 12900 16108
rect 12855 16068 12900 16096
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 13096 16096 13124 16192
rect 14734 16164 14740 16176
rect 14695 16136 14740 16164
rect 14734 16124 14740 16136
rect 14792 16124 14798 16176
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13096 16068 13369 16096
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 15565 16099 15623 16105
rect 15565 16096 15577 16099
rect 13357 16059 13415 16065
rect 14568 16068 15577 16096
rect 14568 16040 14596 16068
rect 15565 16065 15577 16068
rect 15611 16065 15623 16099
rect 16040 16096 16068 16195
rect 17586 16192 17592 16244
rect 17644 16232 17650 16244
rect 17681 16235 17739 16241
rect 17681 16232 17693 16235
rect 17644 16204 17693 16232
rect 17644 16192 17650 16204
rect 17681 16201 17693 16204
rect 17727 16201 17739 16235
rect 17681 16195 17739 16201
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 18012 16204 18061 16232
rect 18012 16192 18018 16204
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 16298 16096 16304 16108
rect 16040 16068 16304 16096
rect 15565 16059 15623 16065
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 18690 16096 18696 16108
rect 18651 16068 18696 16096
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 4212 16000 4844 16028
rect 4908 16000 7849 16028
rect 4212 15988 4218 16000
rect 4908 15904 4936 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 8754 16028 8760 16040
rect 8444 16000 8760 16028
rect 8444 15988 8450 16000
rect 8754 15988 8760 16000
rect 8812 16028 8818 16040
rect 9033 16031 9091 16037
rect 9033 16028 9045 16031
rect 8812 16000 9045 16028
rect 8812 15988 8818 16000
rect 9033 15997 9045 16000
rect 9079 15997 9091 16031
rect 9033 15991 9091 15997
rect 12805 16031 12863 16037
rect 12805 15997 12817 16031
rect 12851 15997 12863 16031
rect 12805 15991 12863 15997
rect 13624 16031 13682 16037
rect 13624 15997 13636 16031
rect 13670 16028 13682 16031
rect 14550 16028 14556 16040
rect 13670 16000 14556 16028
rect 13670 15997 13682 16000
rect 13624 15991 13682 15997
rect 5629 15963 5687 15969
rect 5629 15929 5641 15963
rect 5675 15960 5687 15963
rect 6273 15963 6331 15969
rect 6273 15960 6285 15963
rect 5675 15932 6285 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 6273 15929 6285 15932
rect 6319 15929 6331 15963
rect 6273 15923 6331 15929
rect 9300 15963 9358 15969
rect 9300 15929 9312 15963
rect 9346 15960 9358 15963
rect 9766 15960 9772 15972
rect 9346 15932 9772 15960
rect 9346 15929 9358 15932
rect 9300 15923 9358 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 11882 15920 11888 15972
rect 11940 15960 11946 15972
rect 12820 15960 12848 15991
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 16209 16031 16267 16037
rect 16209 15997 16221 16031
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 15286 15960 15292 15972
rect 11940 15932 12756 15960
rect 12820 15932 15292 15960
rect 11940 15920 11946 15932
rect 3970 15892 3976 15904
rect 3931 15864 3976 15892
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 4890 15892 4896 15904
rect 4663 15864 4896 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5718 15892 5724 15904
rect 5679 15864 5724 15892
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 7469 15895 7527 15901
rect 7469 15892 7481 15895
rect 7340 15864 7481 15892
rect 7340 15852 7346 15864
rect 7469 15861 7481 15864
rect 7515 15861 7527 15895
rect 7469 15855 7527 15861
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 12400 15864 12541 15892
rect 12400 15852 12406 15864
rect 12529 15861 12541 15864
rect 12575 15861 12587 15895
rect 12728 15892 12756 15932
rect 15286 15920 15292 15932
rect 15344 15960 15350 15972
rect 16224 15960 16252 15991
rect 15344 15932 16252 15960
rect 16568 15963 16626 15969
rect 15344 15920 15350 15932
rect 16568 15929 16580 15963
rect 16614 15960 16626 15963
rect 17126 15960 17132 15972
rect 16614 15932 17132 15960
rect 16614 15929 16626 15932
rect 16568 15923 16626 15929
rect 17126 15920 17132 15932
rect 17184 15920 17190 15972
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 18509 15963 18567 15969
rect 18509 15960 18521 15963
rect 18012 15932 18521 15960
rect 18012 15920 18018 15932
rect 18509 15929 18521 15932
rect 18555 15929 18567 15963
rect 18509 15923 18567 15929
rect 13998 15892 14004 15904
rect 12728 15864 14004 15892
rect 12529 15855 12587 15861
rect 13998 15852 14004 15864
rect 14056 15892 14062 15904
rect 15381 15895 15439 15901
rect 15381 15892 15393 15895
rect 14056 15864 15393 15892
rect 14056 15852 14062 15864
rect 15381 15861 15393 15864
rect 15427 15861 15439 15895
rect 15381 15855 15439 15861
rect 15473 15895 15531 15901
rect 15473 15861 15485 15895
rect 15519 15892 15531 15895
rect 15654 15892 15660 15904
rect 15519 15864 15660 15892
rect 15519 15861 15531 15864
rect 15473 15855 15531 15861
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 18414 15892 18420 15904
rect 18375 15864 18420 15892
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 2130 15688 2136 15700
rect 1627 15660 2136 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 3234 15688 3240 15700
rect 3195 15660 3240 15688
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 5810 15648 5816 15700
rect 5868 15688 5874 15700
rect 6181 15691 6239 15697
rect 6181 15688 6193 15691
rect 5868 15660 6193 15688
rect 5868 15648 5874 15660
rect 6181 15657 6193 15660
rect 6227 15657 6239 15691
rect 6181 15651 6239 15657
rect 6457 15691 6515 15697
rect 6457 15657 6469 15691
rect 6503 15657 6515 15691
rect 6457 15651 6515 15657
rect 6825 15691 6883 15697
rect 6825 15657 6837 15691
rect 6871 15688 6883 15691
rect 7006 15688 7012 15700
rect 6871 15660 7012 15688
rect 6871 15657 6883 15660
rect 6825 15651 6883 15657
rect 1762 15580 1768 15632
rect 1820 15620 1826 15632
rect 2225 15623 2283 15629
rect 2225 15620 2237 15623
rect 1820 15592 2237 15620
rect 1820 15580 1826 15592
rect 2225 15589 2237 15592
rect 2271 15589 2283 15623
rect 4982 15620 4988 15632
rect 2225 15583 2283 15589
rect 4816 15592 4988 15620
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 1959 15555 2017 15561
rect 1959 15521 1971 15555
rect 2005 15521 2017 15555
rect 1959 15515 2017 15521
rect 1964 15348 1992 15515
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4816 15493 4844 15592
rect 4982 15580 4988 15592
rect 5040 15620 5046 15632
rect 6472 15620 6500 15651
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15688 7895 15691
rect 8202 15688 8208 15700
rect 7883 15660 8208 15688
rect 7883 15657 7895 15660
rect 7837 15651 7895 15657
rect 7190 15620 7196 15632
rect 5040 15592 6500 15620
rect 7151 15592 7196 15620
rect 5040 15580 5046 15592
rect 7190 15580 7196 15592
rect 7248 15580 7254 15632
rect 5068 15555 5126 15561
rect 5068 15521 5080 15555
rect 5114 15552 5126 15555
rect 6178 15552 6184 15564
rect 5114 15524 6184 15552
rect 5114 15521 5126 15524
rect 5068 15515 5126 15521
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 7852 15552 7880 15651
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9079 15660 9689 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 10318 15688 10324 15700
rect 10183 15660 10324 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12986 15688 12992 15700
rect 12124 15660 12909 15688
rect 12947 15660 12992 15688
rect 12124 15648 12130 15660
rect 11232 15623 11290 15629
rect 11232 15589 11244 15623
rect 11278 15620 11290 15623
rect 12250 15620 12256 15632
rect 11278 15592 12256 15620
rect 11278 15589 11290 15592
rect 11232 15583 11290 15589
rect 12250 15580 12256 15592
rect 12308 15580 12314 15632
rect 12881 15620 12909 15660
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14001 15691 14059 15697
rect 14001 15688 14013 15691
rect 13964 15660 14013 15688
rect 13964 15648 13970 15660
rect 14001 15657 14013 15660
rect 14047 15657 14059 15691
rect 14458 15688 14464 15700
rect 14419 15660 14464 15688
rect 14001 15651 14059 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 15286 15648 15292 15700
rect 15344 15688 15350 15700
rect 15473 15691 15531 15697
rect 15473 15688 15485 15691
rect 15344 15660 15485 15688
rect 15344 15648 15350 15660
rect 15473 15657 15485 15660
rect 15519 15657 15531 15691
rect 17126 15688 17132 15700
rect 17087 15660 17132 15688
rect 15473 15651 15531 15657
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 17954 15688 17960 15700
rect 17915 15660 17960 15688
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 18969 15691 19027 15697
rect 18969 15688 18981 15691
rect 18472 15660 18981 15688
rect 18472 15648 18478 15660
rect 18969 15657 18981 15660
rect 19015 15657 19027 15691
rect 18969 15651 19027 15657
rect 14369 15623 14427 15629
rect 14369 15620 14381 15623
rect 12881 15592 14381 15620
rect 14369 15589 14381 15592
rect 14415 15620 14427 15623
rect 15102 15620 15108 15632
rect 14415 15592 15108 15620
rect 14415 15589 14427 15592
rect 14369 15583 14427 15589
rect 15102 15580 15108 15592
rect 15160 15620 15166 15632
rect 16016 15623 16074 15629
rect 15160 15592 15884 15620
rect 15160 15580 15166 15592
rect 6687 15524 7880 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 7926 15512 7932 15564
rect 7984 15552 7990 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7984 15524 8033 15552
rect 7984 15512 7990 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8941 15555 8999 15561
rect 8941 15521 8953 15555
rect 8987 15552 8999 15555
rect 9674 15552 9680 15564
rect 8987 15524 9680 15552
rect 8987 15521 8999 15524
rect 8941 15515 8999 15521
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4212 15456 4813 15484
rect 4212 15444 4218 15456
rect 4801 15453 4813 15456
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 8478 15484 8484 15496
rect 7515 15456 8484 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15484 9275 15487
rect 9766 15484 9772 15496
rect 9263 15456 9772 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 3510 15376 3516 15428
rect 3568 15416 3574 15428
rect 3786 15416 3792 15428
rect 3568 15388 3792 15416
rect 3568 15376 3574 15388
rect 3786 15376 3792 15388
rect 3844 15376 3850 15428
rect 8573 15419 8631 15425
rect 8573 15416 8585 15419
rect 5736 15388 8585 15416
rect 5736 15348 5764 15388
rect 8573 15385 8585 15388
rect 8619 15385 8631 15419
rect 8573 15379 8631 15385
rect 1964 15320 5764 15348
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 10060 15348 10088 15515
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 10928 15524 10977 15552
rect 10928 15512 10934 15524
rect 10965 15521 10977 15524
rect 11011 15552 11023 15555
rect 12342 15552 12348 15564
rect 11011 15524 12348 15552
rect 11011 15521 11023 15524
rect 10965 15515 11023 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 13357 15555 13415 15561
rect 13357 15552 13369 15555
rect 12860 15524 13369 15552
rect 12860 15512 12866 15524
rect 13357 15521 13369 15524
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 13538 15512 13544 15564
rect 13596 15552 13602 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 13596 15524 15669 15552
rect 13596 15512 13602 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15856 15552 15884 15592
rect 16016 15589 16028 15623
rect 16062 15620 16074 15623
rect 16666 15620 16672 15632
rect 16062 15592 16672 15620
rect 16062 15589 16074 15592
rect 16016 15583 16074 15589
rect 16666 15580 16672 15592
rect 16724 15580 16730 15632
rect 15856 15524 17540 15552
rect 15657 15515 15715 15521
rect 10226 15484 10232 15496
rect 10187 15456 10232 15484
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 13446 15484 13452 15496
rect 13407 15456 13452 15484
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13648 15416 13676 15447
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 14608 15456 14653 15484
rect 14608 15444 14614 15456
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15528 15456 15761 15484
rect 15528 15444 15534 15456
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 17402 15484 17408 15496
rect 17363 15456 17408 15484
rect 15749 15447 15807 15453
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 17512 15484 17540 15524
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18325 15555 18383 15561
rect 18325 15552 18337 15555
rect 18012 15524 18337 15552
rect 18012 15512 18018 15524
rect 18325 15521 18337 15524
rect 18371 15521 18383 15555
rect 18325 15515 18383 15521
rect 18417 15487 18475 15493
rect 18417 15484 18429 15487
rect 17512 15456 18429 15484
rect 18417 15453 18429 15456
rect 18463 15453 18475 15487
rect 18598 15484 18604 15496
rect 18511 15456 18604 15484
rect 18417 15447 18475 15453
rect 18598 15444 18604 15456
rect 18656 15484 18662 15496
rect 19242 15484 19248 15496
rect 18656 15456 19248 15484
rect 18656 15444 18662 15456
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 14568 15416 14596 15444
rect 13648 15388 14596 15416
rect 6696 15320 10088 15348
rect 6696 15308 6702 15320
rect 11882 15308 11888 15360
rect 11940 15348 11946 15360
rect 12345 15351 12403 15357
rect 12345 15348 12357 15351
rect 11940 15320 12357 15348
rect 11940 15308 11946 15320
rect 12345 15317 12357 15320
rect 12391 15317 12403 15351
rect 12345 15311 12403 15317
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 2682 15144 2688 15156
rect 1627 15116 2688 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 2958 15144 2964 15156
rect 2792 15116 2964 15144
rect 2792 15017 2820 15116
rect 2958 15104 2964 15116
rect 3016 15144 3022 15156
rect 4154 15144 4160 15156
rect 3016 15116 4160 15144
rect 3016 15104 3022 15116
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 5629 15147 5687 15153
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 5718 15144 5724 15156
rect 5675 15116 5724 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 5828 15116 9720 15144
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 5828 15076 5856 15116
rect 3844 15048 5856 15076
rect 9692 15076 9720 15116
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 9824 15116 10149 15144
rect 9824 15104 9830 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 13354 15144 13360 15156
rect 13315 15116 13360 15144
rect 10137 15107 10195 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 15746 15144 15752 15156
rect 13648 15116 15752 15144
rect 12894 15076 12900 15088
rect 9692 15048 12900 15076
rect 3844 15036 3850 15048
rect 12894 15036 12900 15048
rect 12952 15036 12958 15088
rect 2133 15011 2191 15017
rect 2133 15008 2145 15011
rect 1412 14980 2145 15008
rect 1412 14949 1440 14980
rect 2133 14977 2145 14980
rect 2179 14977 2191 15011
rect 2133 14971 2191 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 6178 15008 6184 15020
rect 6139 14980 6184 15008
rect 2777 14971 2835 14977
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 6270 14968 6276 15020
rect 6328 15008 6334 15020
rect 6328 14980 6684 15008
rect 6328 14968 6334 14980
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 1959 14943 2017 14949
rect 1959 14909 1971 14943
rect 2005 14909 2017 14943
rect 1959 14903 2017 14909
rect 3044 14943 3102 14949
rect 3044 14909 3056 14943
rect 3090 14940 3102 14943
rect 3970 14940 3976 14952
rect 3090 14912 3976 14940
rect 3090 14909 3102 14912
rect 3044 14903 3102 14909
rect 1964 14872 1992 14903
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6546 14940 6552 14952
rect 6135 14912 6552 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 6454 14872 6460 14884
rect 1964 14844 6460 14872
rect 6454 14832 6460 14844
rect 6512 14832 6518 14884
rect 6656 14872 6684 14980
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 8757 15011 8815 15017
rect 8757 15008 8769 15011
rect 8444 14980 8769 15008
rect 8444 14968 8450 14980
rect 8757 14977 8769 14980
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 11882 15008 11888 15020
rect 10008 14980 11744 15008
rect 11843 14980 11888 15008
rect 10008 14968 10014 14980
rect 6730 14900 6736 14952
rect 6788 14940 6794 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6788 14912 6837 14940
rect 6788 14900 6794 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 7092 14943 7150 14949
rect 7092 14909 7104 14943
rect 7138 14940 7150 14943
rect 8478 14940 8484 14952
rect 7138 14912 8484 14940
rect 7138 14909 7150 14912
rect 7092 14903 7150 14909
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 9024 14943 9082 14949
rect 9024 14909 9036 14943
rect 9070 14940 9082 14943
rect 9766 14940 9772 14952
rect 9070 14912 9772 14940
rect 9070 14909 9082 14912
rect 9024 14903 9082 14909
rect 9766 14900 9772 14912
rect 9824 14940 9830 14952
rect 10226 14940 10232 14952
rect 9824 14912 10232 14940
rect 9824 14900 9830 14912
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 11716 14940 11744 14980
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 11793 14943 11851 14949
rect 11793 14940 11805 14943
rect 11716 14912 11805 14940
rect 11793 14909 11805 14912
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 13648 14940 13676 15116
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 16574 15144 16580 15156
rect 16535 15116 16580 15144
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 19705 15147 19763 15153
rect 19705 15144 19717 15147
rect 18748 15116 19717 15144
rect 18748 15104 18754 15116
rect 19705 15113 19717 15116
rect 19751 15113 19763 15147
rect 19705 15107 19763 15113
rect 15194 15076 15200 15088
rect 14016 15048 15200 15076
rect 14016 15017 14044 15048
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 15470 15036 15476 15088
rect 15528 15076 15534 15088
rect 15528 15048 18368 15076
rect 15528 15036 15534 15048
rect 18340 15020 18368 15048
rect 14001 15011 14059 15017
rect 14001 14977 14013 15011
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 14608 14980 14933 15008
rect 14608 14968 14614 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 16209 15011 16267 15017
rect 16209 14977 16221 15011
rect 16255 15008 16267 15011
rect 16574 15008 16580 15020
rect 16255 14980 16580 15008
rect 16255 14977 16267 14980
rect 16209 14971 16267 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 17126 15008 17132 15020
rect 17087 14980 17132 15008
rect 17126 14968 17132 14980
rect 17184 14968 17190 15020
rect 18322 15008 18328 15020
rect 18235 14980 18328 15008
rect 18322 14968 18328 14980
rect 18380 14968 18386 15020
rect 12207 14912 13676 14940
rect 13725 14943 13783 14949
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 13725 14909 13737 14943
rect 13771 14940 13783 14943
rect 15010 14940 15016 14952
rect 13771 14912 15016 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15120 14912 16037 14940
rect 8570 14872 8576 14884
rect 6656 14844 8576 14872
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 8938 14832 8944 14884
rect 8996 14872 9002 14884
rect 11701 14875 11759 14881
rect 11701 14872 11713 14875
rect 8996 14844 11713 14872
rect 8996 14832 9002 14844
rect 11701 14841 11713 14844
rect 11747 14841 11759 14875
rect 11701 14835 11759 14841
rect 4154 14804 4160 14816
rect 4115 14776 4160 14804
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 5997 14807 6055 14813
rect 5997 14804 6009 14807
rect 5776 14776 6009 14804
rect 5776 14764 5782 14776
rect 5997 14773 6009 14776
rect 6043 14804 6055 14807
rect 6638 14804 6644 14816
rect 6043 14776 6644 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11606 14804 11612 14816
rect 11379 14776 11612 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11716 14804 11744 14835
rect 14458 14832 14464 14884
rect 14516 14872 14522 14884
rect 14829 14875 14887 14881
rect 14829 14872 14841 14875
rect 14516 14844 14841 14872
rect 14516 14832 14522 14844
rect 14829 14841 14841 14844
rect 14875 14872 14887 14875
rect 15120 14872 15148 14912
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 16945 14943 17003 14949
rect 16945 14909 16957 14943
rect 16991 14940 17003 14943
rect 17402 14940 17408 14952
rect 16991 14912 17408 14940
rect 16991 14909 17003 14912
rect 16945 14903 17003 14909
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 18598 14949 18604 14952
rect 18592 14940 18604 14949
rect 18559 14912 18604 14940
rect 18592 14903 18604 14912
rect 18598 14900 18604 14903
rect 18656 14900 18662 14952
rect 17037 14875 17095 14881
rect 17037 14872 17049 14875
rect 14875 14844 15148 14872
rect 15580 14844 17049 14872
rect 14875 14841 14887 14844
rect 14829 14835 14887 14841
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 11716 14776 12173 14804
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 13814 14804 13820 14816
rect 13775 14776 13820 14804
rect 12161 14767 12219 14773
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14182 14764 14188 14816
rect 14240 14804 14246 14816
rect 14369 14807 14427 14813
rect 14369 14804 14381 14807
rect 14240 14776 14381 14804
rect 14240 14764 14246 14776
rect 14369 14773 14381 14776
rect 14415 14773 14427 14807
rect 14369 14767 14427 14773
rect 14737 14807 14795 14813
rect 14737 14773 14749 14807
rect 14783 14804 14795 14807
rect 15102 14804 15108 14816
rect 14783 14776 15108 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15580 14813 15608 14844
rect 17037 14841 17049 14844
rect 17083 14841 17095 14875
rect 17037 14835 17095 14841
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14773 15623 14807
rect 15930 14804 15936 14816
rect 15891 14776 15936 14804
rect 15565 14767 15623 14773
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 1765 14603 1823 14609
rect 1765 14600 1777 14603
rect 1728 14572 1777 14600
rect 1728 14560 1734 14572
rect 1765 14569 1777 14572
rect 1811 14569 1823 14603
rect 2961 14603 3019 14609
rect 2961 14600 2973 14603
rect 1765 14563 1823 14569
rect 2516 14572 2973 14600
rect 1394 14492 1400 14544
rect 1452 14532 1458 14544
rect 2409 14535 2467 14541
rect 2409 14532 2421 14535
rect 1452 14504 2421 14532
rect 1452 14492 1458 14504
rect 2409 14501 2421 14504
rect 2455 14501 2467 14535
rect 2409 14495 2467 14501
rect 1578 14464 1584 14476
rect 1539 14436 1584 14464
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 2516 14464 2544 14572
rect 2961 14569 2973 14572
rect 3007 14569 3019 14603
rect 2961 14563 3019 14569
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14600 5503 14603
rect 7558 14600 7564 14612
rect 5491 14572 7564 14600
rect 5491 14569 5503 14572
rect 5445 14563 5503 14569
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4310 14535 4368 14541
rect 4310 14532 4322 14535
rect 4212 14504 4322 14532
rect 4212 14492 4218 14504
rect 4310 14501 4322 14504
rect 4356 14501 4368 14535
rect 4310 14495 4368 14501
rect 3326 14464 3332 14476
rect 2179 14436 2544 14464
rect 3287 14436 3332 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 3326 14424 3332 14436
rect 3384 14424 3390 14476
rect 5460 14464 5488 14563
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8757 14603 8815 14609
rect 8757 14600 8769 14603
rect 8352 14572 8769 14600
rect 8352 14560 8358 14572
rect 8757 14569 8769 14572
rect 8803 14569 8815 14603
rect 9674 14600 9680 14612
rect 9635 14572 9680 14600
rect 8757 14563 8815 14569
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 11974 14600 11980 14612
rect 11204 14572 11980 14600
rect 11204 14560 11210 14572
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 13262 14600 13268 14612
rect 12667 14572 13268 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 14829 14603 14887 14609
rect 14829 14569 14841 14603
rect 14875 14600 14887 14603
rect 15194 14600 15200 14612
rect 14875 14572 15200 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 17313 14603 17371 14609
rect 17313 14600 17325 14603
rect 15887 14572 17325 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 17313 14569 17325 14572
rect 17359 14569 17371 14603
rect 17313 14563 17371 14569
rect 6181 14535 6239 14541
rect 6181 14501 6193 14535
rect 6227 14532 6239 14535
rect 7190 14532 7196 14544
rect 6227 14504 7196 14532
rect 6227 14501 6239 14504
rect 6181 14495 6239 14501
rect 7190 14492 7196 14504
rect 7248 14492 7254 14544
rect 7282 14492 7288 14544
rect 7340 14532 7346 14544
rect 8665 14535 8723 14541
rect 8665 14532 8677 14535
rect 7340 14504 8677 14532
rect 7340 14492 7346 14504
rect 8665 14501 8677 14504
rect 8711 14501 8723 14535
rect 8665 14495 8723 14501
rect 10864 14535 10922 14541
rect 10864 14501 10876 14535
rect 10910 14532 10922 14535
rect 11882 14532 11888 14544
rect 10910 14504 11888 14532
rect 10910 14501 10922 14504
rect 10864 14495 10922 14501
rect 11882 14492 11888 14504
rect 11940 14532 11946 14544
rect 13280 14532 13308 14560
rect 15102 14532 15108 14544
rect 11940 14504 12848 14532
rect 13280 14504 15108 14532
rect 11940 14492 11946 14504
rect 6730 14464 6736 14476
rect 3620 14436 5488 14464
rect 6656 14436 6736 14464
rect 3418 14396 3424 14408
rect 3379 14368 3424 14396
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 3620 14405 3648 14436
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14365 3663 14399
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 3605 14359 3663 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 5074 14356 5080 14408
rect 5132 14396 5138 14408
rect 6656 14405 6684 14436
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 6908 14467 6966 14473
rect 6908 14433 6920 14467
rect 6954 14464 6966 14467
rect 8202 14464 8208 14476
rect 6954 14436 8208 14464
rect 6954 14433 6966 14436
rect 6908 14427 6966 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 12342 14464 12348 14476
rect 10643 14436 12348 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 12342 14424 12348 14436
rect 12400 14464 12406 14476
rect 12710 14464 12716 14476
rect 12400 14436 12572 14464
rect 12671 14436 12716 14464
rect 12400 14424 12406 14436
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 5132 14368 6653 14396
rect 5132 14356 5138 14368
rect 6641 14365 6653 14368
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 8220 14328 8248 14424
rect 8849 14399 8907 14405
rect 8849 14365 8861 14399
rect 8895 14365 8907 14399
rect 8849 14359 8907 14365
rect 8864 14328 8892 14359
rect 12544 14328 12572 14436
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 12820 14405 12848 14504
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 16206 14532 16212 14544
rect 16167 14504 16212 14532
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 18690 14541 18696 14544
rect 18684 14532 18696 14541
rect 18651 14504 18696 14532
rect 18684 14495 18696 14504
rect 18690 14492 18696 14495
rect 18748 14492 18754 14544
rect 13716 14467 13774 14473
rect 13716 14433 13728 14467
rect 13762 14464 13774 14467
rect 14458 14464 14464 14476
rect 13762 14436 14464 14464
rect 13762 14433 13774 14436
rect 13716 14427 13774 14433
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 15746 14424 15752 14476
rect 15804 14464 15810 14476
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 15804 14436 16313 14464
rect 15804 14424 15810 14436
rect 16301 14433 16313 14436
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 17865 14467 17923 14473
rect 17865 14464 17877 14467
rect 17267 14436 17877 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 17865 14433 17877 14436
rect 17911 14433 17923 14467
rect 17865 14427 17923 14433
rect 18322 14424 18328 14476
rect 18380 14464 18386 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 18380 14436 18429 14464
rect 18380 14424 18386 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 13464 14328 13492 14359
rect 8220 14300 8892 14328
rect 11808 14300 12388 14328
rect 12544 14300 13492 14328
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 6270 14260 6276 14272
rect 3660 14232 6276 14260
rect 3660 14220 3666 14232
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 6546 14220 6552 14272
rect 6604 14260 6610 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 6604 14232 8033 14260
rect 6604 14220 6610 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8294 14260 8300 14272
rect 8255 14232 8300 14260
rect 8021 14223 8079 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 11808 14260 11836 14300
rect 11974 14260 11980 14272
rect 8628 14232 11836 14260
rect 11935 14232 11980 14260
rect 8628 14220 8634 14232
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12250 14260 12256 14272
rect 12211 14232 12256 14260
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12360 14260 12388 14300
rect 15930 14260 15936 14272
rect 12360 14232 15936 14260
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16298 14220 16304 14272
rect 16356 14260 16362 14272
rect 16500 14260 16528 14359
rect 17402 14356 17408 14408
rect 17460 14396 17466 14408
rect 17460 14368 17505 14396
rect 17460 14356 17466 14368
rect 16850 14328 16856 14340
rect 16811 14300 16856 14328
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 19797 14263 19855 14269
rect 19797 14260 19809 14263
rect 16356 14232 19809 14260
rect 16356 14220 16362 14232
rect 19797 14229 19809 14232
rect 19843 14229 19855 14263
rect 19797 14223 19855 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1762 14056 1768 14068
rect 1627 14028 1768 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 3476 14028 3617 14056
rect 3476 14016 3482 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3605 14019 3663 14025
rect 3988 14028 5948 14056
rect 1578 13880 1584 13932
rect 1636 13920 1642 13932
rect 2133 13923 2191 13929
rect 2133 13920 2145 13923
rect 1636 13892 2145 13920
rect 1636 13880 1642 13892
rect 2133 13889 2145 13892
rect 2179 13889 2191 13923
rect 2133 13883 2191 13889
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3326 13920 3332 13932
rect 3191 13892 3332 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13852 2007 13855
rect 3988 13852 4016 14028
rect 5920 13988 5948 14028
rect 6178 14016 6184 14068
rect 6236 14056 6242 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6236 14028 6377 14056
rect 6236 14016 6242 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6365 14019 6423 14025
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6512 14028 6837 14056
rect 6512 14016 6518 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 7282 14056 7288 14068
rect 6825 14019 6883 14025
rect 7024 14028 7288 14056
rect 6914 13988 6920 14000
rect 5920 13960 6920 13988
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 4154 13920 4160 13932
rect 4115 13892 4160 13920
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 4982 13920 4988 13932
rect 4943 13892 4988 13920
rect 4982 13880 4988 13892
rect 5040 13880 5046 13932
rect 6730 13920 6736 13932
rect 6472 13892 6736 13920
rect 6472 13852 6500 13892
rect 6730 13880 6736 13892
rect 6788 13920 6794 13932
rect 7024 13920 7052 14028
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 9766 14056 9772 14068
rect 7616 14028 9352 14056
rect 9727 14028 9772 14056
rect 7616 14016 7622 14028
rect 8294 13988 8300 14000
rect 7300 13960 8300 13988
rect 7300 13929 7328 13960
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 9324 13988 9352 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 11882 14056 11888 14068
rect 9876 14028 11888 14056
rect 9876 13988 9904 14028
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 13538 14056 13544 14068
rect 13499 14028 13544 14056
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 9324 13960 9904 13988
rect 11149 13991 11207 13997
rect 11149 13957 11161 13991
rect 11195 13988 11207 13991
rect 12710 13988 12716 14000
rect 11195 13960 12716 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 6788 13892 7052 13920
rect 7285 13923 7343 13929
rect 6788 13880 6794 13892
rect 7285 13889 7297 13923
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 8386 13920 8392 13932
rect 8347 13892 8392 13920
rect 7377 13883 7435 13889
rect 1995 13824 4016 13852
rect 5184 13824 6500 13852
rect 1995 13821 2007 13824
rect 1949 13815 2007 13821
rect 3973 13787 4031 13793
rect 3973 13753 3985 13787
rect 4019 13784 4031 13787
rect 5184 13784 5212 13824
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 7392 13852 7420 13883
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 11790 13920 11796 13932
rect 11703 13892 11796 13920
rect 11790 13880 11796 13892
rect 11848 13920 11854 13932
rect 11974 13920 11980 13932
rect 11848 13892 11980 13920
rect 11848 13880 11854 13892
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 13078 13920 13084 13932
rect 13039 13892 13084 13920
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 14550 13920 14556 13932
rect 13556 13892 14412 13920
rect 14511 13892 14556 13920
rect 11517 13855 11575 13861
rect 6604 13824 7420 13852
rect 8588 13824 8984 13852
rect 6604 13812 6610 13824
rect 4019 13756 5212 13784
rect 5252 13787 5310 13793
rect 4019 13753 4031 13756
rect 3973 13747 4031 13753
rect 5252 13753 5264 13787
rect 5298 13784 5310 13787
rect 5442 13784 5448 13796
rect 5298 13756 5448 13784
rect 5298 13753 5310 13756
rect 5252 13747 5310 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 7190 13784 7196 13796
rect 7151 13756 7196 13784
rect 7190 13744 7196 13756
rect 7248 13744 7254 13796
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 8588 13784 8616 13824
rect 7340 13756 8616 13784
rect 8656 13787 8714 13793
rect 7340 13744 7346 13756
rect 8656 13753 8668 13787
rect 8702 13784 8714 13787
rect 8846 13784 8852 13796
rect 8702 13756 8852 13784
rect 8702 13753 8714 13756
rect 8656 13747 8714 13753
rect 8846 13744 8852 13756
rect 8904 13744 8910 13796
rect 8956 13784 8984 13824
rect 11517 13821 11529 13855
rect 11563 13852 11575 13855
rect 11606 13852 11612 13864
rect 11563 13824 11612 13852
rect 11563 13821 11575 13824
rect 11517 13815 11575 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12216 13824 13001 13852
rect 12216 13812 12222 13824
rect 12989 13821 13001 13824
rect 13035 13852 13047 13855
rect 13556 13852 13584 13892
rect 13722 13852 13728 13864
rect 13035 13824 13584 13852
rect 13683 13824 13728 13852
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14384 13861 14412 13892
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 16025 13923 16083 13929
rect 16025 13920 16037 13923
rect 15528 13892 16037 13920
rect 15528 13880 15534 13892
rect 16025 13889 16037 13892
rect 16071 13889 16083 13923
rect 16025 13883 16083 13889
rect 16298 13861 16304 13864
rect 14277 13855 14335 13861
rect 14277 13852 14289 13855
rect 14056 13824 14289 13852
rect 14056 13812 14062 13824
rect 14277 13821 14289 13824
rect 14323 13821 14335 13855
rect 14277 13815 14335 13821
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 16292 13852 16304 13861
rect 14415 13824 15240 13852
rect 16259 13824 16304 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 12802 13784 12808 13796
rect 8956 13756 12808 13784
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 12897 13787 12955 13793
rect 12897 13753 12909 13787
rect 12943 13784 12955 13787
rect 13446 13784 13452 13796
rect 12943 13756 13452 13784
rect 12943 13753 12955 13756
rect 12897 13747 12955 13753
rect 13446 13744 13452 13756
rect 13504 13744 13510 13796
rect 15212 13784 15240 13824
rect 16292 13815 16304 13824
rect 16298 13812 16304 13815
rect 16356 13812 16362 13864
rect 15654 13784 15660 13796
rect 15212 13756 15660 13784
rect 15654 13744 15660 13756
rect 15712 13784 15718 13796
rect 16206 13784 16212 13796
rect 15712 13756 16212 13784
rect 15712 13744 15718 13756
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 4065 13719 4123 13725
rect 4065 13716 4077 13719
rect 3936 13688 4077 13716
rect 3936 13676 3942 13688
rect 4065 13685 4077 13688
rect 4111 13685 4123 13719
rect 4065 13679 4123 13685
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 10226 13716 10232 13728
rect 4764 13688 10232 13716
rect 4764 13676 4770 13688
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 11609 13719 11667 13725
rect 11609 13685 11621 13719
rect 11655 13716 11667 13719
rect 12250 13716 12256 13728
rect 11655 13688 12256 13716
rect 11655 13685 11667 13688
rect 11609 13679 11667 13685
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 12526 13716 12532 13728
rect 12487 13688 12532 13716
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 13906 13716 13912 13728
rect 13867 13688 13912 13716
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5491 13484 6009 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 5997 13475 6055 13481
rect 6457 13515 6515 13521
rect 6457 13481 6469 13515
rect 6503 13512 6515 13515
rect 6822 13512 6828 13524
rect 6503 13484 6828 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 6972 13484 8217 13512
rect 6972 13472 6978 13484
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 12066 13512 12072 13524
rect 8205 13475 8263 13481
rect 9416 13484 12072 13512
rect 1394 13404 1400 13456
rect 1452 13444 1458 13456
rect 2317 13447 2375 13453
rect 2317 13444 2329 13447
rect 1452 13416 2329 13444
rect 1452 13404 1458 13416
rect 2317 13413 2329 13416
rect 2363 13413 2375 13447
rect 2317 13407 2375 13413
rect 4982 13404 4988 13456
rect 5040 13444 5046 13456
rect 5813 13447 5871 13453
rect 5813 13444 5825 13447
rect 5040 13416 5825 13444
rect 5040 13404 5046 13416
rect 5813 13413 5825 13416
rect 5859 13413 5871 13447
rect 8938 13444 8944 13456
rect 5813 13407 5871 13413
rect 7668 13416 8944 13444
rect 2051 13379 2109 13385
rect 2051 13345 2063 13379
rect 2097 13345 2109 13379
rect 2051 13339 2109 13345
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 6270 13376 6276 13388
rect 5399 13348 6276 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 2056 13240 2084 13339
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 7668 13376 7696 13416
rect 8938 13404 8944 13416
rect 8996 13404 9002 13456
rect 9416 13385 9444 13484
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 12492 13484 12633 13512
rect 12492 13472 12498 13484
rect 12621 13481 12633 13484
rect 12667 13481 12679 13515
rect 12621 13475 12679 13481
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 13081 13515 13139 13521
rect 13081 13512 13093 13515
rect 12768 13484 13093 13512
rect 12768 13472 12774 13484
rect 13081 13481 13093 13484
rect 13127 13481 13139 13515
rect 13814 13512 13820 13524
rect 13775 13484 13820 13512
rect 13081 13475 13139 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 13964 13484 14289 13512
rect 13964 13472 13970 13484
rect 14277 13481 14289 13484
rect 14323 13481 14335 13515
rect 14277 13475 14335 13481
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 15068 13484 15301 13512
rect 15068 13472 15074 13484
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 10137 13447 10195 13453
rect 10137 13413 10149 13447
rect 10183 13444 10195 13447
rect 10183 13416 11284 13444
rect 10183 13413 10195 13416
rect 10137 13407 10195 13413
rect 6411 13348 7696 13376
rect 7745 13379 7803 13385
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 7745 13345 7757 13379
rect 7791 13376 7803 13379
rect 8573 13379 8631 13385
rect 8573 13376 8585 13379
rect 7791 13348 8585 13376
rect 7791 13345 7803 13348
rect 7745 13339 7803 13345
rect 8573 13345 8585 13348
rect 8619 13345 8631 13379
rect 8573 13339 8631 13345
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13345 9459 13379
rect 10226 13376 10232 13388
rect 10187 13348 10232 13376
rect 9401 13339 9459 13345
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 10778 13376 10784 13388
rect 10739 13348 10784 13376
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 11256 13376 11284 13416
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 12989 13447 13047 13453
rect 12989 13444 13001 13447
rect 11664 13416 13001 13444
rect 11664 13404 11670 13416
rect 12989 13413 13001 13416
rect 13035 13413 13047 13447
rect 14182 13444 14188 13456
rect 14143 13416 14188 13444
rect 12989 13407 13047 13413
rect 14182 13404 14188 13416
rect 14240 13404 14246 13456
rect 17120 13447 17178 13453
rect 17120 13413 17132 13447
rect 17166 13444 17178 13447
rect 17402 13444 17408 13456
rect 17166 13416 17408 13444
rect 17166 13413 17178 13416
rect 17120 13407 17178 13413
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 12434 13376 12440 13388
rect 11256 13348 12440 13376
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 13814 13336 13820 13388
rect 13872 13376 13878 13388
rect 14090 13376 14096 13388
rect 13872 13348 14096 13376
rect 13872 13336 13878 13348
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 14826 13336 14832 13388
rect 14884 13376 14890 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14884 13348 15669 13376
rect 14884 13336 14890 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 16942 13376 16948 13388
rect 16899 13348 16948 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4120 13280 5120 13308
rect 4120 13268 4126 13280
rect 4985 13243 5043 13249
rect 4985 13240 4997 13243
rect 2056 13212 4997 13240
rect 4985 13209 4997 13212
rect 5031 13209 5043 13243
rect 5092 13240 5120 13280
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 5537 13311 5595 13317
rect 5537 13308 5549 13311
rect 5500 13280 5549 13308
rect 5500 13268 5506 13280
rect 5537 13277 5549 13280
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 5859 13280 6561 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 6549 13271 6607 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 8846 13308 8852 13320
rect 8807 13280 8852 13308
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 11054 13308 11060 13320
rect 10459 13280 11060 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 11054 13268 11060 13280
rect 11112 13308 11118 13320
rect 11790 13308 11796 13320
rect 11112 13280 11796 13308
rect 11112 13268 11118 13280
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 12032 13280 13185 13308
rect 12032 13268 12038 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 14366 13308 14372 13320
rect 14327 13280 14372 13308
rect 13173 13271 13231 13277
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 14458 13268 14464 13320
rect 14516 13308 14522 13320
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 14516 13280 15761 13308
rect 14516 13268 14522 13280
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 12618 13240 12624 13252
rect 5092 13212 12624 13240
rect 4985 13203 5043 13209
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 14384 13240 14412 13268
rect 15856 13240 15884 13271
rect 14384 13212 15884 13240
rect 4062 13132 4068 13184
rect 4120 13172 4126 13184
rect 7282 13172 7288 13184
rect 4120 13144 7288 13172
rect 4120 13132 4126 13144
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 9217 13175 9275 13181
rect 9217 13172 9229 13175
rect 7800 13144 9229 13172
rect 7800 13132 7806 13144
rect 9217 13141 9229 13144
rect 9263 13141 9275 13175
rect 9217 13135 9275 13141
rect 9769 13175 9827 13181
rect 9769 13141 9781 13175
rect 9815 13172 9827 13175
rect 11606 13172 11612 13184
rect 9815 13144 11612 13172
rect 9815 13141 9827 13144
rect 9769 13135 9827 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 13722 13172 13728 13184
rect 12124 13144 13728 13172
rect 12124 13132 12130 13144
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 18598 13172 18604 13184
rect 18279 13144 18604 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 2866 12968 2872 12980
rect 2547 12940 2872 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 5442 12928 5448 12980
rect 5500 12968 5506 12980
rect 6089 12971 6147 12977
rect 6089 12968 6101 12971
rect 5500 12940 6101 12968
rect 5500 12928 5506 12940
rect 6089 12937 6101 12940
rect 6135 12937 6147 12971
rect 6089 12931 6147 12937
rect 8846 12928 8852 12980
rect 8904 12968 8910 12980
rect 9493 12971 9551 12977
rect 9493 12968 9505 12971
rect 8904 12940 9505 12968
rect 8904 12928 8910 12940
rect 9493 12937 9505 12940
rect 9539 12937 9551 12971
rect 9493 12931 9551 12937
rect 14366 12928 14372 12980
rect 14424 12968 14430 12980
rect 14553 12971 14611 12977
rect 14553 12968 14565 12971
rect 14424 12940 14565 12968
rect 14424 12928 14430 12940
rect 14553 12937 14565 12940
rect 14599 12937 14611 12971
rect 14553 12931 14611 12937
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 16632 12940 16957 12968
rect 16632 12928 16638 12940
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 16945 12931 17003 12937
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3605 12903 3663 12909
rect 3605 12900 3617 12903
rect 2832 12872 3617 12900
rect 2832 12860 2838 12872
rect 3605 12869 3617 12872
rect 3651 12869 3663 12903
rect 3605 12863 3663 12869
rect 18049 12903 18107 12909
rect 18049 12869 18061 12903
rect 18095 12900 18107 12903
rect 19426 12900 19432 12912
rect 18095 12872 19432 12900
rect 18095 12869 18107 12872
rect 18049 12863 18107 12869
rect 19426 12860 19432 12872
rect 19484 12860 19490 12912
rect 4154 12832 4160 12844
rect 4115 12804 4160 12832
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6328 12804 6837 12832
rect 6328 12792 6334 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 7742 12832 7748 12844
rect 6825 12795 6883 12801
rect 7484 12804 7748 12832
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 1946 12764 1952 12776
rect 1811 12736 1952 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 2314 12764 2320 12776
rect 2275 12736 2320 12764
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 2866 12764 2872 12776
rect 2827 12736 2872 12764
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 7484 12773 7512 12804
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 12492 12804 12537 12832
rect 12492 12792 12498 12804
rect 14366 12792 14372 12844
rect 14424 12832 14430 12844
rect 14550 12832 14556 12844
rect 14424 12804 14556 12832
rect 14424 12792 14430 12804
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 14826 12832 14832 12844
rect 14787 12804 14832 12832
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 3936 12736 4721 12764
rect 3936 12724 3942 12736
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 8113 12767 8171 12773
rect 8113 12733 8125 12767
rect 8159 12764 8171 12767
rect 8202 12764 8208 12776
rect 8159 12736 8208 12764
rect 8159 12733 8171 12736
rect 8113 12727 8171 12733
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 11422 12764 11428 12776
rect 10643 12736 11428 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 11422 12724 11428 12736
rect 11480 12764 11486 12776
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 11480 12736 13185 12764
rect 11480 12724 11486 12736
rect 13173 12733 13185 12736
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 13440 12767 13498 12773
rect 13440 12733 13452 12767
rect 13486 12764 13498 12767
rect 14384 12764 14412 12792
rect 13486 12736 14412 12764
rect 15565 12767 15623 12773
rect 13486 12733 13498 12736
rect 13440 12727 13498 12733
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 16942 12764 16948 12776
rect 15611 12736 16948 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12764 18475 12767
rect 19702 12764 19708 12776
rect 18463 12736 19708 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 3973 12699 4031 12705
rect 3973 12665 3985 12699
rect 4019 12696 4031 12699
rect 4246 12696 4252 12708
rect 4019 12668 4252 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 4982 12705 4988 12708
rect 4976 12696 4988 12705
rect 4943 12668 4988 12696
rect 4976 12659 4988 12668
rect 5040 12696 5046 12708
rect 5350 12696 5356 12708
rect 5040 12668 5356 12696
rect 4982 12656 4988 12659
rect 5040 12656 5046 12668
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 8380 12699 8438 12705
rect 8380 12665 8392 12699
rect 8426 12696 8438 12699
rect 9122 12696 9128 12708
rect 8426 12668 9128 12696
rect 8426 12665 8438 12668
rect 8380 12659 8438 12665
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 10864 12699 10922 12705
rect 10864 12665 10876 12699
rect 10910 12696 10922 12699
rect 11054 12696 11060 12708
rect 10910 12668 11060 12696
rect 10910 12665 10922 12668
rect 10864 12659 10922 12665
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 15832 12699 15890 12705
rect 15832 12665 15844 12699
rect 15878 12696 15890 12699
rect 16114 12696 16120 12708
rect 15878 12668 16120 12696
rect 15878 12665 15890 12668
rect 15832 12659 15890 12665
rect 16114 12656 16120 12668
rect 16172 12656 16178 12708
rect 16206 12656 16212 12708
rect 16264 12696 16270 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 16264 12668 18521 12696
rect 16264 12656 16270 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 6822 12628 6828 12640
rect 4111 12600 6828 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7285 12631 7343 12637
rect 7285 12597 7297 12631
rect 7331 12628 7343 12631
rect 7558 12628 7564 12640
rect 7331 12600 7564 12628
rect 7331 12597 7343 12600
rect 7285 12591 7343 12597
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 11974 12628 11980 12640
rect 11935 12600 11980 12628
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 14182 12628 14188 12640
rect 13504 12600 14188 12628
rect 13504 12588 13510 12600
rect 14182 12588 14188 12600
rect 14240 12628 14246 12640
rect 18616 12628 18644 12736
rect 19702 12724 19708 12736
rect 19760 12724 19766 12776
rect 14240 12600 18644 12628
rect 14240 12588 14246 12600
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2056 12396 5120 12424
rect 2056 12297 2084 12396
rect 2314 12356 2320 12368
rect 2275 12328 2320 12356
rect 2314 12316 2320 12328
rect 2372 12316 2378 12368
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 3053 12359 3111 12365
rect 3053 12356 3065 12359
rect 2924 12328 3065 12356
rect 2924 12316 2930 12328
rect 3053 12325 3065 12328
rect 3099 12325 3111 12359
rect 3053 12319 3111 12325
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 4310 12359 4368 12365
rect 4310 12356 4322 12359
rect 4212 12328 4322 12356
rect 4212 12316 4218 12328
rect 4310 12325 4322 12328
rect 4356 12325 4368 12359
rect 5092 12356 5120 12396
rect 5350 12384 5356 12436
rect 5408 12424 5414 12436
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 5408 12396 5457 12424
rect 5408 12384 5414 12396
rect 5445 12393 5457 12396
rect 5491 12393 5503 12427
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 5445 12387 5503 12393
rect 5552 12396 7481 12424
rect 5552 12356 5580 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 7469 12387 7527 12393
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 8662 12424 8668 12436
rect 8619 12396 8668 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 14182 12424 14188 12436
rect 14143 12396 14188 12424
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15562 12424 15568 12436
rect 15519 12396 15568 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 16942 12424 16948 12436
rect 16855 12396 16948 12424
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 18966 12424 18972 12436
rect 18927 12396 18972 12424
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19426 12424 19432 12436
rect 19387 12396 19432 12424
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 5092 12328 5580 12356
rect 5988 12359 6046 12365
rect 4310 12319 4368 12325
rect 5988 12325 6000 12359
rect 6034 12356 6046 12359
rect 6546 12356 6552 12368
rect 6034 12328 6552 12356
rect 6034 12325 6046 12328
rect 5988 12319 6046 12325
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 11692 12359 11750 12365
rect 11692 12325 11704 12359
rect 11738 12356 11750 12359
rect 11974 12356 11980 12368
rect 11738 12328 11980 12356
rect 11738 12325 11750 12328
rect 11692 12319 11750 12325
rect 11974 12316 11980 12328
rect 12032 12316 12038 12368
rect 13538 12316 13544 12368
rect 13596 12356 13602 12368
rect 16960 12356 16988 12384
rect 17862 12356 17868 12368
rect 13596 12328 14964 12356
rect 16960 12328 17868 12356
rect 13596 12316 13602 12328
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 3694 12248 3700 12300
rect 3752 12288 3758 12300
rect 4706 12288 4712 12300
rect 3752 12260 4712 12288
rect 3752 12248 3758 12260
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 5810 12288 5816 12300
rect 5767 12260 5816 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 6454 12248 6460 12300
rect 6512 12288 6518 12300
rect 7837 12291 7895 12297
rect 7837 12288 7849 12291
rect 6512 12260 7849 12288
rect 6512 12248 6518 12260
rect 7837 12257 7849 12260
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8478 12288 8484 12300
rect 7975 12260 8484 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8938 12288 8944 12300
rect 8899 12260 8944 12288
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 9732 12260 10517 12288
rect 9732 12248 9738 12260
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 13078 12288 13084 12300
rect 10505 12251 10563 12257
rect 10796 12260 13084 12288
rect 10796 12232 10824 12260
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3936 12192 4077 12220
rect 3936 12180 3942 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8846 12220 8852 12232
rect 8159 12192 8852 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12189 10655 12223
rect 10778 12220 10784 12232
rect 10691 12192 10784 12220
rect 10597 12183 10655 12189
rect 10612 12152 10640 12183
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11422 12220 11428 12232
rect 11383 12192 11428 12220
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12820 12161 12848 12260
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 14090 12288 14096 12300
rect 14051 12260 14096 12288
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14936 12297 14964 12328
rect 17328 12297 17356 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 15887 12260 16497 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 17580 12291 17638 12297
rect 17580 12257 17592 12291
rect 17626 12288 17638 12291
rect 18598 12288 18604 12300
rect 17626 12260 18604 12288
rect 17626 12257 17638 12260
rect 17580 12251 17638 12257
rect 14366 12220 14372 12232
rect 14279 12192 14372 12220
rect 14366 12180 14372 12192
rect 14424 12220 14430 12232
rect 14734 12220 14740 12232
rect 14424 12192 14740 12220
rect 14424 12180 14430 12192
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15344 12192 15945 12220
rect 15344 12180 15350 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 15933 12183 15991 12189
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 6748 12124 10640 12152
rect 12805 12155 12863 12161
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 6748 12084 6776 12124
rect 12805 12121 12817 12155
rect 12851 12121 12863 12155
rect 12805 12115 12863 12121
rect 13725 12155 13783 12161
rect 13725 12121 13737 12155
rect 13771 12152 13783 12155
rect 14458 12152 14464 12164
rect 13771 12124 14464 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 14458 12112 14464 12124
rect 14516 12112 14522 12164
rect 17144 12152 17172 12251
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 19334 12288 19340 12300
rect 19295 12260 19340 12288
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 14752 12124 17172 12152
rect 18708 12192 19533 12220
rect 7098 12084 7104 12096
rect 4120 12056 6776 12084
rect 7059 12056 7104 12084
rect 4120 12044 4126 12056
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 10137 12087 10195 12093
rect 10137 12053 10149 12087
rect 10183 12084 10195 12087
rect 12618 12084 12624 12096
rect 10183 12056 12624 12084
rect 10183 12053 10195 12056
rect 10137 12047 10195 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 14752 12093 14780 12124
rect 18708 12096 18736 12192
rect 19521 12189 19533 12192
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 14737 12087 14795 12093
rect 14737 12084 14749 12087
rect 12768 12056 14749 12084
rect 12768 12044 12774 12056
rect 14737 12053 14749 12056
rect 14783 12053 14795 12087
rect 18690 12084 18696 12096
rect 18651 12056 18696 12084
rect 14737 12047 14795 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 3878 11880 3884 11892
rect 2792 11852 3884 11880
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2792 11753 2820 11852
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4154 11880 4160 11892
rect 4115 11852 4160 11880
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4304 11852 4445 11880
rect 4304 11840 4310 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 6822 11880 6828 11892
rect 6783 11852 6828 11880
rect 4433 11843 4491 11849
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 8202 11880 8208 11892
rect 7524 11852 8208 11880
rect 7524 11840 7530 11852
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 4028 11784 7512 11812
rect 4028 11772 4034 11784
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4212 11716 4905 11744
rect 4212 11704 4218 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11744 5043 11747
rect 7098 11744 7104 11756
rect 5031 11716 7104 11744
rect 5031 11713 5043 11716
rect 4985 11707 5043 11713
rect 1762 11676 1768 11688
rect 1723 11648 1768 11676
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 3044 11679 3102 11685
rect 3044 11645 3056 11679
rect 3090 11676 3102 11679
rect 5000 11676 5028 11707
rect 7098 11704 7104 11716
rect 7156 11744 7162 11756
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 7156 11716 7389 11744
rect 7156 11704 7162 11716
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 3090 11648 5028 11676
rect 3090 11645 3102 11648
rect 3044 11639 3102 11645
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 7064 11648 7297 11676
rect 7064 11636 7070 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7484 11676 7512 11784
rect 7944 11753 7972 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9309 11883 9367 11889
rect 9309 11880 9321 11883
rect 9180 11852 9321 11880
rect 9180 11840 9186 11852
rect 9309 11849 9321 11852
rect 9355 11849 9367 11883
rect 9309 11843 9367 11849
rect 11977 11883 12035 11889
rect 11977 11849 11989 11883
rect 12023 11880 12035 11883
rect 15194 11880 15200 11892
rect 12023 11852 13032 11880
rect 12023 11849 12035 11852
rect 11977 11843 12035 11849
rect 12710 11812 12716 11824
rect 12268 11784 12716 11812
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9732 11716 9777 11744
rect 9732 11704 9738 11716
rect 9030 11676 9036 11688
rect 7484 11648 9036 11676
rect 7285 11639 7343 11645
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 10008 11648 10149 11676
rect 10008 11636 10014 11648
rect 10137 11645 10149 11648
rect 10183 11645 10195 11679
rect 10137 11639 10195 11645
rect 10404 11679 10462 11685
rect 10404 11645 10416 11679
rect 10450 11676 10462 11679
rect 10778 11676 10784 11688
rect 10450 11648 10784 11676
rect 10450 11645 10462 11648
rect 10404 11639 10462 11645
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11974 11676 11980 11688
rect 10879 11648 11980 11676
rect 3326 11568 3332 11620
rect 3384 11608 3390 11620
rect 8196 11611 8254 11617
rect 3384 11580 7328 11608
rect 3384 11568 3390 11580
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4580 11512 4813 11540
rect 4580 11500 4586 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 7190 11540 7196 11552
rect 7151 11512 7196 11540
rect 4801 11503 4859 11509
rect 7190 11500 7196 11512
rect 7248 11500 7254 11552
rect 7300 11540 7328 11580
rect 8196 11577 8208 11611
rect 8242 11608 8254 11611
rect 8846 11608 8852 11620
rect 8242 11580 8852 11608
rect 8242 11577 8254 11580
rect 8196 11571 8254 11577
rect 8846 11568 8852 11580
rect 8904 11568 8910 11620
rect 10879 11540 10907 11648
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12268 11685 12296 11784
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 13004 11753 13032 11852
rect 13740 11852 15200 11880
rect 13740 11753 13768 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 17221 11883 17279 11889
rect 17221 11880 17233 11883
rect 16172 11852 17233 11880
rect 16172 11840 16178 11852
rect 17221 11849 17233 11852
rect 17267 11849 17279 11883
rect 17221 11843 17279 11849
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 19334 11880 19340 11892
rect 18095 11852 19340 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 15565 11815 15623 11821
rect 15565 11781 15577 11815
rect 15611 11812 15623 11815
rect 15657 11815 15715 11821
rect 15657 11812 15669 11815
rect 15611 11784 15669 11812
rect 15611 11781 15623 11784
rect 15565 11775 15623 11781
rect 15657 11781 15669 11784
rect 15703 11781 15715 11815
rect 15657 11775 15715 11781
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 17920 11784 19748 11812
rect 17920 11772 17926 11784
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12584 11716 12909 11744
rect 12584 11704 12590 11716
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11713 13783 11747
rect 18598 11744 18604 11756
rect 13725 11707 13783 11713
rect 15212 11716 15976 11744
rect 18559 11716 18604 11744
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 12253 11639 12311 11645
rect 12452 11648 13461 11676
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 11664 11580 12112 11608
rect 11664 11568 11670 11580
rect 7300 11512 10907 11540
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 12084 11549 12112 11580
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 11204 11512 11529 11540
rect 11204 11500 11210 11512
rect 11517 11509 11529 11512
rect 11563 11540 11575 11543
rect 11977 11543 12035 11549
rect 11977 11540 11989 11543
rect 11563 11512 11989 11540
rect 11563 11509 11575 11512
rect 11517 11503 11575 11509
rect 11977 11509 11989 11512
rect 12023 11509 12035 11543
rect 11977 11503 12035 11509
rect 12069 11543 12127 11549
rect 12069 11509 12081 11543
rect 12115 11540 12127 11543
rect 12158 11540 12164 11552
rect 12115 11512 12164 11540
rect 12115 11509 12127 11512
rect 12069 11503 12127 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12452 11549 12480 11648
rect 13449 11645 13461 11648
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14231 11648 14688 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 12676 11580 12817 11608
rect 12676 11568 12682 11580
rect 12805 11577 12817 11580
rect 12851 11577 12863 11611
rect 12805 11571 12863 11577
rect 14452 11611 14510 11617
rect 14452 11577 14464 11611
rect 14498 11608 14510 11611
rect 14550 11608 14556 11620
rect 14498 11580 14556 11608
rect 14498 11577 14510 11580
rect 14452 11571 14510 11577
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 14660 11608 14688 11648
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 15212 11676 15240 11716
rect 15746 11676 15752 11688
rect 14792 11648 15240 11676
rect 15304 11648 15752 11676
rect 14792 11636 14798 11648
rect 15304 11608 15332 11648
rect 15746 11636 15752 11648
rect 15804 11676 15810 11688
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 15804 11648 15853 11676
rect 15804 11636 15810 11648
rect 15841 11645 15853 11648
rect 15887 11645 15899 11679
rect 15948 11676 15976 11716
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 19720 11753 19748 11784
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 15948 11648 19012 11676
rect 15841 11639 15899 11645
rect 14660 11580 15332 11608
rect 15657 11611 15715 11617
rect 15657 11577 15669 11611
rect 15703 11608 15715 11611
rect 15930 11608 15936 11620
rect 15703 11580 15936 11608
rect 15703 11577 15715 11580
rect 15657 11571 15715 11577
rect 15930 11568 15936 11580
rect 15988 11608 15994 11620
rect 16086 11611 16144 11617
rect 16086 11608 16098 11611
rect 15988 11580 16098 11608
rect 15988 11568 15994 11580
rect 16086 11577 16098 11580
rect 16132 11577 16144 11611
rect 16086 11571 16144 11577
rect 17497 11611 17555 11617
rect 17497 11577 17509 11611
rect 17543 11608 17555 11611
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 17543 11580 18429 11608
rect 17543 11577 17555 11580
rect 17497 11571 17555 11577
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18417 11571 18475 11577
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11509 12495 11543
rect 12437 11503 12495 11509
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 18509 11543 18567 11549
rect 18509 11540 18521 11543
rect 13228 11512 18521 11540
rect 13228 11500 13234 11512
rect 18509 11509 18521 11512
rect 18555 11540 18567 11543
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18555 11512 18889 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18984 11540 19012 11648
rect 19978 11617 19984 11620
rect 19972 11608 19984 11617
rect 19939 11580 19984 11608
rect 19972 11571 19984 11580
rect 19978 11568 19984 11571
rect 20036 11568 20042 11620
rect 21085 11543 21143 11549
rect 21085 11540 21097 11543
rect 18984 11512 21097 11540
rect 18877 11503 18935 11509
rect 21085 11509 21097 11512
rect 21131 11509 21143 11543
rect 21085 11503 21143 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 2958 11336 2964 11348
rect 1627 11308 2964 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 4522 11336 4528 11348
rect 4483 11308 4528 11336
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 8846 11336 8852 11348
rect 7760 11308 8064 11336
rect 8807 11308 8852 11336
rect 4246 11268 4252 11280
rect 1964 11240 4252 11268
rect 1964 11209 1992 11240
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 6825 11271 6883 11277
rect 6825 11237 6837 11271
rect 6871 11268 6883 11271
rect 7760 11268 7788 11308
rect 6871 11240 7788 11268
rect 8036 11268 8064 11308
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 9088 11308 11161 11336
rect 9088 11296 9094 11308
rect 11149 11305 11161 11308
rect 11195 11305 11207 11339
rect 11149 11299 11207 11305
rect 11885 11339 11943 11345
rect 11885 11305 11897 11339
rect 11931 11305 11943 11339
rect 11885 11299 11943 11305
rect 9125 11271 9183 11277
rect 9125 11268 9137 11271
rect 8036 11240 9137 11268
rect 6871 11237 6883 11240
rect 6825 11231 6883 11237
rect 9125 11237 9137 11240
rect 9171 11237 9183 11271
rect 9125 11231 9183 11237
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11169 1455 11203
rect 1397 11163 1455 11169
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11169 2007 11203
rect 3234 11200 3240 11212
rect 3195 11172 3240 11200
rect 1949 11163 2007 11169
rect 1412 11132 1440 11163
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 3970 11200 3976 11212
rect 3375 11172 3976 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 7742 11209 7748 11212
rect 7736 11200 7748 11209
rect 7116 11172 7748 11200
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1412 11104 2145 11132
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 3694 11132 3700 11144
rect 3559 11104 3700 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 3694 11092 3700 11104
rect 3752 11092 3758 11144
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 7116 11141 7144 11172
rect 7736 11163 7748 11172
rect 7742 11160 7748 11163
rect 7800 11160 7806 11212
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11200 11299 11203
rect 11900 11200 11928 11299
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 13170 11336 13176 11348
rect 12032 11308 13176 11336
rect 12032 11296 12038 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 13998 11336 14004 11348
rect 13771 11308 14004 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 12253 11271 12311 11277
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 12434 11268 12440 11280
rect 12299 11240 12440 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 12434 11228 12440 11240
rect 12492 11228 12498 11280
rect 13280 11268 13308 11299
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 14458 11268 14464 11280
rect 13280 11240 14464 11268
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 15102 11228 15108 11280
rect 15160 11268 15166 11280
rect 15749 11271 15807 11277
rect 15749 11268 15761 11271
rect 15160 11240 15761 11268
rect 15160 11228 15166 11240
rect 15749 11237 15761 11240
rect 15795 11237 15807 11271
rect 15749 11231 15807 11237
rect 11287 11172 11836 11200
rect 11900 11172 12940 11200
rect 11287 11169 11299 11172
rect 11241 11163 11299 11169
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 4212 11104 6929 11132
rect 4212 11092 4218 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11101 7159 11135
rect 7466 11132 7472 11144
rect 7427 11104 7472 11132
rect 7101 11095 7159 11101
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11132 11483 11135
rect 11606 11132 11612 11144
rect 11471 11104 11612 11132
rect 11471 11101 11483 11104
rect 11425 11095 11483 11101
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 11808 11132 11836 11172
rect 12250 11132 12256 11144
rect 11808 11104 12256 11132
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12912 11132 12940 11172
rect 12986 11160 12992 11212
rect 13044 11200 13050 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 13044 11172 13645 11200
rect 13044 11160 13050 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 15654 11200 15660 11212
rect 15615 11172 15660 11200
rect 13633 11163 13691 11169
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 13722 11132 13728 11144
rect 12912 11104 13728 11132
rect 12437 11095 12495 11101
rect 6454 11064 6460 11076
rect 6415 11036 6460 11064
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 7190 11064 7196 11076
rect 6840 11036 7196 11064
rect 2866 10996 2872 11008
rect 2827 10968 2872 10996
rect 2866 10956 2872 10968
rect 2924 10956 2930 11008
rect 4890 10956 4896 11008
rect 4948 10996 4954 11008
rect 6840 10996 6868 11036
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 4948 10968 6868 10996
rect 4948 10956 4954 10968
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7484 10996 7512 11092
rect 10781 11067 10839 11073
rect 10781 11033 10793 11067
rect 10827 11064 10839 11067
rect 12360 11064 12388 11095
rect 10827 11036 12388 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 6972 10968 7512 10996
rect 6972 10956 6978 10968
rect 12342 10956 12348 11008
rect 12400 10996 12406 11008
rect 12452 10996 12480 11095
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11101 13875 11135
rect 15930 11132 15936 11144
rect 15891 11104 15936 11132
rect 13817 11095 13875 11101
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13832 11064 13860 11095
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 13504 11036 13860 11064
rect 13504 11024 13510 11036
rect 12400 10968 12480 10996
rect 12400 10956 12406 10968
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 1820 10764 2053 10792
rect 1820 10752 1826 10764
rect 2041 10761 2053 10764
rect 2087 10761 2099 10795
rect 7558 10792 7564 10804
rect 2041 10755 2099 10761
rect 6012 10764 7564 10792
rect 3053 10727 3111 10733
rect 3053 10724 3065 10727
rect 2516 10696 3065 10724
rect 2516 10656 2544 10696
rect 3053 10693 3065 10696
rect 3099 10693 3111 10727
rect 3053 10687 3111 10693
rect 2682 10656 2688 10668
rect 2424 10628 2544 10656
rect 2643 10628 2688 10656
rect 2424 10597 2452 10628
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3694 10656 3700 10668
rect 3655 10628 3700 10656
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4062 10656 4068 10668
rect 3936 10628 4068 10656
rect 3936 10616 3942 10628
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 4706 10656 4712 10668
rect 4667 10628 4712 10656
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2866 10588 2872 10600
rect 2547 10560 2872 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3510 10548 3516 10600
rect 3568 10588 3574 10600
rect 6012 10597 6040 10764
rect 7558 10752 7564 10764
rect 7616 10792 7622 10804
rect 7616 10764 8616 10792
rect 7616 10752 7622 10764
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7892 10696 8217 10724
rect 7892 10684 7898 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8478 10724 8484 10736
rect 8439 10696 8484 10724
rect 8205 10687 8263 10693
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 8220 10656 8248 10687
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 8588 10724 8616 10764
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 12986 10792 12992 10804
rect 8720 10764 12992 10792
rect 8720 10752 8726 10764
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 14550 10792 14556 10804
rect 14511 10764 14556 10792
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 9674 10724 9680 10736
rect 8588 10696 9680 10724
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 11425 10727 11483 10733
rect 11425 10693 11437 10727
rect 11471 10724 11483 10727
rect 11606 10724 11612 10736
rect 11471 10696 11612 10724
rect 11471 10693 11483 10696
rect 11425 10687 11483 10693
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8220 10628 9045 10656
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 9950 10656 9956 10668
rect 9640 10628 9956 10656
rect 9640 10616 9646 10628
rect 9950 10616 9956 10628
rect 10008 10656 10014 10668
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 10008 10628 10057 10656
rect 10008 10616 10014 10628
rect 10045 10625 10057 10628
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12492 10628 12537 10656
rect 12492 10616 12498 10628
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 17920 10628 18061 10656
rect 17920 10616 17926 10628
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 4525 10591 4583 10597
rect 4525 10588 4537 10591
rect 3568 10560 4537 10588
rect 3568 10548 3574 10560
rect 4525 10557 4537 10560
rect 4571 10557 4583 10591
rect 4525 10551 4583 10557
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10557 6055 10591
rect 5997 10551 6055 10557
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10312 10591 10370 10597
rect 9732 10560 9777 10588
rect 9732 10548 9738 10560
rect 10312 10557 10324 10591
rect 10358 10588 10370 10591
rect 11146 10588 11152 10600
rect 10358 10560 11152 10588
rect 10358 10557 10370 10560
rect 10312 10551 10370 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 12308 10560 13185 10588
rect 12308 10548 12314 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 15746 10588 15752 10600
rect 15659 10560 15752 10588
rect 13173 10551 13231 10557
rect 15746 10548 15752 10560
rect 15804 10588 15810 10600
rect 17880 10588 17908 10616
rect 15804 10560 17908 10588
rect 18316 10591 18374 10597
rect 15804 10548 15810 10560
rect 18316 10557 18328 10591
rect 18362 10588 18374 10591
rect 18690 10588 18696 10600
rect 18362 10560 18696 10588
rect 18362 10557 18374 10560
rect 18316 10551 18374 10557
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 7098 10529 7104 10532
rect 7092 10520 7104 10529
rect 7059 10492 7104 10520
rect 7092 10483 7104 10492
rect 7098 10480 7104 10483
rect 7156 10480 7162 10532
rect 7190 10480 7196 10532
rect 7248 10520 7254 10532
rect 8846 10520 8852 10532
rect 7248 10492 8852 10520
rect 7248 10480 7254 10492
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 8941 10523 8999 10529
rect 8941 10489 8953 10523
rect 8987 10520 8999 10523
rect 11698 10520 11704 10532
rect 8987 10492 11704 10520
rect 8987 10489 8999 10492
rect 8941 10483 8999 10489
rect 11698 10480 11704 10492
rect 11756 10480 11762 10532
rect 13446 10529 13452 10532
rect 13440 10520 13452 10529
rect 13407 10492 13452 10520
rect 13440 10483 13452 10492
rect 13446 10480 13452 10483
rect 13504 10480 13510 10532
rect 15654 10520 15660 10532
rect 14016 10492 15660 10520
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 3568 10424 3613 10452
rect 3568 10412 3574 10424
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 4028 10424 4077 10452
rect 4028 10412 4034 10424
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4890 10452 4896 10464
rect 4479 10424 4896 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5810 10452 5816 10464
rect 5771 10424 5816 10452
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 9306 10452 9312 10464
rect 8260 10424 9312 10452
rect 8260 10412 8266 10424
rect 9306 10412 9312 10424
rect 9364 10452 9370 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 9364 10424 9505 10452
rect 9364 10412 9370 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 14016 10452 14044 10492
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 16022 10529 16028 10532
rect 16016 10520 16028 10529
rect 15935 10492 16028 10520
rect 16016 10483 16028 10492
rect 16080 10520 16086 10532
rect 16080 10492 17540 10520
rect 16022 10480 16028 10483
rect 16080 10480 16086 10492
rect 9640 10424 14044 10452
rect 9640 10412 9646 10424
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 14829 10455 14887 10461
rect 14829 10452 14841 10455
rect 14424 10424 14841 10452
rect 14424 10412 14430 10424
rect 14829 10421 14841 10424
rect 14875 10421 14887 10455
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 14829 10415 14887 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17402 10452 17408 10464
rect 17363 10424 17408 10452
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17512 10452 17540 10492
rect 19429 10455 19487 10461
rect 19429 10452 19441 10455
rect 17512 10424 19441 10452
rect 19429 10421 19441 10424
rect 19475 10421 19487 10455
rect 19429 10415 19487 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 3752 10220 5457 10248
rect 3752 10208 3758 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 12342 10248 12348 10260
rect 5445 10211 5503 10217
rect 5552 10220 12112 10248
rect 12303 10220 12348 10248
rect 2032 10115 2090 10121
rect 2032 10081 2044 10115
rect 2078 10112 2090 10115
rect 3712 10112 3740 10208
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 5552 10180 5580 10220
rect 4028 10152 5580 10180
rect 8389 10183 8447 10189
rect 4028 10140 4034 10152
rect 8389 10149 8401 10183
rect 8435 10180 8447 10183
rect 9674 10180 9680 10192
rect 8435 10152 9680 10180
rect 8435 10149 8447 10152
rect 8389 10143 8447 10149
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 11232 10183 11290 10189
rect 11232 10149 11244 10183
rect 11278 10180 11290 10183
rect 11606 10180 11612 10192
rect 11278 10152 11612 10180
rect 11278 10149 11290 10152
rect 11232 10143 11290 10149
rect 11606 10140 11612 10152
rect 11664 10140 11670 10192
rect 4062 10112 4068 10124
rect 2078 10084 3740 10112
rect 4023 10084 4068 10112
rect 2078 10081 2090 10084
rect 2032 10075 2090 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4332 10115 4390 10121
rect 4332 10081 4344 10115
rect 4378 10112 4390 10115
rect 4706 10112 4712 10124
rect 4378 10084 4712 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 5810 10112 5816 10124
rect 5767 10084 5816 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 5988 10115 6046 10121
rect 5988 10081 6000 10115
rect 6034 10112 6046 10115
rect 8481 10115 8539 10121
rect 6034 10084 8064 10112
rect 6034 10081 6046 10084
rect 5988 10075 6046 10081
rect 1670 10004 1676 10056
rect 1728 10044 1734 10056
rect 1765 10047 1823 10053
rect 1765 10044 1777 10047
rect 1728 10016 1777 10044
rect 1728 10004 1734 10016
rect 1765 10013 1777 10016
rect 1811 10013 1823 10047
rect 8036 10044 8064 10084
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 10410 10112 10416 10124
rect 8527 10084 10416 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10112 11023 10115
rect 12084 10112 12112 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12584 10220 13032 10248
rect 12584 10208 12590 10220
rect 12360 10180 12388 10208
rect 12866 10183 12924 10189
rect 12866 10180 12878 10183
rect 12360 10152 12878 10180
rect 12866 10149 12878 10152
rect 12912 10149 12924 10183
rect 13004 10180 13032 10220
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 14001 10251 14059 10257
rect 14001 10248 14013 10251
rect 13504 10220 14013 10248
rect 13504 10208 13510 10220
rect 14001 10217 14013 10220
rect 14047 10217 14059 10251
rect 14001 10211 14059 10217
rect 15381 10251 15439 10257
rect 15381 10217 15393 10251
rect 15427 10248 15439 10251
rect 17034 10248 17040 10260
rect 15427 10220 17040 10248
rect 15427 10217 15439 10220
rect 15381 10211 15439 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 15841 10183 15899 10189
rect 15841 10180 15853 10183
rect 13004 10152 15853 10180
rect 12866 10143 12924 10149
rect 15841 10149 15853 10152
rect 15887 10149 15899 10183
rect 15841 10143 15899 10149
rect 16660 10183 16718 10189
rect 16660 10149 16672 10183
rect 16706 10180 16718 10183
rect 17126 10180 17132 10192
rect 16706 10152 17132 10180
rect 16706 10149 16718 10152
rect 16660 10143 16718 10149
rect 17126 10140 17132 10152
rect 17184 10140 17190 10192
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 11011 10084 12020 10112
rect 12084 10084 15761 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 8662 10044 8668 10056
rect 8036 10016 8668 10044
rect 1765 10007 1823 10013
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 11992 10044 12020 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 17862 10112 17868 10124
rect 16439 10084 17868 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 12250 10044 12256 10056
rect 11992 10016 12256 10044
rect 12250 10004 12256 10016
rect 12308 10044 12314 10056
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 12308 10016 12633 10044
rect 12308 10004 12314 10016
rect 12621 10013 12633 10016
rect 12667 10013 12679 10047
rect 16022 10044 16028 10056
rect 15983 10016 16028 10044
rect 12621 10007 12679 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 6656 9948 8156 9976
rect 2682 9868 2688 9920
rect 2740 9908 2746 9920
rect 3145 9911 3203 9917
rect 3145 9908 3157 9911
rect 2740 9880 3157 9908
rect 2740 9868 2746 9880
rect 3145 9877 3157 9880
rect 3191 9877 3203 9911
rect 3145 9871 3203 9877
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 6656 9908 6684 9948
rect 7098 9908 7104 9920
rect 4764 9880 6684 9908
rect 7059 9880 7104 9908
rect 4764 9868 4770 9880
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8128 9908 8156 9948
rect 13924 9948 15516 9976
rect 13924 9908 13952 9948
rect 8128 9880 13952 9908
rect 15488 9908 15516 9948
rect 17773 9911 17831 9917
rect 17773 9908 17785 9911
rect 15488 9880 17785 9908
rect 17773 9877 17785 9880
rect 17819 9877 17831 9911
rect 17773 9871 17831 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 3053 9707 3111 9713
rect 3053 9673 3065 9707
rect 3099 9704 3111 9707
rect 3510 9704 3516 9716
rect 3099 9676 3516 9704
rect 3099 9673 3111 9676
rect 3053 9667 3111 9673
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 8720 9676 9720 9704
rect 8720 9664 8726 9676
rect 3234 9596 3240 9648
rect 3292 9636 3298 9648
rect 4065 9639 4123 9645
rect 4065 9636 4077 9639
rect 3292 9608 4077 9636
rect 3292 9596 3298 9608
rect 4065 9605 4077 9608
rect 4111 9605 4123 9639
rect 4065 9599 4123 9605
rect 4246 9596 4252 9648
rect 4304 9636 4310 9648
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 4304 9608 5733 9636
rect 4304 9596 4310 9608
rect 5721 9605 5733 9608
rect 5767 9605 5779 9639
rect 5721 9599 5779 9605
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 4706 9568 4712 9580
rect 3743 9540 4712 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 7098 9568 7104 9580
rect 6411 9540 7104 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 8680 9568 8708 9664
rect 9692 9636 9720 9676
rect 10137 9639 10195 9645
rect 10137 9636 10149 9639
rect 9692 9608 10149 9636
rect 10137 9605 10149 9608
rect 10183 9605 10195 9639
rect 10410 9636 10416 9648
rect 10371 9608 10416 9636
rect 10137 9599 10195 9605
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 14001 9639 14059 9645
rect 14001 9605 14013 9639
rect 14047 9636 14059 9639
rect 14274 9636 14280 9648
rect 14047 9608 14280 9636
rect 14047 9605 14059 9608
rect 14001 9599 14059 9605
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 16577 9639 16635 9645
rect 16577 9605 16589 9639
rect 16623 9636 16635 9639
rect 16758 9636 16764 9648
rect 16623 9608 16764 9636
rect 16623 9605 16635 9608
rect 16577 9599 16635 9605
rect 16758 9596 16764 9608
rect 16816 9596 16822 9648
rect 7515 9540 8708 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10284 9540 10977 9568
rect 10284 9528 10290 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 14550 9568 14556 9580
rect 14511 9540 14556 9568
rect 10965 9531 11023 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 17126 9568 17132 9580
rect 17087 9540 17132 9568
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 4798 9500 4804 9512
rect 3559 9472 4804 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 4798 9460 4804 9472
rect 4856 9500 4862 9512
rect 4982 9500 4988 9512
rect 4856 9472 4988 9500
rect 4856 9460 4862 9472
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 8018 9500 8024 9512
rect 6227 9472 8024 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 8260 9472 8769 9500
rect 8260 9460 8266 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 9024 9503 9082 9509
rect 9024 9469 9036 9503
rect 9070 9500 9082 9503
rect 10244 9500 10272 9528
rect 14366 9500 14372 9512
rect 9070 9472 10272 9500
rect 14327 9472 14372 9500
rect 9070 9469 9082 9472
rect 9024 9463 9082 9469
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 17034 9500 17040 9512
rect 14516 9472 14561 9500
rect 16995 9472 17040 9500
rect 14516 9460 14522 9472
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 3234 9392 3240 9444
rect 3292 9432 3298 9444
rect 4433 9435 4491 9441
rect 3292 9404 4384 9432
rect 3292 9392 3298 9404
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9364 3482 9376
rect 4154 9364 4160 9376
rect 3476 9336 4160 9364
rect 3476 9324 3482 9336
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 4356 9364 4384 9404
rect 4433 9401 4445 9435
rect 4479 9432 4491 9435
rect 5534 9432 5540 9444
rect 4479 9404 5540 9432
rect 4479 9401 4491 9404
rect 4433 9395 4491 9401
rect 5534 9392 5540 9404
rect 5592 9432 5598 9444
rect 5994 9432 6000 9444
rect 5592 9404 6000 9432
rect 5592 9392 5598 9404
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 6135 9404 6868 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 4525 9367 4583 9373
rect 4525 9364 4537 9367
rect 4356 9336 4537 9364
rect 4525 9333 4537 9336
rect 4571 9364 4583 9367
rect 5718 9364 5724 9376
rect 4571 9336 5724 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 6840 9373 6868 9404
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 10873 9435 10931 9441
rect 7064 9404 7328 9432
rect 7064 9392 7070 9404
rect 7300 9376 7328 9404
rect 10873 9401 10885 9435
rect 10919 9432 10931 9435
rect 10962 9432 10968 9444
rect 10919 9404 10968 9432
rect 10919 9401 10931 9404
rect 10873 9395 10931 9401
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 16945 9435 17003 9441
rect 16945 9401 16957 9435
rect 16991 9432 17003 9435
rect 17402 9432 17408 9444
rect 16991 9404 17408 9432
rect 16991 9401 17003 9404
rect 16945 9395 17003 9401
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9333 6883 9367
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 6825 9327 6883 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7340 9336 7385 9364
rect 7340 9324 7346 9336
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8938 9364 8944 9376
rect 7800 9336 8944 9364
rect 7800 9324 7806 9336
rect 8938 9324 8944 9336
rect 8996 9364 9002 9376
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 8996 9336 10793 9364
rect 8996 9324 9002 9336
rect 10781 9333 10793 9336
rect 10827 9333 10839 9367
rect 10781 9327 10839 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1912 9132 1961 9160
rect 1912 9120 1918 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 1949 9123 2007 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 5074 9160 5080 9172
rect 4663 9132 5080 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 5074 9120 5080 9132
rect 5132 9160 5138 9172
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 5132 9132 5181 9160
rect 5132 9120 5138 9132
rect 5169 9129 5181 9132
rect 5215 9129 5227 9163
rect 5169 9123 5227 9129
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 7190 9160 7196 9172
rect 6411 9132 7196 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8202 9160 8208 9172
rect 7944 9132 8208 9160
rect 1762 9024 1768 9036
rect 1723 8996 1768 9024
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2317 9027 2375 9033
rect 2317 9024 2329 9027
rect 1912 8996 2329 9024
rect 1912 8984 1918 8996
rect 2317 8993 2329 8996
rect 2363 8993 2375 9027
rect 2317 8987 2375 8993
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 3660 8996 5089 9024
rect 3660 8984 3666 8996
rect 5077 8993 5089 8996
rect 5123 9024 5135 9027
rect 7742 9024 7748 9036
rect 5123 8996 7748 9024
rect 5123 8993 5135 8996
rect 5077 8987 5135 8993
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 7944 9033 7972 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10137 9095 10195 9101
rect 10137 9092 10149 9095
rect 8036 9064 10149 9092
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 3510 8916 3516 8968
rect 3568 8956 3574 8968
rect 5258 8956 5264 8968
rect 3568 8928 5264 8956
rect 3568 8916 3574 8928
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 8036 8956 8064 9064
rect 10137 9061 10149 9064
rect 10183 9061 10195 9095
rect 10137 9055 10195 9061
rect 8202 9033 8208 9036
rect 8196 9024 8208 9033
rect 8163 8996 8208 9024
rect 8196 8987 8208 8996
rect 8202 8984 8208 8987
rect 8260 8984 8266 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9398 9024 9404 9036
rect 8536 8996 9404 9024
rect 8536 8984 8542 8996
rect 9398 8984 9404 8996
rect 9456 9024 9462 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9456 8996 10057 9024
rect 9456 8984 9462 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 10226 8956 10232 8968
rect 6420 8928 8064 8956
rect 10187 8928 10232 8956
rect 6420 8916 6426 8928
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 9309 8891 9367 8897
rect 9309 8857 9321 8891
rect 9355 8888 9367 8891
rect 10244 8888 10272 8916
rect 9355 8860 10272 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 4706 8820 4712 8832
rect 4667 8792 4712 8820
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 17954 8820 17960 8832
rect 9640 8792 17960 8820
rect 9640 8780 9646 8792
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 4798 8616 4804 8628
rect 1412 8588 4804 8616
rect 1412 8421 1440 8588
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 4065 8551 4123 8557
rect 4065 8517 4077 8551
rect 4111 8548 4123 8551
rect 4522 8548 4528 8560
rect 4111 8520 4528 8548
rect 4111 8517 4123 8520
rect 4065 8511 4123 8517
rect 4522 8508 4528 8520
rect 4580 8508 4586 8560
rect 5074 8508 5080 8560
rect 5132 8548 5138 8560
rect 5810 8548 5816 8560
rect 5132 8520 5816 8548
rect 5132 8508 5138 8520
rect 5810 8508 5816 8520
rect 5868 8548 5874 8560
rect 6730 8548 6736 8560
rect 5868 8520 6736 8548
rect 5868 8508 5874 8520
rect 6730 8508 6736 8520
rect 6788 8548 6794 8560
rect 6788 8520 7144 8548
rect 6788 8508 6794 8520
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1854 8480 1860 8492
rect 1719 8452 1860 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4304 8452 4629 8480
rect 4304 8440 4310 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 5258 8440 5264 8492
rect 5316 8480 5322 8492
rect 7116 8489 7144 8520
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 8481 8551 8539 8557
rect 8481 8548 8493 8551
rect 8260 8520 8493 8548
rect 8260 8508 8266 8520
rect 8481 8517 8493 8520
rect 8527 8517 8539 8551
rect 8481 8511 8539 8517
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5316 8452 5641 8480
rect 5316 8440 5322 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 9306 8480 9312 8492
rect 9267 8452 9312 8480
rect 7101 8443 7159 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 2133 8415 2191 8421
rect 2133 8381 2145 8415
rect 2179 8381 2191 8415
rect 2133 8375 2191 8381
rect 2400 8415 2458 8421
rect 2400 8381 2412 8415
rect 2446 8412 2458 8415
rect 2682 8412 2688 8424
rect 2446 8384 2688 8412
rect 2446 8381 2458 8384
rect 2400 8375 2458 8381
rect 1670 8304 1676 8356
rect 1728 8344 1734 8356
rect 2148 8344 2176 8375
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 4706 8412 4712 8424
rect 4571 8384 4712 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8412 4951 8415
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 4939 8384 5549 8412
rect 4939 8381 4951 8384
rect 4893 8375 4951 8381
rect 5537 8381 5549 8384
rect 5583 8412 5595 8415
rect 6362 8412 6368 8424
rect 5583 8384 6368 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8904 8384 9137 8412
rect 8904 8372 8910 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8412 9275 8415
rect 9950 8412 9956 8424
rect 9263 8384 9956 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 2958 8344 2964 8356
rect 1728 8316 2964 8344
rect 1728 8304 1734 8316
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4433 8347 4491 8353
rect 3752 8316 4384 8344
rect 3752 8304 3758 8316
rect 3510 8276 3516 8288
rect 3471 8248 3516 8276
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 4356 8276 4384 8316
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 7368 8347 7426 8353
rect 4479 8316 5120 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 5092 8285 5120 8316
rect 7368 8313 7380 8347
rect 7414 8344 7426 8347
rect 7742 8344 7748 8356
rect 7414 8316 7748 8344
rect 7414 8313 7426 8316
rect 7368 8307 7426 8313
rect 7742 8304 7748 8316
rect 7800 8304 7806 8356
rect 4893 8279 4951 8285
rect 4893 8276 4905 8279
rect 4356 8248 4905 8276
rect 4893 8245 4905 8248
rect 4939 8245 4951 8279
rect 4893 8239 4951 8245
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8245 5135 8279
rect 5077 8239 5135 8245
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5316 8248 5457 8276
rect 5316 8236 5322 8248
rect 5445 8245 5457 8248
rect 5491 8276 5503 8279
rect 8478 8276 8484 8288
rect 5491 8248 8484 8276
rect 5491 8245 5503 8248
rect 5445 8239 5503 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8754 8276 8760 8288
rect 8715 8248 8760 8276
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 4522 8072 4528 8084
rect 4483 8044 4528 8072
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7800 8044 8125 8072
rect 7800 8032 7806 8044
rect 8113 8041 8125 8044
rect 8159 8072 8171 8075
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 8159 8044 8217 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 8849 8075 8907 8081
rect 8849 8072 8861 8075
rect 8812 8044 8861 8072
rect 8812 8032 8818 8044
rect 8849 8041 8861 8044
rect 8895 8041 8907 8075
rect 8849 8035 8907 8041
rect 18601 8075 18659 8081
rect 18601 8041 18613 8075
rect 18647 8072 18659 8075
rect 19518 8072 19524 8084
rect 18647 8044 19524 8072
rect 18647 8041 18659 8044
rect 18601 8035 18659 8041
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 1762 7964 1768 8016
rect 1820 8004 1826 8016
rect 2317 8007 2375 8013
rect 2317 8004 2329 8007
rect 1820 7976 2329 8004
rect 1820 7964 1826 7976
rect 2317 7973 2329 7976
rect 2363 7973 2375 8007
rect 2317 7967 2375 7973
rect 3878 7964 3884 8016
rect 3936 8004 3942 8016
rect 3936 7976 18460 8004
rect 3936 7964 3942 7976
rect 2030 7939 2088 7945
rect 2030 7936 2042 7939
rect 1964 7908 2042 7936
rect 1964 7732 1992 7908
rect 2030 7905 2042 7908
rect 2076 7905 2088 7939
rect 2030 7899 2088 7905
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 5350 7945 5356 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4212 7908 4445 7936
rect 4212 7896 4218 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 5344 7936 5356 7945
rect 4433 7899 4491 7905
rect 4724 7908 5356 7936
rect 4724 7877 4752 7908
rect 5344 7899 5356 7908
rect 5350 7896 5356 7899
rect 5408 7896 5414 7948
rect 7000 7939 7058 7945
rect 7000 7936 7012 7939
rect 6472 7908 7012 7936
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 5074 7868 5080 7880
rect 5035 7840 5080 7868
rect 4709 7831 4767 7837
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 6472 7809 6500 7908
rect 7000 7905 7012 7908
rect 7046 7936 7058 7939
rect 7046 7908 8064 7936
rect 7046 7905 7058 7908
rect 7000 7899 7058 7905
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 6457 7803 6515 7809
rect 6457 7769 6469 7803
rect 6503 7769 6515 7803
rect 8036 7800 8064 7908
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 18432 7945 18460 7976
rect 8757 7939 8815 7945
rect 8757 7936 8769 7939
rect 8352 7908 8769 7936
rect 8352 7896 8358 7908
rect 8757 7905 8769 7908
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 18423 7939 18481 7945
rect 18423 7905 18435 7939
rect 18469 7905 18481 7939
rect 18423 7899 18481 7905
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8251 7840 8953 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 8846 7800 8852 7812
rect 8036 7772 8852 7800
rect 6457 7763 6515 7769
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 1964 7704 4077 7732
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 4065 7695 4123 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4304 7500 4353 7528
rect 4304 7488 4310 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 2958 7392 2964 7404
rect 2919 7364 2964 7392
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 4356 7392 4384 7491
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5997 7531 6055 7537
rect 5997 7528 6009 7531
rect 5408 7500 6009 7528
rect 5408 7488 5414 7500
rect 5997 7497 6009 7500
rect 6043 7497 6055 7531
rect 5997 7491 6055 7497
rect 19153 7531 19211 7537
rect 19153 7497 19165 7531
rect 19199 7528 19211 7531
rect 19794 7528 19800 7540
rect 19199 7500 19800 7528
rect 19199 7497 19211 7500
rect 19153 7491 19211 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 5644 7432 8800 7460
rect 4356 7364 4752 7392
rect 2976 7256 3004 7352
rect 4724 7336 4752 7364
rect 3228 7327 3286 7333
rect 3228 7293 3240 7327
rect 3274 7324 3286 7327
rect 3510 7324 3516 7336
rect 3274 7296 3516 7324
rect 3274 7293 3286 7296
rect 3228 7287 3286 7293
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 4632 7256 4660 7287
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 4873 7327 4931 7333
rect 4873 7324 4885 7327
rect 4764 7296 4885 7324
rect 4764 7284 4770 7296
rect 4873 7293 4885 7296
rect 4919 7293 4931 7327
rect 4873 7287 4931 7293
rect 5074 7256 5080 7268
rect 2976 7228 5080 7256
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 5644 7256 5672 7432
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8772 7401 8800 7432
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7800 7364 7849 7392
rect 7800 7352 7806 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8846 7352 8852 7404
rect 8904 7392 8910 7404
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8904 7364 8953 7392
rect 8904 7352 8910 7364
rect 8941 7361 8953 7364
rect 8987 7392 8999 7395
rect 9306 7392 9312 7404
rect 8987 7364 9312 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 5500 7228 5672 7256
rect 5736 7296 8677 7324
rect 5500 7216 5506 7228
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 5736 7188 5764 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 12400 7296 18981 7324
rect 12400 7284 12406 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 6825 7259 6883 7265
rect 6825 7225 6837 7259
rect 6871 7256 6883 7259
rect 7653 7259 7711 7265
rect 7653 7256 7665 7259
rect 6871 7228 7665 7256
rect 6871 7225 6883 7228
rect 6825 7219 6883 7225
rect 7653 7225 7665 7228
rect 7699 7225 7711 7259
rect 7653 7219 7711 7225
rect 3476 7160 5764 7188
rect 7285 7191 7343 7197
rect 3476 7148 3482 7160
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7466 7188 7472 7200
rect 7331 7160 7472 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 7745 7191 7803 7197
rect 7745 7157 7757 7191
rect 7791 7188 7803 7191
rect 8297 7191 8355 7197
rect 8297 7188 8309 7191
rect 7791 7160 8309 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 8297 7157 8309 7160
rect 8343 7157 8355 7191
rect 8297 7151 8355 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5442 6984 5448 6996
rect 5040 6956 5448 6984
rect 5040 6944 5046 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 8573 6987 8631 6993
rect 8573 6984 8585 6987
rect 5592 6956 8585 6984
rect 5592 6944 5598 6956
rect 8573 6953 8585 6956
rect 8619 6953 8631 6987
rect 8573 6947 8631 6953
rect 5718 6876 5724 6928
rect 5776 6916 5782 6928
rect 8665 6919 8723 6925
rect 8665 6916 8677 6919
rect 5776 6888 8677 6916
rect 5776 6876 5782 6888
rect 8665 6885 8677 6888
rect 8711 6885 8723 6919
rect 8665 6879 8723 6885
rect 8754 6876 8760 6928
rect 8812 6916 8818 6928
rect 12342 6916 12348 6928
rect 8812 6888 12348 6916
rect 8812 6876 8818 6888
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 4479 6820 5089 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 7466 6848 7472 6860
rect 7427 6820 7472 6848
rect 5077 6811 5135 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 8386 6848 8392 6860
rect 7607 6820 8392 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 14568 6820 19441 6848
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 3936 6752 4537 6780
rect 3936 6740 3942 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 4525 6743 4583 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 8110 6780 8116 6792
rect 7791 6752 8116 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 8846 6780 8852 6792
rect 8807 6752 8852 6780
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 4065 6715 4123 6721
rect 4065 6681 4077 6715
rect 4111 6712 4123 6715
rect 4154 6712 4160 6724
rect 4111 6684 4160 6712
rect 4111 6681 4123 6684
rect 4065 6675 4123 6681
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 8205 6715 8263 6721
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 8294 6712 8300 6724
rect 8251 6684 8300 6712
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 7101 6647 7159 6653
rect 7101 6644 7113 6647
rect 4856 6616 7113 6644
rect 4856 6604 4862 6616
rect 7101 6613 7113 6616
rect 7147 6613 7159 6647
rect 7101 6607 7159 6613
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 14568 6644 14596 6820
rect 19429 6817 19441 6820
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 19610 6712 19616 6724
rect 19571 6684 19616 6712
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 7248 6616 14596 6644
rect 7248 6604 7254 6616
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 7282 6440 7288 6452
rect 3936 6412 7288 6440
rect 3936 6400 3942 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 20073 6443 20131 6449
rect 20073 6409 20085 6443
rect 20119 6440 20131 6443
rect 20714 6440 20720 6452
rect 20119 6412 20720 6440
rect 20119 6409 20131 6412
rect 20073 6403 20131 6409
rect 20714 6400 20720 6412
rect 20772 6400 20778 6452
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 19889 6239 19947 6245
rect 19889 6236 19901 6239
rect 4120 6208 19901 6236
rect 4120 6196 4126 6208
rect 19889 6205 19901 6208
rect 19935 6205 19947 6239
rect 19889 6199 19947 6205
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 20441 5899 20499 5905
rect 20441 5865 20453 5899
rect 20487 5896 20499 5899
rect 21174 5896 21180 5908
rect 20487 5868 21180 5896
rect 20487 5865 20499 5868
rect 20441 5859 20499 5865
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 4028 5732 20269 5760
rect 4028 5720 4034 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 14090 5352 14096 5364
rect 2924 5324 14096 5352
rect 2924 5312 2930 5324
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 20898 5352 20904 5364
rect 20763 5324 20904 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 4120 5120 20545 5148
rect 4120 5108 4126 5120
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4982 4128 4988 4140
rect 4028 4100 4988 4128
rect 4028 4088 4034 4100
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 5534 2020 5540 2032
rect 4120 1992 5540 2020
rect 4120 1980 4126 1992
rect 5534 1980 5540 1992
rect 5592 1980 5598 2032
rect 11422 1980 11428 2032
rect 11480 2020 11486 2032
rect 11882 2020 11888 2032
rect 11480 1992 11888 2020
rect 11480 1980 11486 1992
rect 11882 1980 11888 1992
rect 11940 1980 11946 2032
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2872 20000 2924 20052
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 9312 20000 9364 20052
rect 12900 20000 12952 20052
rect 14280 20000 14332 20052
rect 15660 20000 15712 20052
rect 16304 20000 16356 20052
rect 16856 20000 16908 20052
rect 18420 20000 18472 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 6000 19864 6052 19916
rect 9680 19864 9732 19916
rect 13084 19907 13136 19916
rect 13084 19873 13093 19907
rect 13093 19873 13127 19907
rect 13127 19873 13136 19907
rect 13084 19864 13136 19873
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 4896 19796 4948 19848
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 10048 19796 10100 19848
rect 2780 19728 2832 19780
rect 10968 19796 11020 19848
rect 14096 19796 14148 19848
rect 13268 19728 13320 19780
rect 15384 19864 15436 19916
rect 15660 19864 15712 19916
rect 16580 19907 16632 19916
rect 16580 19873 16589 19907
rect 16589 19873 16623 19907
rect 16623 19873 16632 19907
rect 16580 19864 16632 19873
rect 16672 19864 16724 19916
rect 18512 19864 18564 19916
rect 18604 19796 18656 19848
rect 15200 19728 15252 19780
rect 17040 19728 17092 19780
rect 2228 19660 2280 19712
rect 9772 19703 9824 19712
rect 9772 19669 9781 19703
rect 9781 19669 9815 19703
rect 9815 19669 9824 19703
rect 9772 19660 9824 19669
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3056 19456 3108 19508
rect 1768 19320 1820 19372
rect 20352 19363 20404 19372
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 204 19184 256 19236
rect 3056 19184 3108 19236
rect 2964 19116 3016 19168
rect 4988 19252 5040 19304
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 7656 19295 7708 19304
rect 5816 19184 5868 19236
rect 6828 19184 6880 19236
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 8760 19184 8812 19236
rect 3424 19116 3476 19168
rect 3608 19116 3660 19168
rect 4068 19116 4120 19168
rect 4160 19116 4212 19168
rect 4896 19116 4948 19168
rect 8208 19116 8260 19168
rect 9680 19252 9732 19304
rect 9956 19252 10008 19304
rect 12624 19295 12676 19304
rect 12624 19261 12633 19295
rect 12633 19261 12667 19295
rect 12667 19261 12676 19295
rect 12624 19252 12676 19261
rect 13360 19295 13412 19304
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 13820 19252 13872 19304
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 14372 19252 14424 19304
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 16304 19295 16356 19304
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 16856 19252 16908 19304
rect 17960 19252 18012 19304
rect 18972 19252 19024 19304
rect 22100 19252 22152 19304
rect 10140 19227 10192 19236
rect 10140 19193 10174 19227
rect 10174 19193 10192 19227
rect 10140 19184 10192 19193
rect 12072 19184 12124 19236
rect 10324 19116 10376 19168
rect 10968 19116 11020 19168
rect 13912 19184 13964 19236
rect 15660 19184 15712 19236
rect 16580 19184 16632 19236
rect 17408 19184 17460 19236
rect 18880 19184 18932 19236
rect 13452 19116 13504 19168
rect 15292 19116 15344 19168
rect 17592 19116 17644 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 2320 18844 2372 18896
rect 1492 18776 1544 18828
rect 1952 18819 2004 18828
rect 1952 18785 1961 18819
rect 1961 18785 1995 18819
rect 1995 18785 2004 18819
rect 1952 18776 2004 18785
rect 3240 18776 3292 18828
rect 5172 18912 5224 18964
rect 6828 18955 6880 18964
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 6920 18912 6972 18964
rect 11060 18912 11112 18964
rect 11704 18912 11756 18964
rect 12440 18912 12492 18964
rect 13084 18912 13136 18964
rect 14464 18912 14516 18964
rect 16028 18912 16080 18964
rect 5908 18844 5960 18896
rect 7104 18844 7156 18896
rect 10048 18844 10100 18896
rect 13268 18844 13320 18896
rect 13452 18887 13504 18896
rect 13452 18853 13461 18887
rect 13461 18853 13495 18887
rect 13495 18853 13504 18887
rect 13452 18844 13504 18853
rect 16304 18844 16356 18896
rect 16672 18887 16724 18896
rect 16672 18853 16681 18887
rect 16681 18853 16715 18887
rect 16715 18853 16724 18887
rect 16672 18844 16724 18853
rect 18972 18912 19024 18964
rect 18604 18844 18656 18896
rect 3516 18751 3568 18760
rect 3516 18717 3525 18751
rect 3525 18717 3559 18751
rect 3559 18717 3568 18751
rect 3516 18708 3568 18717
rect 4160 18708 4212 18760
rect 4988 18708 5040 18760
rect 9772 18776 9824 18828
rect 10324 18819 10376 18828
rect 10324 18785 10358 18819
rect 10358 18785 10376 18819
rect 10324 18776 10376 18785
rect 12440 18776 12492 18828
rect 12900 18776 12952 18828
rect 14096 18776 14148 18828
rect 15752 18819 15804 18828
rect 15752 18785 15761 18819
rect 15761 18785 15795 18819
rect 15795 18785 15804 18819
rect 15752 18776 15804 18785
rect 16580 18776 16632 18828
rect 16764 18776 16816 18828
rect 7748 18708 7800 18760
rect 8116 18751 8168 18760
rect 8116 18717 8125 18751
rect 8125 18717 8159 18751
rect 8159 18717 8168 18751
rect 8116 18708 8168 18717
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 8484 18708 8536 18760
rect 9956 18708 10008 18760
rect 13728 18708 13780 18760
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 18604 18708 18656 18760
rect 572 18640 624 18692
rect 2136 18572 2188 18624
rect 9680 18640 9732 18692
rect 12808 18640 12860 18692
rect 20352 18640 20404 18692
rect 7104 18572 7156 18624
rect 8760 18572 8812 18624
rect 14648 18572 14700 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18368 2004 18420
rect 8116 18368 8168 18420
rect 10140 18368 10192 18420
rect 13452 18368 13504 18420
rect 2136 18207 2188 18216
rect 2136 18173 2145 18207
rect 2145 18173 2179 18207
rect 2179 18173 2188 18207
rect 2136 18164 2188 18173
rect 4068 18232 4120 18284
rect 5724 18232 5776 18284
rect 5908 18275 5960 18284
rect 5908 18241 5917 18275
rect 5917 18241 5951 18275
rect 5951 18241 5960 18275
rect 5908 18232 5960 18241
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 8944 18232 8996 18284
rect 7104 18207 7156 18216
rect 1676 18096 1728 18148
rect 7104 18173 7113 18207
rect 7113 18173 7147 18207
rect 7147 18173 7156 18207
rect 7104 18164 7156 18173
rect 7748 18164 7800 18216
rect 4160 18096 4212 18148
rect 8852 18164 8904 18216
rect 9772 18164 9824 18216
rect 1768 18071 1820 18080
rect 1768 18037 1777 18071
rect 1777 18037 1811 18071
rect 1811 18037 1820 18071
rect 1768 18028 1820 18037
rect 2964 18028 3016 18080
rect 3424 18028 3476 18080
rect 3516 18028 3568 18080
rect 4068 18028 4120 18080
rect 5724 18071 5776 18080
rect 5724 18037 5733 18071
rect 5733 18037 5767 18071
rect 5767 18037 5776 18071
rect 5724 18028 5776 18037
rect 5816 18028 5868 18080
rect 7748 18028 7800 18080
rect 8392 18028 8444 18080
rect 9404 18096 9456 18148
rect 11888 18164 11940 18216
rect 9956 18096 10008 18148
rect 10232 18096 10284 18148
rect 10416 18096 10468 18148
rect 12164 18096 12216 18148
rect 13452 18232 13504 18284
rect 17868 18368 17920 18420
rect 18512 18232 18564 18284
rect 14648 18207 14700 18216
rect 14648 18173 14657 18207
rect 14657 18173 14691 18207
rect 14691 18173 14700 18207
rect 14648 18164 14700 18173
rect 17408 18207 17460 18216
rect 13084 18096 13136 18148
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 18972 18164 19024 18216
rect 15936 18096 15988 18148
rect 19708 18096 19760 18148
rect 22560 18096 22612 18148
rect 8944 18028 8996 18080
rect 9036 18028 9088 18080
rect 10692 18028 10744 18080
rect 10968 18028 11020 18080
rect 11612 18028 11664 18080
rect 13728 18028 13780 18080
rect 15292 18028 15344 18080
rect 15476 18028 15528 18080
rect 19616 18028 19668 18080
rect 20260 18028 20312 18080
rect 20904 18028 20956 18080
rect 21640 18028 21692 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 3240 17824 3292 17876
rect 5908 17824 5960 17876
rect 9864 17824 9916 17876
rect 12900 17824 12952 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15660 17867 15712 17876
rect 15660 17833 15669 17867
rect 15669 17833 15703 17867
rect 15703 17833 15712 17867
rect 15660 17824 15712 17833
rect 18604 17824 18656 17876
rect 9680 17756 9732 17808
rect 12716 17756 12768 17808
rect 2688 17731 2740 17740
rect 1584 17620 1636 17672
rect 2688 17697 2719 17731
rect 2719 17697 2740 17731
rect 2688 17688 2740 17697
rect 4988 17688 5040 17740
rect 6184 17688 6236 17740
rect 7012 17731 7064 17740
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7012 17688 7064 17697
rect 5172 17620 5224 17672
rect 6368 17620 6420 17672
rect 13176 17688 13228 17740
rect 13728 17756 13780 17808
rect 10416 17620 10468 17672
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 13084 17663 13136 17672
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 10140 17484 10192 17536
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 16948 17620 17000 17672
rect 19432 17620 19484 17672
rect 13452 17484 13504 17536
rect 14556 17484 14608 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 3148 17280 3200 17332
rect 3240 17280 3292 17332
rect 5724 17280 5776 17332
rect 1492 17144 1544 17196
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 6092 17187 6144 17196
rect 6092 17153 6101 17187
rect 6101 17153 6135 17187
rect 6135 17153 6144 17187
rect 6092 17144 6144 17153
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 4068 17076 4120 17128
rect 6368 17076 6420 17128
rect 7104 17008 7156 17060
rect 8208 17076 8260 17128
rect 8760 17076 8812 17128
rect 9772 17076 9824 17128
rect 12624 17280 12676 17332
rect 16948 17323 17000 17332
rect 16948 17289 16957 17323
rect 16957 17289 16991 17323
rect 16991 17289 17000 17323
rect 16948 17280 17000 17289
rect 11060 17212 11112 17264
rect 14464 17212 14516 17264
rect 12256 17144 12308 17196
rect 13176 17144 13228 17196
rect 16028 17144 16080 17196
rect 17592 17187 17644 17196
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 17868 17076 17920 17128
rect 7656 17008 7708 17060
rect 10416 17008 10468 17060
rect 4068 16940 4120 16992
rect 4160 16940 4212 16992
rect 8208 16940 8260 16992
rect 10048 16940 10100 16992
rect 10232 16940 10284 16992
rect 12532 16940 12584 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 19432 16983 19484 16992
rect 12900 16940 12952 16949
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 1584 16600 1636 16652
rect 3884 16736 3936 16788
rect 4252 16736 4304 16788
rect 6184 16736 6236 16788
rect 10048 16779 10100 16788
rect 5172 16668 5224 16720
rect 10048 16745 10057 16779
rect 10057 16745 10091 16779
rect 10091 16745 10100 16779
rect 10048 16736 10100 16745
rect 10140 16779 10192 16788
rect 10140 16745 10149 16779
rect 10149 16745 10183 16779
rect 10183 16745 10192 16779
rect 12532 16779 12584 16788
rect 10140 16736 10192 16745
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 12900 16736 12952 16788
rect 15936 16736 15988 16788
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 4252 16600 4304 16652
rect 5816 16600 5868 16652
rect 7196 16600 7248 16652
rect 8208 16600 8260 16652
rect 1400 16532 1452 16584
rect 3976 16532 4028 16584
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 8116 16532 8168 16584
rect 12900 16643 12952 16652
rect 12900 16609 12909 16643
rect 12909 16609 12943 16643
rect 12943 16609 12952 16643
rect 12900 16600 12952 16609
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 10876 16575 10928 16584
rect 10876 16541 10885 16575
rect 10885 16541 10919 16575
rect 10919 16541 10928 16575
rect 10876 16532 10928 16541
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 19432 16668 19484 16720
rect 13912 16643 13964 16652
rect 13912 16609 13921 16643
rect 13921 16609 13955 16643
rect 13955 16609 13964 16643
rect 13912 16600 13964 16609
rect 15200 16600 15252 16652
rect 16304 16600 16356 16652
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 14004 16575 14056 16584
rect 14004 16541 14013 16575
rect 14013 16541 14047 16575
rect 14047 16541 14056 16575
rect 14004 16532 14056 16541
rect 14740 16532 14792 16584
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 8760 16439 8812 16448
rect 8760 16405 8769 16439
rect 8769 16405 8803 16439
rect 8803 16405 8812 16439
rect 8760 16396 8812 16405
rect 12256 16439 12308 16448
rect 12256 16405 12265 16439
rect 12265 16405 12299 16439
rect 12299 16405 12308 16439
rect 12256 16396 12308 16405
rect 15476 16396 15528 16448
rect 19248 16439 19300 16448
rect 19248 16405 19257 16439
rect 19257 16405 19291 16439
rect 19291 16405 19300 16439
rect 19248 16396 19300 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2964 16192 3016 16244
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 10416 16235 10468 16244
rect 10416 16201 10425 16235
rect 10425 16201 10459 16235
rect 10459 16201 10468 16235
rect 10416 16192 10468 16201
rect 13084 16192 13136 16244
rect 14004 16192 14056 16244
rect 15476 16192 15528 16244
rect 4068 16124 4120 16176
rect 10784 16124 10836 16176
rect 12808 16124 12860 16176
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 5816 16099 5868 16108
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 4160 15988 4212 16040
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 7748 16056 7800 16108
rect 8208 16056 8260 16108
rect 12900 16099 12952 16108
rect 12900 16065 12909 16099
rect 12909 16065 12943 16099
rect 12943 16065 12952 16099
rect 12900 16056 12952 16065
rect 14740 16167 14792 16176
rect 14740 16133 14749 16167
rect 14749 16133 14783 16167
rect 14783 16133 14792 16167
rect 14740 16124 14792 16133
rect 17592 16192 17644 16244
rect 17960 16192 18012 16244
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 8392 15988 8444 16040
rect 8760 15988 8812 16040
rect 9772 15920 9824 15972
rect 11888 15920 11940 15972
rect 14556 15988 14608 16040
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 4896 15852 4948 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 7288 15852 7340 15904
rect 12348 15852 12400 15904
rect 15292 15920 15344 15972
rect 17132 15920 17184 15972
rect 17960 15920 18012 15972
rect 14004 15852 14056 15904
rect 15660 15852 15712 15904
rect 18420 15895 18472 15904
rect 18420 15861 18429 15895
rect 18429 15861 18463 15895
rect 18463 15861 18472 15895
rect 18420 15852 18472 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 2136 15648 2188 15700
rect 3240 15691 3292 15700
rect 3240 15657 3249 15691
rect 3249 15657 3283 15691
rect 3283 15657 3292 15691
rect 3240 15648 3292 15657
rect 5816 15648 5868 15700
rect 1768 15580 1820 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 4160 15444 4212 15496
rect 4988 15580 5040 15632
rect 7012 15648 7064 15700
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 7196 15623 7248 15632
rect 7196 15589 7205 15623
rect 7205 15589 7239 15623
rect 7239 15589 7248 15623
rect 7196 15580 7248 15589
rect 6184 15512 6236 15564
rect 8208 15648 8260 15700
rect 10324 15648 10376 15700
rect 12072 15648 12124 15700
rect 12992 15691 13044 15700
rect 12256 15580 12308 15632
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 13912 15648 13964 15700
rect 14464 15691 14516 15700
rect 14464 15657 14473 15691
rect 14473 15657 14507 15691
rect 14507 15657 14516 15691
rect 14464 15648 14516 15657
rect 15292 15648 15344 15700
rect 17132 15691 17184 15700
rect 17132 15657 17141 15691
rect 17141 15657 17175 15691
rect 17175 15657 17184 15691
rect 17132 15648 17184 15657
rect 17960 15691 18012 15700
rect 17960 15657 17969 15691
rect 17969 15657 18003 15691
rect 18003 15657 18012 15691
rect 17960 15648 18012 15657
rect 18420 15648 18472 15700
rect 15108 15580 15160 15632
rect 7932 15512 7984 15564
rect 9680 15512 9732 15564
rect 8484 15444 8536 15496
rect 9772 15444 9824 15496
rect 3516 15376 3568 15428
rect 3792 15376 3844 15428
rect 6644 15308 6696 15360
rect 10876 15512 10928 15564
rect 12348 15512 12400 15564
rect 12808 15512 12860 15564
rect 13544 15512 13596 15564
rect 16672 15580 16724 15632
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 14556 15487 14608 15496
rect 14556 15453 14565 15487
rect 14565 15453 14599 15487
rect 14599 15453 14608 15487
rect 14556 15444 14608 15453
rect 15476 15444 15528 15496
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 17960 15512 18012 15564
rect 18604 15487 18656 15496
rect 18604 15453 18613 15487
rect 18613 15453 18647 15487
rect 18647 15453 18656 15487
rect 18604 15444 18656 15453
rect 19248 15444 19300 15496
rect 11888 15308 11940 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2688 15104 2740 15156
rect 2964 15104 3016 15156
rect 4160 15104 4212 15156
rect 5724 15104 5776 15156
rect 3792 15036 3844 15088
rect 9772 15104 9824 15156
rect 13360 15147 13412 15156
rect 13360 15113 13369 15147
rect 13369 15113 13403 15147
rect 13403 15113 13412 15147
rect 13360 15104 13412 15113
rect 12900 15036 12952 15088
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 6276 14968 6328 15020
rect 3976 14900 4028 14952
rect 6552 14900 6604 14952
rect 6460 14832 6512 14884
rect 8392 14968 8444 15020
rect 9956 14968 10008 15020
rect 11888 15011 11940 15020
rect 6736 14900 6788 14952
rect 8484 14900 8536 14952
rect 9772 14900 9824 14952
rect 10232 14900 10284 14952
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 15752 15104 15804 15156
rect 16580 15147 16632 15156
rect 16580 15113 16589 15147
rect 16589 15113 16623 15147
rect 16623 15113 16632 15147
rect 16580 15104 16632 15113
rect 18696 15104 18748 15156
rect 15200 15036 15252 15088
rect 15476 15036 15528 15088
rect 14556 14968 14608 15020
rect 16580 14968 16632 15020
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 15016 14900 15068 14952
rect 8576 14832 8628 14884
rect 8944 14832 8996 14884
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 5724 14764 5776 14816
rect 6644 14764 6696 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 11612 14764 11664 14816
rect 14464 14832 14516 14884
rect 17408 14900 17460 14952
rect 18604 14943 18656 14952
rect 18604 14909 18638 14943
rect 18638 14909 18656 14943
rect 18604 14900 18656 14909
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 14188 14764 14240 14816
rect 15108 14764 15160 14816
rect 15936 14807 15988 14816
rect 15936 14773 15945 14807
rect 15945 14773 15979 14807
rect 15979 14773 15988 14807
rect 15936 14764 15988 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14560 1728 14612
rect 1400 14492 1452 14544
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 4160 14492 4212 14544
rect 3332 14467 3384 14476
rect 3332 14433 3341 14467
rect 3341 14433 3375 14467
rect 3375 14433 3384 14467
rect 3332 14424 3384 14433
rect 7564 14560 7616 14612
rect 8300 14560 8352 14612
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 11152 14560 11204 14612
rect 11980 14560 12032 14612
rect 13268 14560 13320 14612
rect 15200 14560 15252 14612
rect 7196 14492 7248 14544
rect 7288 14492 7340 14544
rect 11888 14492 11940 14544
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 5080 14356 5132 14408
rect 6736 14424 6788 14476
rect 8208 14424 8260 14476
rect 12348 14424 12400 14476
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 15108 14492 15160 14544
rect 16212 14535 16264 14544
rect 16212 14501 16221 14535
rect 16221 14501 16255 14535
rect 16255 14501 16264 14535
rect 16212 14492 16264 14501
rect 18696 14535 18748 14544
rect 18696 14501 18730 14535
rect 18730 14501 18748 14535
rect 18696 14492 18748 14501
rect 14464 14424 14516 14476
rect 15752 14424 15804 14476
rect 18328 14424 18380 14476
rect 3608 14220 3660 14272
rect 6276 14220 6328 14272
rect 6552 14220 6604 14272
rect 8300 14263 8352 14272
rect 8300 14229 8309 14263
rect 8309 14229 8343 14263
rect 8343 14229 8352 14263
rect 8300 14220 8352 14229
rect 8576 14220 8628 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 15936 14220 15988 14272
rect 16304 14220 16356 14272
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 16856 14331 16908 14340
rect 16856 14297 16865 14331
rect 16865 14297 16899 14331
rect 16899 14297 16908 14331
rect 16856 14288 16908 14297
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1768 14016 1820 14068
rect 3424 14016 3476 14068
rect 1584 13880 1636 13932
rect 3332 13880 3384 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 6184 14016 6236 14068
rect 6460 14016 6512 14068
rect 6920 13948 6972 14000
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 4988 13923 5040 13932
rect 4988 13889 4997 13923
rect 4997 13889 5031 13923
rect 5031 13889 5040 13923
rect 4988 13880 5040 13889
rect 6736 13880 6788 13932
rect 7288 14016 7340 14068
rect 7564 14016 7616 14068
rect 9772 14059 9824 14068
rect 8300 13948 8352 14000
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 11888 14016 11940 14068
rect 13544 14059 13596 14068
rect 13544 14025 13553 14059
rect 13553 14025 13587 14059
rect 13587 14025 13596 14059
rect 13544 14016 13596 14025
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 12716 13948 12768 14000
rect 8392 13923 8444 13932
rect 6552 13812 6604 13864
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 11980 13880 12032 13932
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 14556 13923 14608 13932
rect 5448 13744 5500 13796
rect 7196 13787 7248 13796
rect 7196 13753 7205 13787
rect 7205 13753 7239 13787
rect 7239 13753 7248 13787
rect 7196 13744 7248 13753
rect 7288 13744 7340 13796
rect 8852 13744 8904 13796
rect 11612 13812 11664 13864
rect 12164 13812 12216 13864
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 14004 13812 14056 13864
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 15476 13880 15528 13932
rect 16304 13855 16356 13864
rect 12808 13744 12860 13796
rect 13452 13744 13504 13796
rect 16304 13821 16338 13855
rect 16338 13821 16356 13855
rect 16304 13812 16356 13821
rect 15660 13744 15712 13796
rect 16212 13744 16264 13796
rect 3884 13676 3936 13728
rect 4712 13676 4764 13728
rect 10232 13676 10284 13728
rect 12256 13676 12308 13728
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 13912 13719 13964 13728
rect 13912 13685 13921 13719
rect 13921 13685 13955 13719
rect 13955 13685 13964 13719
rect 13912 13676 13964 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 6828 13472 6880 13524
rect 6920 13472 6972 13524
rect 12072 13515 12124 13524
rect 1400 13404 1452 13456
rect 4988 13404 5040 13456
rect 6276 13336 6328 13388
rect 8944 13404 8996 13456
rect 12072 13481 12081 13515
rect 12081 13481 12115 13515
rect 12115 13481 12124 13515
rect 12072 13472 12124 13481
rect 12440 13472 12492 13524
rect 12716 13472 12768 13524
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 13912 13472 13964 13524
rect 15016 13472 15068 13524
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 10784 13379 10836 13388
rect 10784 13345 10793 13379
rect 10793 13345 10827 13379
rect 10827 13345 10836 13379
rect 10784 13336 10836 13345
rect 11612 13404 11664 13456
rect 14188 13447 14240 13456
rect 14188 13413 14197 13447
rect 14197 13413 14231 13447
rect 14231 13413 14240 13447
rect 14188 13404 14240 13413
rect 17408 13404 17460 13456
rect 12440 13336 12492 13388
rect 13820 13336 13872 13388
rect 14096 13336 14148 13388
rect 14832 13336 14884 13388
rect 16948 13336 17000 13388
rect 4068 13268 4120 13320
rect 5448 13268 5500 13320
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 8852 13311 8904 13320
rect 8852 13277 8861 13311
rect 8861 13277 8895 13311
rect 8895 13277 8904 13311
rect 8852 13268 8904 13277
rect 11060 13268 11112 13320
rect 11796 13268 11848 13320
rect 11980 13268 12032 13320
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 14464 13268 14516 13320
rect 12624 13200 12676 13252
rect 4068 13132 4120 13184
rect 7288 13132 7340 13184
rect 7748 13132 7800 13184
rect 11612 13132 11664 13184
rect 12072 13132 12124 13184
rect 13728 13132 13780 13184
rect 18604 13132 18656 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 2872 12928 2924 12980
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 5448 12928 5500 12980
rect 8852 12928 8904 12980
rect 14372 12928 14424 12980
rect 16580 12928 16632 12980
rect 2780 12860 2832 12912
rect 19432 12860 19484 12912
rect 4160 12835 4212 12844
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 6276 12792 6328 12844
rect 1952 12724 2004 12776
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 3884 12724 3936 12776
rect 7748 12792 7800 12844
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 14372 12792 14424 12844
rect 14556 12792 14608 12844
rect 14832 12835 14884 12844
rect 14832 12801 14841 12835
rect 14841 12801 14875 12835
rect 14875 12801 14884 12835
rect 14832 12792 14884 12801
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 8208 12724 8260 12776
rect 11428 12724 11480 12776
rect 16948 12724 17000 12776
rect 4252 12656 4304 12708
rect 4988 12699 5040 12708
rect 4988 12665 5022 12699
rect 5022 12665 5040 12699
rect 4988 12656 5040 12665
rect 5356 12656 5408 12708
rect 9128 12656 9180 12708
rect 11060 12656 11112 12708
rect 16120 12656 16172 12708
rect 16212 12656 16264 12708
rect 6828 12588 6880 12640
rect 7564 12588 7616 12640
rect 11980 12631 12032 12640
rect 11980 12597 11989 12631
rect 11989 12597 12023 12631
rect 12023 12597 12032 12631
rect 11980 12588 12032 12597
rect 13452 12588 13504 12640
rect 14188 12588 14240 12640
rect 19708 12724 19760 12776
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2320 12359 2372 12368
rect 2320 12325 2329 12359
rect 2329 12325 2363 12359
rect 2363 12325 2372 12359
rect 2320 12316 2372 12325
rect 2872 12316 2924 12368
rect 4160 12316 4212 12368
rect 5356 12384 5408 12436
rect 8668 12384 8720 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 14188 12427 14240 12436
rect 14188 12393 14197 12427
rect 14197 12393 14231 12427
rect 14231 12393 14240 12427
rect 14188 12384 14240 12393
rect 15568 12384 15620 12436
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 18972 12427 19024 12436
rect 18972 12393 18981 12427
rect 18981 12393 19015 12427
rect 19015 12393 19024 12427
rect 18972 12384 19024 12393
rect 19432 12427 19484 12436
rect 19432 12393 19441 12427
rect 19441 12393 19475 12427
rect 19475 12393 19484 12427
rect 19432 12384 19484 12393
rect 6552 12316 6604 12368
rect 11980 12316 12032 12368
rect 13544 12316 13596 12368
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 3700 12248 3752 12300
rect 4712 12248 4764 12300
rect 5816 12248 5868 12300
rect 6460 12248 6512 12300
rect 8484 12248 8536 12300
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 9680 12248 9732 12300
rect 3884 12180 3936 12232
rect 8852 12180 8904 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 13084 12248 13136 12300
rect 14096 12291 14148 12300
rect 14096 12257 14105 12291
rect 14105 12257 14139 12291
rect 14139 12257 14148 12291
rect 14096 12248 14148 12257
rect 17868 12316 17920 12368
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 14740 12180 14792 12232
rect 15292 12180 15344 12232
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 4068 12044 4120 12096
rect 14464 12112 14516 12164
rect 18604 12248 18656 12300
rect 19340 12291 19392 12300
rect 19340 12257 19349 12291
rect 19349 12257 19383 12291
rect 19383 12257 19392 12291
rect 19340 12248 19392 12257
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 12624 12044 12676 12096
rect 12716 12044 12768 12096
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 3884 11840 3936 11892
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 4252 11840 4304 11892
rect 6828 11883 6880 11892
rect 6828 11849 6837 11883
rect 6837 11849 6871 11883
rect 6871 11849 6880 11883
rect 6828 11840 6880 11849
rect 7472 11840 7524 11892
rect 3976 11772 4028 11824
rect 4160 11704 4212 11756
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 7104 11704 7156 11756
rect 7012 11636 7064 11688
rect 8208 11840 8260 11892
rect 9128 11840 9180 11892
rect 9680 11747 9732 11756
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 9036 11636 9088 11688
rect 9956 11636 10008 11688
rect 10784 11636 10836 11688
rect 3332 11568 3384 11620
rect 4528 11500 4580 11552
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 8852 11568 8904 11620
rect 11980 11636 12032 11688
rect 12716 11772 12768 11824
rect 12532 11704 12584 11756
rect 15200 11840 15252 11892
rect 16120 11840 16172 11892
rect 19340 11840 19392 11892
rect 17868 11772 17920 11824
rect 18604 11747 18656 11756
rect 11612 11568 11664 11620
rect 11152 11500 11204 11552
rect 12164 11500 12216 11552
rect 12624 11568 12676 11620
rect 14556 11568 14608 11620
rect 14740 11636 14792 11688
rect 15752 11636 15804 11688
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 15936 11568 15988 11620
rect 13176 11500 13228 11552
rect 19984 11611 20036 11620
rect 19984 11577 20018 11611
rect 20018 11577 20036 11611
rect 19984 11568 20036 11577
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2964 11296 3016 11348
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 8852 11339 8904 11348
rect 4252 11228 4304 11280
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 9036 11296 9088 11348
rect 3240 11203 3292 11212
rect 3240 11169 3249 11203
rect 3249 11169 3283 11203
rect 3283 11169 3292 11203
rect 3240 11160 3292 11169
rect 3976 11160 4028 11212
rect 7748 11203 7800 11212
rect 3700 11092 3752 11144
rect 4160 11092 4212 11144
rect 7748 11169 7782 11203
rect 7782 11169 7800 11203
rect 7748 11160 7800 11169
rect 11980 11296 12032 11348
rect 13176 11296 13228 11348
rect 12440 11228 12492 11280
rect 14004 11296 14056 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 14464 11228 14516 11280
rect 15108 11228 15160 11280
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 11612 11092 11664 11144
rect 12256 11092 12308 11144
rect 12992 11160 13044 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 6460 11067 6512 11076
rect 6460 11033 6469 11067
rect 6469 11033 6503 11067
rect 6503 11033 6512 11067
rect 6460 11024 6512 11033
rect 2872 10999 2924 11008
rect 2872 10965 2881 10999
rect 2881 10965 2915 10999
rect 2915 10965 2924 10999
rect 2872 10956 2924 10965
rect 4896 10956 4948 11008
rect 7196 11024 7248 11076
rect 6920 10956 6972 11008
rect 12348 10956 12400 11008
rect 13728 11092 13780 11144
rect 15936 11135 15988 11144
rect 13452 11024 13504 11076
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1768 10752 1820 10804
rect 2688 10659 2740 10668
rect 2688 10625 2697 10659
rect 2697 10625 2731 10659
rect 2731 10625 2740 10659
rect 2688 10616 2740 10625
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 3884 10616 3936 10668
rect 4068 10616 4120 10668
rect 4712 10659 4764 10668
rect 4712 10625 4721 10659
rect 4721 10625 4755 10659
rect 4755 10625 4764 10659
rect 4712 10616 4764 10625
rect 2872 10548 2924 10600
rect 3516 10548 3568 10600
rect 7564 10752 7616 10804
rect 7840 10684 7892 10736
rect 8484 10727 8536 10736
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 8484 10693 8493 10727
rect 8493 10693 8527 10727
rect 8527 10693 8536 10727
rect 8484 10684 8536 10693
rect 8668 10752 8720 10804
rect 12992 10752 13044 10804
rect 14556 10795 14608 10804
rect 14556 10761 14565 10795
rect 14565 10761 14599 10795
rect 14599 10761 14608 10795
rect 14556 10752 14608 10761
rect 9680 10684 9732 10736
rect 11612 10684 11664 10736
rect 9588 10616 9640 10668
rect 9956 10616 10008 10668
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 17868 10616 17920 10668
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 11152 10548 11204 10600
rect 12256 10548 12308 10600
rect 15752 10591 15804 10600
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 18696 10548 18748 10600
rect 7104 10523 7156 10532
rect 7104 10489 7138 10523
rect 7138 10489 7156 10523
rect 7104 10480 7156 10489
rect 7196 10480 7248 10532
rect 8852 10523 8904 10532
rect 8852 10489 8861 10523
rect 8861 10489 8895 10523
rect 8895 10489 8904 10523
rect 8852 10480 8904 10489
rect 11704 10480 11756 10532
rect 13452 10523 13504 10532
rect 13452 10489 13486 10523
rect 13486 10489 13504 10523
rect 13452 10480 13504 10489
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 3516 10412 3568 10421
rect 3976 10412 4028 10464
rect 4896 10412 4948 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 8208 10412 8260 10464
rect 9312 10412 9364 10464
rect 9588 10412 9640 10464
rect 15660 10480 15712 10532
rect 16028 10523 16080 10532
rect 16028 10489 16062 10523
rect 16062 10489 16080 10523
rect 16028 10480 16080 10489
rect 14372 10412 14424 10464
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 3700 10208 3752 10260
rect 12348 10251 12400 10260
rect 3976 10140 4028 10192
rect 9680 10140 9732 10192
rect 11612 10140 11664 10192
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 4712 10072 4764 10124
rect 5816 10072 5868 10124
rect 1676 10004 1728 10056
rect 10416 10072 10468 10124
rect 12348 10217 12357 10251
rect 12357 10217 12391 10251
rect 12391 10217 12400 10251
rect 12348 10208 12400 10217
rect 12532 10208 12584 10260
rect 13452 10208 13504 10260
rect 17040 10208 17092 10260
rect 17132 10140 17184 10192
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 17868 10072 17920 10124
rect 12256 10004 12308 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 2688 9868 2740 9920
rect 4712 9868 4764 9920
rect 7104 9911 7156 9920
rect 7104 9877 7113 9911
rect 7113 9877 7147 9911
rect 7147 9877 7156 9911
rect 7104 9868 7156 9877
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 3516 9664 3568 9716
rect 8668 9664 8720 9716
rect 3240 9596 3292 9648
rect 4252 9596 4304 9648
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 7104 9528 7156 9580
rect 10416 9639 10468 9648
rect 10416 9605 10425 9639
rect 10425 9605 10459 9639
rect 10459 9605 10468 9639
rect 10416 9596 10468 9605
rect 14280 9596 14332 9648
rect 16764 9596 16816 9648
rect 10232 9528 10284 9580
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 4804 9460 4856 9512
rect 4988 9460 5040 9512
rect 8024 9460 8076 9512
rect 8208 9460 8260 9512
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 17040 9503 17092 9512
rect 14464 9460 14516 9469
rect 17040 9469 17049 9503
rect 17049 9469 17083 9503
rect 17083 9469 17092 9503
rect 17040 9460 17092 9469
rect 3240 9392 3292 9444
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4160 9324 4212 9376
rect 5540 9392 5592 9444
rect 6000 9392 6052 9444
rect 5724 9324 5776 9376
rect 7012 9392 7064 9444
rect 10968 9392 11020 9444
rect 17408 9392 17460 9444
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 7748 9324 7800 9376
rect 8944 9324 8996 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 1860 9120 1912 9172
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 5080 9120 5132 9172
rect 7196 9120 7248 9172
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 1860 8984 1912 9036
rect 3608 8984 3660 9036
rect 7748 8984 7800 9036
rect 8208 9120 8260 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 3516 8916 3568 8968
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 6368 8916 6420 8968
rect 8208 9027 8260 9036
rect 8208 8993 8242 9027
rect 8242 8993 8260 9027
rect 8208 8984 8260 8993
rect 8484 8984 8536 9036
rect 9404 8984 9456 9036
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 4712 8823 4764 8832
rect 4712 8789 4721 8823
rect 4721 8789 4755 8823
rect 4755 8789 4764 8823
rect 4712 8780 4764 8789
rect 9588 8780 9640 8832
rect 17960 8780 18012 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 4804 8576 4856 8628
rect 4528 8508 4580 8560
rect 5080 8508 5132 8560
rect 5816 8508 5868 8560
rect 6736 8508 6788 8560
rect 1860 8440 1912 8492
rect 4252 8440 4304 8492
rect 5264 8440 5316 8492
rect 8208 8508 8260 8560
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 1676 8304 1728 8356
rect 2688 8372 2740 8424
rect 4712 8372 4764 8424
rect 6368 8372 6420 8424
rect 8852 8372 8904 8424
rect 9956 8372 10008 8424
rect 2964 8304 3016 8356
rect 3700 8304 3752 8356
rect 3516 8279 3568 8288
rect 3516 8245 3525 8279
rect 3525 8245 3559 8279
rect 3559 8245 3568 8279
rect 3516 8236 3568 8245
rect 7748 8304 7800 8356
rect 5264 8236 5316 8288
rect 8484 8236 8536 8288
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 7748 8032 7800 8084
rect 8760 8032 8812 8084
rect 19524 8032 19576 8084
rect 1768 7964 1820 8016
rect 3884 7964 3936 8016
rect 4160 7896 4212 7948
rect 5356 7939 5408 7948
rect 5356 7905 5390 7939
rect 5390 7905 5408 7939
rect 5356 7896 5408 7905
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 8300 7896 8352 7948
rect 8852 7760 8904 7812
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 4252 7488 4304 7540
rect 2964 7395 3016 7404
rect 2964 7361 2973 7395
rect 2973 7361 3007 7395
rect 3007 7361 3016 7395
rect 2964 7352 3016 7361
rect 5356 7488 5408 7540
rect 19800 7488 19852 7540
rect 3516 7284 3568 7336
rect 4712 7284 4764 7336
rect 5080 7216 5132 7268
rect 5448 7216 5500 7268
rect 7748 7352 7800 7404
rect 8852 7352 8904 7404
rect 9312 7352 9364 7404
rect 3424 7148 3476 7200
rect 12348 7284 12400 7336
rect 7472 7148 7524 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 4988 6944 5040 6996
rect 5448 6944 5500 6996
rect 5540 6944 5592 6996
rect 5724 6876 5776 6928
rect 8760 6876 8812 6928
rect 12348 6876 12400 6928
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 8392 6808 8444 6860
rect 3884 6740 3936 6792
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 8116 6740 8168 6792
rect 8852 6783 8904 6792
rect 8852 6749 8861 6783
rect 8861 6749 8895 6783
rect 8895 6749 8904 6783
rect 8852 6740 8904 6749
rect 4160 6672 4212 6724
rect 8300 6672 8352 6724
rect 4804 6604 4856 6656
rect 7196 6604 7248 6656
rect 19616 6715 19668 6724
rect 19616 6681 19625 6715
rect 19625 6681 19659 6715
rect 19659 6681 19668 6715
rect 19616 6672 19668 6681
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 3884 6400 3936 6452
rect 7288 6400 7340 6452
rect 20720 6400 20772 6452
rect 4068 6196 4120 6248
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 21180 5856 21232 5908
rect 3976 5720 4028 5772
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2872 5312 2924 5364
rect 14096 5312 14148 5364
rect 20904 5312 20956 5364
rect 4068 5108 4120 5160
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3976 4088 4028 4140
rect 4988 4088 5040 4140
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 4068 1980 4120 2032
rect 5540 1980 5592 2032
rect 11428 1980 11480 2032
rect 11888 1980 11940 2032
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 1030 22320 1086 22800
rect 1490 22320 1546 22800
rect 1950 22320 2006 22800
rect 2134 22536 2190 22545
rect 2134 22471 2190 22480
rect 216 19242 244 22320
rect 204 19236 256 19242
rect 204 19178 256 19184
rect 584 18698 612 22320
rect 572 18692 624 18698
rect 572 18634 624 18640
rect 1044 18193 1072 22320
rect 1504 18986 1532 22320
rect 1582 20224 1638 20233
rect 1582 20159 1638 20168
rect 1412 18958 1532 18986
rect 1596 18970 1624 20159
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1780 19378 1808 19858
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1584 18964 1636 18970
rect 1412 18737 1440 18958
rect 1584 18906 1636 18912
rect 1492 18828 1544 18834
rect 1492 18770 1544 18776
rect 1398 18728 1454 18737
rect 1398 18663 1454 18672
rect 1030 18184 1086 18193
rect 1030 18119 1086 18128
rect 1504 17202 1532 18770
rect 1582 18320 1638 18329
rect 1582 18255 1638 18264
rect 1596 17882 1624 18255
rect 1688 18154 1716 19246
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1780 17921 1808 18022
rect 1766 17912 1822 17921
rect 1584 17876 1636 17882
rect 1766 17847 1822 17856
rect 1584 17818 1636 17824
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1412 16590 1440 17070
rect 1596 16658 1624 17614
rect 1674 16960 1730 16969
rect 1674 16895 1730 16904
rect 1688 16794 1716 16895
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1768 16040 1820 16046
rect 1674 16008 1730 16017
rect 1768 15982 1820 15988
rect 1674 15943 1730 15952
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 14550 1440 15506
rect 1688 14618 1716 15943
rect 1780 15638 1808 15982
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1400 14544 1452 14550
rect 1400 14486 1452 14492
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1596 13938 1624 14418
rect 1872 14226 1900 19751
rect 1964 19009 1992 22320
rect 1950 19000 2006 19009
rect 1950 18935 2006 18944
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 18426 1992 18770
rect 2148 18714 2176 22471
rect 2410 22320 2466 22800
rect 2870 22320 2926 22800
rect 3330 22320 3386 22800
rect 3790 22320 3846 22800
rect 4250 22320 4306 22800
rect 4710 22320 4766 22800
rect 5170 22320 5226 22800
rect 5630 22320 5686 22800
rect 6090 22320 6146 22800
rect 6550 22320 6606 22800
rect 7010 22320 7066 22800
rect 7470 22320 7526 22800
rect 7930 22320 7986 22800
rect 8390 22320 8446 22800
rect 8850 22320 8906 22800
rect 9310 22320 9366 22800
rect 9770 22320 9826 22800
rect 10230 22320 10286 22800
rect 10690 22320 10746 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12438 22320 12494 22800
rect 12898 22320 12954 22800
rect 13358 22320 13414 22800
rect 13818 22320 13874 22800
rect 14278 22320 14334 22800
rect 14738 22320 14794 22800
rect 15198 22320 15254 22800
rect 15658 22320 15714 22800
rect 16118 22320 16174 22800
rect 16578 22320 16634 22800
rect 17038 22320 17094 22800
rect 17498 22320 17554 22800
rect 17958 22320 18014 22800
rect 18418 22320 18474 22800
rect 18878 22320 18934 22800
rect 19338 22320 19394 22800
rect 19798 22320 19854 22800
rect 20258 22320 20314 22800
rect 20718 22320 20774 22800
rect 21178 22320 21234 22800
rect 21638 22320 21694 22800
rect 22098 22320 22154 22800
rect 22558 22320 22614 22800
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2240 19310 2268 19654
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2332 18902 2360 19858
rect 2424 19145 2452 22320
rect 2884 21706 2912 22320
rect 3146 22128 3202 22137
rect 3146 22063 3202 22072
rect 2884 21678 3096 21706
rect 2962 21584 3018 21593
rect 2962 21519 3018 21528
rect 2870 21176 2926 21185
rect 2870 21111 2926 21120
rect 2778 20632 2834 20641
rect 2778 20567 2834 20576
rect 2792 19786 2820 20567
rect 2884 20058 2912 21111
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2870 19272 2926 19281
rect 2870 19207 2926 19216
rect 2410 19136 2466 19145
rect 2410 19071 2466 19080
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2148 18686 2268 18714
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 2148 18222 2176 18566
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1964 16250 1992 16487
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2240 15722 2268 18686
rect 2686 17776 2742 17785
rect 2686 17711 2688 17720
rect 2740 17711 2742 17720
rect 2688 17682 2740 17688
rect 2148 15706 2268 15722
rect 2136 15700 2268 15706
rect 2188 15694 2268 15700
rect 2136 15642 2188 15648
rect 2792 15178 2820 18799
rect 2884 18170 2912 19207
rect 2976 19174 3004 21519
rect 3068 19514 3096 21678
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3054 19272 3110 19281
rect 3054 19207 3056 19216
rect 3108 19207 3110 19216
rect 3056 19178 3108 19184
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2884 18142 3096 18170
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 17377 2912 17478
rect 2870 17368 2926 17377
rect 2870 17303 2926 17312
rect 2976 17202 3004 18022
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2976 16250 3004 17138
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2870 15600 2926 15609
rect 2870 15535 2926 15544
rect 2700 15162 2820 15178
rect 2688 15156 2820 15162
rect 2740 15150 2820 15156
rect 2688 15098 2740 15104
rect 2502 14648 2558 14657
rect 2502 14583 2558 14592
rect 1780 14198 1900 14226
rect 1780 14074 1808 14198
rect 1858 14104 1914 14113
rect 1768 14068 1820 14074
rect 1858 14039 1914 14048
rect 1768 14010 1820 14016
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 13462 1440 13806
rect 1400 13456 1452 13462
rect 1400 13398 1452 13404
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1780 10810 1808 11630
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 8362 1716 9998
rect 1872 9178 1900 14039
rect 1950 13696 2006 13705
rect 1950 13631 2006 13640
rect 1964 12986 1992 13631
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 1964 11762 1992 12718
rect 2332 12374 2360 12718
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2516 9178 2544 14583
rect 2884 12986 2912 15535
rect 2976 15162 3004 16186
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2962 15056 3018 15065
rect 2962 14991 3018 15000
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2792 12306 2820 12854
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12374 2912 12718
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2976 11354 3004 14991
rect 3068 12986 3096 18142
rect 3160 17338 3188 22063
rect 3344 19258 3372 22320
rect 3344 19230 3648 19258
rect 3620 19174 3648 19230
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3252 17882 3280 18770
rect 3436 18086 3464 19110
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3528 18086 3556 18702
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3252 16776 3280 17274
rect 3160 16748 3280 16776
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 9926 2728 10610
rect 2884 10606 2912 10950
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1780 8022 1808 8978
rect 1872 8498 1900 8978
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 2700 8430 2728 9862
rect 3160 9489 3188 16748
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3252 15706 3280 16594
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3804 15434 3832 22320
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4080 18290 4108 19110
rect 4172 18766 4200 19110
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4172 18154 4200 18702
rect 4160 18148 4212 18154
rect 4160 18090 4212 18096
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4080 17134 4108 18022
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3792 15428 3844 15434
rect 3792 15370 3844 15376
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3344 13938 3372 14418
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 14074 3464 14350
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 9654 3280 11154
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3146 9480 3202 9489
rect 3146 9415 3202 9424
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 2976 7410 3004 8298
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2884 4321 2912 5306
rect 2870 4312 2926 4321
rect 2870 4247 2926 4256
rect 3252 1057 3280 9386
rect 3344 8129 3372 11562
rect 3528 10606 3556 15370
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3436 10266 3464 10406
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3528 9722 3556 10406
rect 3620 10033 3648 14214
rect 3698 12336 3754 12345
rect 3698 12271 3700 12280
rect 3752 12271 3754 12280
rect 3700 12242 3752 12248
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3712 10674 3740 11086
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3712 10266 3740 10610
rect 3804 10282 3832 15030
rect 3896 13734 3924 16730
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3988 15910 4016 16526
rect 4080 16182 4108 16934
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4172 16046 4200 16934
rect 4264 16794 4292 22320
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4264 16250 4292 16594
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4724 16114 4752 22320
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4908 19174 4936 19790
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 5000 18766 5028 19246
rect 5184 18970 5212 22320
rect 5644 20058 5672 22320
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5828 19242 5856 19790
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5908 18896 5960 18902
rect 5446 18864 5502 18873
rect 5908 18838 5960 18844
rect 5446 18799 5502 18808
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5000 17746 5028 18702
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5000 16590 5028 17682
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 16726 5212 17614
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 3988 14958 4016 15846
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 15162 4200 15438
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 3976 14952 4028 14958
rect 4172 14906 4200 15098
rect 3976 14894 4028 14900
rect 4080 14878 4200 14906
rect 4080 14414 4108 14878
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14550 4200 14758
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4172 13938 4200 14486
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4068 13320 4120 13326
rect 4066 13288 4068 13297
rect 4120 13288 4122 13297
rect 4066 13223 4122 13232
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3884 12776 3936 12782
rect 4080 12753 4108 13126
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3884 12718 3936 12724
rect 4066 12744 4122 12753
rect 3896 12238 3924 12718
rect 4066 12679 4122 12688
rect 4172 12374 4200 12786
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11898 3924 12174
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3896 10674 3924 11834
rect 3976 11824 4028 11830
rect 4080 11801 4108 12038
rect 4172 11898 4200 12310
rect 4264 11898 4292 12650
rect 4724 12306 4752 13670
rect 4908 12356 4936 15846
rect 5000 15638 5028 16526
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 5000 14362 5028 15574
rect 5080 14408 5132 14414
rect 5000 14356 5080 14362
rect 5000 14350 5132 14356
rect 5000 14334 5120 14350
rect 5000 13938 5028 14334
rect 5460 14226 5488 18799
rect 5920 18290 5948 18838
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5736 18170 5764 18226
rect 5736 18142 5856 18170
rect 5828 18086 5856 18142
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5736 17338 5764 18022
rect 5920 17882 5948 18226
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5828 16114 5856 16594
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5736 15162 5764 15846
rect 5828 15706 5856 16050
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5092 14198 5488 14226
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4988 13456 5040 13462
rect 4988 13398 5040 13404
rect 5000 12714 5028 13398
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 4816 12328 4936 12356
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 3976 11766 4028 11772
rect 4066 11792 4122 11801
rect 3988 11393 4016 11766
rect 4066 11727 4122 11736
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3988 10470 4016 11154
rect 4172 11150 4200 11698
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4540 11354 4568 11494
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3700 10260 3752 10266
rect 3804 10254 3924 10282
rect 3700 10202 3752 10208
rect 3606 10024 3662 10033
rect 3606 9959 3662 9968
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3330 8120 3386 8129
rect 3330 8055 3386 8064
rect 3436 7206 3464 9318
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3528 8294 3556 8910
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 7342 3556 8230
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3436 3913 3464 7142
rect 3422 3904 3478 3913
rect 3422 3839 3478 3848
rect 3238 1048 3294 1057
rect 3238 983 3294 992
rect 3620 649 3648 8978
rect 3896 8537 3924 10254
rect 3976 10192 4028 10198
rect 4080 10169 4108 10610
rect 3976 10134 4028 10140
rect 4066 10160 4122 10169
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3712 1601 3740 8298
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3896 7177 3924 7958
rect 3988 7585 4016 10134
rect 4066 10095 4068 10104
rect 4120 10095 4122 10104
rect 4068 10066 4120 10072
rect 4172 9382 4200 11086
rect 4264 9654 4292 11222
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4724 10130 4752 10610
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4724 9926 4752 10066
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4724 9586 4752 9862
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4816 9518 4844 12328
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10470 4936 10950
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3974 7576 4030 7585
rect 3974 7511 4030 7520
rect 3882 7168 3938 7177
rect 3882 7103 3938 7112
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 6458 3924 6734
rect 4172 6730 4200 7890
rect 4264 7546 4292 8434
rect 4540 8090 4568 8502
rect 4724 8430 4752 8774
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4724 6798 4752 7278
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4816 6662 4844 8570
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3896 3505 3924 6394
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4080 5817 4108 6190
rect 4066 5808 4122 5817
rect 3976 5772 4028 5778
rect 4066 5743 4122 5752
rect 3976 5714 4028 5720
rect 3988 5273 4016 5714
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 3974 5264 4030 5273
rect 3974 5199 4030 5208
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4865 4108 5102
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3882 3496 3938 3505
rect 3882 3431 3938 3440
rect 3988 2961 4016 4082
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 3974 2952 4030 2961
rect 4908 2938 4936 10406
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5000 7002 5028 9454
rect 5092 9178 5120 14198
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13326 5488 13738
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12986 5488 13262
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5368 12442 5396 12650
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 5092 7886 5120 8502
rect 5276 8498 5304 8910
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5092 7274 5120 7822
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5000 4146 5028 6938
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 3974 2887 4030 2896
rect 4724 2910 4936 2938
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4068 2032 4120 2038
rect 4066 2000 4068 2009
rect 4120 2000 4122 2009
rect 4066 1935 4122 1944
rect 3698 1592 3754 1601
rect 3698 1527 3754 1536
rect 3606 640 3662 649
rect 3606 575 3662 584
rect 4724 241 4752 2910
rect 5276 2553 5304 8230
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5368 7546 5396 7890
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 7002 5488 7210
rect 5552 7002 5580 9386
rect 5736 9382 5764 14758
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5828 10470 5856 12242
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10169 5856 10406
rect 5814 10160 5870 10169
rect 5814 10095 5816 10104
rect 5868 10095 5870 10104
rect 5816 10066 5868 10072
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5262 2544 5318 2553
rect 5262 2479 5318 2488
rect 5552 2038 5580 6938
rect 5736 6934 5764 9318
rect 5828 8566 5856 10066
rect 6012 9450 6040 19858
rect 6104 17202 6132 22320
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6196 17202 6224 17682
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6196 16794 6224 17138
rect 6380 17134 6408 17614
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6196 15026 6224 15506
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6196 14074 6224 14962
rect 6288 14278 6316 14962
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6288 12850 6316 13330
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6380 8974 6408 17070
rect 6564 14958 6592 22320
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6840 18970 6868 19178
rect 6918 19000 6974 19009
rect 6828 18964 6880 18970
rect 6918 18935 6920 18944
rect 6828 18906 6880 18912
rect 6972 18935 6974 18944
rect 6920 18906 6972 18912
rect 7024 18034 7052 22320
rect 7102 19136 7158 19145
rect 7102 19071 7158 19080
rect 7116 18902 7144 19071
rect 7104 18896 7156 18902
rect 7104 18838 7156 18844
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18222 7144 18566
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 6840 18006 7052 18034
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 6472 14074 6500 14826
rect 6656 14822 6684 15302
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6748 14482 6776 14894
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6564 13870 6592 14214
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6564 12374 6592 13806
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6472 11082 6500 12242
rect 6748 11540 6776 13874
rect 6840 13530 6868 18006
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7024 15706 7052 17682
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 7116 16590 7144 17002
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7208 15638 7236 16594
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15706 7328 15846
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7484 14634 7512 22320
rect 7944 20346 7972 22320
rect 7944 20318 8248 20346
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 8220 19258 8248 20318
rect 7668 17066 7696 19246
rect 8220 19230 8340 19258
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8220 18766 8248 19110
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 7760 18222 7788 18702
rect 8128 18426 8156 18702
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7760 16114 7788 18022
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17134 8248 18702
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8220 16658 8248 16934
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8128 15994 8156 16526
rect 8220 16114 8248 16594
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8128 15966 8248 15994
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15706 8248 15966
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7944 14906 7972 15506
rect 7024 14606 7512 14634
rect 7760 14878 7972 14906
rect 7564 14612 7616 14618
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6932 13530 6960 13942
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 11898 6868 12582
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 7024 11694 7052 14606
rect 7564 14554 7616 14560
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7208 13802 7236 14486
rect 7300 14074 7328 14486
rect 7576 14074 7604 14554
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 13190 7328 13738
rect 7760 13190 7788 14878
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14482 8248 14758
rect 8312 14618 8340 19230
rect 8404 18086 8432 22320
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8496 17785 8524 18702
rect 8772 18630 8800 19178
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8772 18290 8800 18566
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8864 18222 8892 22320
rect 9324 20058 9352 22320
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9692 19310 9720 19858
rect 9784 19802 9812 22320
rect 10048 19848 10100 19854
rect 9784 19774 9904 19802
rect 10100 19796 10180 19802
rect 10048 19790 10180 19796
rect 10060 19774 10180 19790
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9784 18834 9812 19654
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8852 18216 8904 18222
rect 8956 18193 8984 18226
rect 8852 18158 8904 18164
rect 8942 18184 8998 18193
rect 8942 18119 8998 18128
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 8482 17776 8538 17785
rect 8482 17711 8538 17720
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8772 16454 8800 17070
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8404 15026 8432 15982
rect 8496 15502 8524 16390
rect 8772 16046 8800 16390
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8312 14006 8340 14214
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8404 13938 8432 14962
rect 8496 14958 8524 15438
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8956 14890 8984 18022
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8588 14278 8616 14826
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8864 13326 8892 13738
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12850 7788 13126
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11762 7144 12038
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7196 11552 7248 11558
rect 6748 11512 7052 11540
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6828 10668 6880 10674
rect 6932 10656 6960 10950
rect 6880 10628 6960 10656
rect 6828 10610 6880 10616
rect 7024 9450 7052 11512
rect 7196 11494 7248 11500
rect 7208 11082 7236 11494
rect 7484 11150 7512 11834
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7208 10538 7236 11018
rect 7576 10810 7604 12582
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8220 11898 8248 12718
rect 8680 12442 8708 13262
rect 8864 12986 8892 13262
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8956 12306 8984 13398
rect 9048 12442 9076 18022
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 11098 7788 11154
rect 7760 11070 7880 11098
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7852 10742 7880 11070
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7116 9926 7144 10474
rect 8220 10470 8248 11834
rect 8496 10742 8524 12242
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8864 11626 8892 12174
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11354 8892 11562
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8484 10736 8536 10742
rect 8680 10713 8708 10746
rect 8484 10678 8536 10684
rect 8666 10704 8722 10713
rect 8666 10639 8722 10648
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7116 9586 7144 9862
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 8036 9518 8064 9862
rect 8220 9518 8248 10406
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8680 9722 8708 9998
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7208 9178 7236 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 6380 8430 6408 8910
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6748 7886 6776 8502
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6225 7236 6598
rect 7300 6458 7328 9318
rect 7760 9042 7788 9318
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8220 9178 8248 9454
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8220 8566 8248 8978
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7760 8090 7788 8298
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7760 7410 7788 8026
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 6866 7512 7142
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8220 6882 8248 8502
rect 8496 8294 8524 8978
rect 8864 8430 8892 10474
rect 8956 9382 8984 12242
rect 9140 12238 9168 12650
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11898 9168 12174
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9048 11354 9076 11630
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9310 10704 9366 10713
rect 9310 10639 9366 10648
rect 9324 10470 9352 10639
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9416 9042 9444 18090
rect 9692 17814 9720 18634
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9784 17134 9812 18158
rect 9876 17882 9904 19774
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9968 18766 9996 19246
rect 10152 19242 10180 19774
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 10046 19000 10102 19009
rect 10046 18935 10102 18944
rect 10060 18902 10088 18935
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9968 18154 9996 18702
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9772 17128 9824 17134
rect 10060 17082 10088 18838
rect 10152 18426 10180 19178
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10244 18306 10272 22320
rect 10414 19272 10470 19281
rect 10414 19207 10470 19216
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10336 18834 10364 19110
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10244 18278 10364 18306
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 9772 17070 9824 17076
rect 9968 17054 10088 17082
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 14618 9720 15506
rect 9784 15502 9812 15914
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9784 15162 9812 15438
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9968 15026 9996 17054
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16794 10088 16934
rect 10152 16794 10180 17478
rect 10244 16998 10272 18090
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10244 16590 10272 16934
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10336 15706 10364 18278
rect 10428 18154 10456 19207
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10704 18086 10732 22320
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10980 19174 11008 19790
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10428 17066 10456 17614
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10428 16250 10456 17002
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 10244 14958 10272 15438
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9784 14074 9812 14894
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13394 10272 13670
rect 10796 13394 10824 16118
rect 10888 15570 10916 16526
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 11762 9720 12242
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 10796 11694 10824 12174
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 9680 10736 9732 10742
rect 9586 10704 9642 10713
rect 9680 10678 9732 10684
rect 9586 10639 9588 10648
rect 9640 10639 9642 10648
rect 9588 10610 9640 10616
rect 9692 10606 9720 10678
rect 9968 10674 9996 11630
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9680 10600 9732 10606
rect 9586 10568 9642 10577
rect 9680 10542 9732 10548
rect 9586 10503 9642 10512
rect 9600 10470 9628 10503
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9692 9178 9720 10134
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10428 9654 10456 10066
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 9954 9480 10010 9489
rect 9954 9415 10010 9424
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9588 8832 9640 8838
rect 9586 8800 9588 8809
rect 9640 8800 9642 8809
rect 9586 8735 9642 8744
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 8090 8800 8230
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 8128 6854 8248 6882
rect 8128 6798 8156 6854
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8312 6730 8340 7890
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 6866 8432 7686
rect 8864 7410 8892 7754
rect 9324 7410 9352 8434
rect 9968 8430 9996 9415
rect 10244 8974 10272 9522
rect 10980 9450 11008 18022
rect 11072 17270 11100 18906
rect 11164 17320 11192 22320
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11624 18086 11652 22320
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11716 18873 11744 18906
rect 11702 18864 11758 18873
rect 11702 18799 11758 18808
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11164 17292 11744 17320
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12714 11100 13262
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 11164 11642 11192 14554
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11624 13870 11652 14758
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11624 13190 11652 13398
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11440 12238 11468 12718
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11440 12084 11468 12174
rect 11440 12056 11652 12084
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11072 11614 11192 11642
rect 11624 11626 11652 12056
rect 11612 11620 11664 11626
rect 11072 9761 11100 11614
rect 11612 11562 11664 11568
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 10606 11192 11494
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 10742 11652 11086
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11624 10198 11652 10678
rect 11716 10538 11744 17292
rect 11900 15978 11928 18158
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11900 15026 11928 15302
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14550 11928 14962
rect 11992 14618 12020 22320
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 12084 15706 12112 19178
rect 12452 18970 12480 22320
rect 12912 20058 12940 22320
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11808 13326 11836 13874
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11058 9752 11114 9761
rect 11252 9744 11548 9764
rect 11058 9687 11114 9696
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8772 6769 8800 6870
rect 8864 6798 8892 7346
rect 8852 6792 8904 6798
rect 8758 6760 8814 6769
rect 8300 6724 8352 6730
rect 8852 6734 8904 6740
rect 8758 6695 8814 6704
rect 8300 6666 8352 6672
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7194 6216 7250 6225
rect 7194 6151 7250 6160
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11900 2038 11928 14010
rect 11992 13938 12020 14214
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12176 13870 12204 18090
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12268 16454 12296 17138
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12268 15638 12296 16390
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 12360 15570 12388 15846
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12360 14482 12388 15506
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12268 13734 12296 14214
rect 12346 14104 12402 14113
rect 12346 14039 12402 14048
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 12646 12020 13262
rect 12084 13190 12112 13466
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11992 12374 12020 12582
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11992 11354 12020 11630
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 12176 10962 12204 11494
rect 12360 11370 12388 14039
rect 12452 13530 12480 18770
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12544 17082 12572 17614
rect 12636 17338 12664 19246
rect 13096 18970 13124 19858
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13280 18902 13308 19722
rect 13372 19394 13400 22320
rect 13832 20074 13860 22320
rect 13832 20046 13952 20074
rect 14292 20058 14320 22320
rect 14752 20482 14780 22320
rect 15212 20618 15240 22320
rect 15212 20590 15332 20618
rect 14752 20454 15240 20482
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13372 19366 13492 19394
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13268 18896 13320 18902
rect 13268 18838 13320 18844
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12544 17054 12664 17082
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16794 12572 16934
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12452 12850 12480 13330
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12544 11762 12572 13670
rect 12636 13258 12664 17054
rect 12728 14482 12756 17750
rect 12820 16182 12848 18634
rect 12912 17882 12940 18770
rect 13266 18728 13322 18737
rect 13266 18663 13322 18672
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 13096 17678 13124 18090
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16794 12940 16934
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12912 16114 12940 16594
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 13004 15706 13032 16526
rect 13096 16250 13124 17614
rect 13188 17202 13216 17682
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12728 14113 12756 14418
rect 12714 14104 12770 14113
rect 12714 14039 12770 14048
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12728 13530 12756 13942
rect 12820 13802 12848 15506
rect 12900 15088 12952 15094
rect 12898 15056 12900 15065
rect 12952 15056 12954 15065
rect 12898 14991 12954 15000
rect 13280 14618 13308 18663
rect 13372 15162 13400 19246
rect 13464 19174 13492 19366
rect 13832 19310 13860 19858
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13924 19242 13952 20046
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14108 19310 14136 19790
rect 15212 19786 15240 20454
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13464 18426 13492 18838
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13464 17542 13492 18226
rect 13740 18086 13768 18702
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13740 17814 13768 18022
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 15706 13952 16594
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 14016 16250 14044 16526
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 13096 12306 13124 13874
rect 13464 13802 13492 15438
rect 13556 14074 13584 15506
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13452 13796 13504 13802
rect 13452 13738 13504 13744
rect 13464 12646 13492 13738
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13556 12374 13584 14010
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13740 13190 13768 13806
rect 13832 13530 13860 14758
rect 14016 13870 14044 15846
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13530 13952 13670
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12636 11626 12664 12038
rect 12728 11830 12756 12038
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12360 11342 12572 11370
rect 13188 11354 13216 11494
rect 12256 11144 12308 11150
rect 12360 11132 12388 11342
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12308 11104 12388 11132
rect 12256 11086 12308 11092
rect 12348 11008 12400 11014
rect 12176 10934 12296 10962
rect 12348 10950 12400 10956
rect 12268 10606 12296 10934
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12268 10062 12296 10542
rect 12360 10266 12388 10950
rect 12452 10674 12480 11222
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12544 10266 12572 11342
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 13004 10810 13032 11154
rect 13728 11144 13780 11150
rect 13832 11098 13860 13330
rect 14016 11354 14044 13806
rect 14108 13394 14136 18770
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14200 13462 14228 14758
rect 14384 14260 14412 19246
rect 15304 19174 15332 20590
rect 15672 20058 15700 22320
rect 16132 20618 16160 22320
rect 16132 20590 16344 20618
rect 16316 20058 16344 20590
rect 16592 20074 16620 22320
rect 16592 20058 16896 20074
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 16304 20052 16356 20058
rect 16592 20052 16908 20058
rect 16592 20046 16856 20052
rect 16304 19994 16356 20000
rect 16856 19994 16908 20000
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14462 19000 14518 19009
rect 14684 18992 14980 19012
rect 14462 18935 14464 18944
rect 14516 18935 14518 18944
rect 14464 18906 14516 18912
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14660 18222 14688 18566
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 15304 17882 15332 18022
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14476 15706 14504 17206
rect 14568 16046 14596 17478
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 16182 14780 16526
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14476 14890 14504 15642
rect 14568 15502 14596 15982
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14292 14232 14412 14260
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 12442 14228 12582
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13780 11092 13860 11098
rect 13728 11086 13860 11092
rect 13452 11076 13504 11082
rect 13740 11070 13860 11086
rect 13452 11018 13504 11024
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13464 10538 13492 11018
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13464 10266 13492 10474
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12360 6934 12388 7278
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 14108 5370 14136 12242
rect 14292 9654 14320 14232
rect 14476 13410 14504 14418
rect 14568 13938 14596 14962
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14384 13382 14504 13410
rect 14384 13326 14412 13382
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14384 12986 14412 13262
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14384 12238 14412 12786
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14476 12170 14504 13262
rect 14568 12850 14596 13874
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15028 13530 15056 14894
rect 15120 14822 15148 15574
rect 15212 15094 15240 16594
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 15706 15332 15914
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15212 14618 15240 15030
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15108 14544 15160 14550
rect 15396 14498 15424 19858
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 16454 15516 18022
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16250 15516 16390
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15488 15502 15516 16186
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 15094 15516 15438
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 15108 14486 15160 14492
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14844 12850 14872 13330
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14752 11694 14780 12174
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14384 9518 14412 10406
rect 14476 9518 14504 11222
rect 14568 10810 14596 11562
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15120 11286 15148 14486
rect 15212 14470 15424 14498
rect 15212 11898 15240 14470
rect 15488 13938 15516 15030
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15580 12442 15608 19246
rect 15672 19242 15700 19858
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15658 18728 15714 18737
rect 15658 18663 15714 18672
rect 15672 17882 15700 18663
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 13802 15700 15846
rect 15764 15162 15792 18770
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15948 18154 15976 18702
rect 15936 18148 15988 18154
rect 15936 18090 15988 18096
rect 15948 17678 15976 18090
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15948 16794 15976 17614
rect 16040 17202 16068 18906
rect 16316 18902 16344 19246
rect 16592 19242 16620 19858
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16684 18902 16712 19858
rect 17052 19786 17080 22320
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 17512 19258 17540 22320
rect 17972 19394 18000 22320
rect 18432 20058 18460 22320
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17880 19366 18000 19394
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16316 16114 16344 16594
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16592 15162 16620 18770
rect 16672 15632 16724 15638
rect 16672 15574 16724 15580
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 15764 14482 15792 15098
rect 16210 15056 16266 15065
rect 16684 15042 16712 15574
rect 16592 15026 16712 15042
rect 16210 14991 16266 15000
rect 16580 15020 16712 15026
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15948 14278 15976 14758
rect 16224 14550 16252 14991
rect 16632 15014 16712 15020
rect 16580 14962 16632 14968
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 13870 16344 14214
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16224 12714 16252 13738
rect 16592 12986 16620 14962
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 16132 12238 16160 12650
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15304 11354 15332 12174
rect 16132 11898 16160 12174
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14568 9586 14596 10746
rect 15672 10538 15700 11154
rect 15764 10606 15792 11630
rect 15936 11620 15988 11626
rect 15936 11562 15988 11568
rect 15948 11150 15976 11562
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 16040 10062 16068 10474
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16776 9654 16804 18770
rect 16868 14346 16896 19246
rect 17408 19236 17460 19242
rect 17512 19230 17632 19258
rect 17408 19178 17460 19184
rect 17420 18222 17448 19178
rect 17604 19174 17632 19230
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17880 18426 17908 19366
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16960 17338 16988 17614
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17604 16250 17632 17138
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16658 17908 17070
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17972 16250 18000 19246
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18524 18290 18552 19858
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18616 18902 18644 19790
rect 18892 19242 18920 22320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18984 18970 19012 19246
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18616 17882 18644 18702
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17144 15706 17172 15914
rect 17972 15706 18000 15914
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18432 15706 18460 15846
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 17144 15026 17172 15642
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17420 14958 17448 15438
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 17420 14074 17448 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17420 13462 17448 14010
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16960 12782 16988 13330
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16960 12442 16988 12718
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17880 11830 17908 12310
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17880 10674 17908 11766
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 17052 9518 17080 10202
rect 17144 10198 17172 10406
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17144 9586 17172 10134
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17420 9450 17448 10406
rect 17880 10130 17908 10610
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 17972 8838 18000 15506
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18340 14482 18368 14962
rect 18616 14958 18644 15438
rect 18708 15162 18736 16050
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18708 14550 18736 15098
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18616 12850 18644 13126
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18616 12306 18644 12786
rect 18984 12442 19012 18158
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19260 15502 19288 16390
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19352 13818 19380 22320
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19444 16998 19472 17614
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19444 16726 19472 16934
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19352 13790 19564 13818
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19444 12442 19472 12854
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18616 11762 18644 12242
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18708 10606 18736 12038
rect 19352 11898 19380 12242
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 19536 8090 19564 13790
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 19628 6730 19656 18022
rect 19720 12782 19748 18090
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19812 7546 19840 22320
rect 20272 18086 20300 22320
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20364 18698 20392 19314
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19996 11529 20024 11562
rect 19982 11520 20038 11529
rect 19982 11455 20038 11464
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 20732 6458 20760 22320
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 20916 5370 20944 18022
rect 21192 5914 21220 22320
rect 21652 18086 21680 22320
rect 22112 19310 22140 22320
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22572 18154 22600 22320
rect 22560 18148 22612 18154
rect 22560 18090 22612 18096
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 11888 2032 11940 2038
rect 11888 1974 11940 1980
rect 11440 480 11468 1974
rect 4710 232 4766 241
rect 4710 167 4766 176
rect 11426 0 11482 480
<< via2 >>
rect 2134 22480 2190 22536
rect 1582 20168 1638 20224
rect 1858 19760 1914 19816
rect 1398 18672 1454 18728
rect 1030 18128 1086 18184
rect 1582 18264 1638 18320
rect 1766 17856 1822 17912
rect 1674 16904 1730 16960
rect 1674 15952 1730 16008
rect 1950 18944 2006 19000
rect 3146 22072 3202 22128
rect 2962 21528 3018 21584
rect 2870 21120 2926 21176
rect 2778 20576 2834 20632
rect 2870 19216 2926 19272
rect 2410 19080 2466 19136
rect 2778 18808 2834 18864
rect 1950 16496 2006 16552
rect 2686 17740 2742 17776
rect 2686 17720 2688 17740
rect 2688 17720 2740 17740
rect 2740 17720 2742 17740
rect 3054 19236 3110 19272
rect 3054 19216 3056 19236
rect 3056 19216 3108 19236
rect 3108 19216 3110 19236
rect 2870 17312 2926 17368
rect 2870 15544 2926 15600
rect 2502 14592 2558 14648
rect 1858 14048 1914 14104
rect 1950 13640 2006 13696
rect 2962 15000 3018 15056
rect 3146 9424 3202 9480
rect 2870 4256 2926 4312
rect 3698 12300 3754 12336
rect 3698 12280 3700 12300
rect 3700 12280 3752 12300
rect 3752 12280 3754 12300
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 5446 18808 5502 18864
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4066 13268 4068 13288
rect 4068 13268 4120 13288
rect 4120 13268 4122 13288
rect 4066 13232 4122 13268
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4066 12688 4122 12744
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 11736 4122 11792
rect 3974 11328 4030 11384
rect 3606 9968 3662 10024
rect 3330 8064 3386 8120
rect 3422 3848 3478 3904
rect 3238 992 3294 1048
rect 3882 8472 3938 8528
rect 4066 10124 4122 10160
rect 4066 10104 4068 10124
rect 4068 10104 4120 10124
rect 4120 10104 4122 10124
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 3974 7520 4030 7576
rect 3882 7112 3938 7168
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4066 5752 4122 5808
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 3974 5208 4030 5264
rect 4066 4800 4122 4856
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 3882 3440 3938 3496
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 3974 2896 4030 2952
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4066 1980 4068 2000
rect 4068 1980 4120 2000
rect 4120 1980 4122 2000
rect 4066 1944 4122 1980
rect 3698 1536 3754 1592
rect 3606 584 3662 640
rect 5814 10124 5870 10160
rect 5814 10104 5816 10124
rect 5816 10104 5868 10124
rect 5868 10104 5870 10124
rect 5262 2488 5318 2544
rect 6918 18964 6974 19000
rect 6918 18944 6920 18964
rect 6920 18944 6972 18964
rect 6972 18944 6974 18964
rect 7102 19080 7158 19136
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 8942 18128 8998 18184
rect 8482 17720 8538 17776
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8666 10648 8722 10704
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 9310 10648 9366 10704
rect 10046 18944 10102 19000
rect 10414 19216 10470 19272
rect 9586 10668 9642 10704
rect 9586 10648 9588 10668
rect 9588 10648 9640 10668
rect 9640 10648 9642 10668
rect 9586 10512 9642 10568
rect 9954 9424 10010 9480
rect 9586 8780 9588 8800
rect 9588 8780 9640 8800
rect 9640 8780 9642 8800
rect 9586 8744 9642 8780
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11702 18808 11758 18864
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11058 9696 11114 9752
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 8758 6704 8814 6760
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 7194 6160 7250 6216
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12346 14048 12402 14104
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 13266 18672 13322 18728
rect 12714 14048 12770 14104
rect 12898 15036 12900 15056
rect 12900 15036 12952 15056
rect 12952 15036 12954 15056
rect 12898 15000 12954 15036
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14462 18964 14518 19000
rect 14462 18944 14464 18964
rect 14464 18944 14516 18964
rect 14516 18944 14518 18964
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 15658 18672 15714 18728
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 16210 15000 16266 15056
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 19982 11464 20038 11520
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 4710 176 4766 232
<< metal3 >>
rect 0 22538 480 22568
rect 2129 22538 2195 22541
rect 0 22536 2195 22538
rect 0 22480 2134 22536
rect 2190 22480 2195 22536
rect 0 22478 2195 22480
rect 0 22448 480 22478
rect 2129 22475 2195 22478
rect 0 22130 480 22160
rect 3141 22130 3207 22133
rect 0 22128 3207 22130
rect 0 22072 3146 22128
rect 3202 22072 3207 22128
rect 0 22070 3207 22072
rect 0 22040 480 22070
rect 3141 22067 3207 22070
rect 0 21586 480 21616
rect 2957 21586 3023 21589
rect 0 21584 3023 21586
rect 0 21528 2962 21584
rect 3018 21528 3023 21584
rect 0 21526 3023 21528
rect 0 21496 480 21526
rect 2957 21523 3023 21526
rect 0 21178 480 21208
rect 2865 21178 2931 21181
rect 0 21176 2931 21178
rect 0 21120 2870 21176
rect 2926 21120 2931 21176
rect 0 21118 2931 21120
rect 0 21088 480 21118
rect 2865 21115 2931 21118
rect 0 20634 480 20664
rect 2773 20634 2839 20637
rect 0 20632 2839 20634
rect 0 20576 2778 20632
rect 2834 20576 2839 20632
rect 0 20574 2839 20576
rect 0 20544 480 20574
rect 2773 20571 2839 20574
rect 0 20226 480 20256
rect 1577 20226 1643 20229
rect 0 20224 1643 20226
rect 0 20168 1582 20224
rect 1638 20168 1643 20224
rect 0 20166 1643 20168
rect 0 20136 480 20166
rect 1577 20163 1643 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 480 19758
rect 1853 19755 1919 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 2865 19274 2931 19277
rect 0 19272 2931 19274
rect 0 19216 2870 19272
rect 2926 19216 2931 19272
rect 0 19214 2931 19216
rect 0 19184 480 19214
rect 2865 19211 2931 19214
rect 3049 19274 3115 19277
rect 10409 19274 10475 19277
rect 3049 19272 10475 19274
rect 3049 19216 3054 19272
rect 3110 19216 10414 19272
rect 10470 19216 10475 19272
rect 3049 19214 10475 19216
rect 3049 19211 3115 19214
rect 10409 19211 10475 19214
rect 2405 19138 2471 19141
rect 7097 19138 7163 19141
rect 2405 19136 7163 19138
rect 2405 19080 2410 19136
rect 2466 19080 7102 19136
rect 7158 19080 7163 19136
rect 2405 19078 7163 19080
rect 2405 19075 2471 19078
rect 7097 19075 7163 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 1945 19002 2011 19005
rect 6913 19002 6979 19005
rect 1945 19000 6979 19002
rect 1945 18944 1950 19000
rect 2006 18944 6918 19000
rect 6974 18944 6979 19000
rect 1945 18942 6979 18944
rect 1945 18939 2011 18942
rect 6913 18939 6979 18942
rect 10041 19002 10107 19005
rect 14457 19002 14523 19005
rect 10041 19000 14523 19002
rect 10041 18944 10046 19000
rect 10102 18944 14462 19000
rect 14518 18944 14523 19000
rect 10041 18942 14523 18944
rect 10041 18939 10107 18942
rect 14457 18939 14523 18942
rect 0 18866 480 18896
rect 2773 18866 2839 18869
rect 0 18864 2839 18866
rect 0 18808 2778 18864
rect 2834 18808 2839 18864
rect 0 18806 2839 18808
rect 0 18776 480 18806
rect 2773 18803 2839 18806
rect 5441 18866 5507 18869
rect 11697 18866 11763 18869
rect 5441 18864 11763 18866
rect 5441 18808 5446 18864
rect 5502 18808 11702 18864
rect 11758 18808 11763 18864
rect 5441 18806 11763 18808
rect 5441 18803 5507 18806
rect 11697 18803 11763 18806
rect 1393 18730 1459 18733
rect 13261 18730 13327 18733
rect 15653 18730 15719 18733
rect 1393 18728 15719 18730
rect 1393 18672 1398 18728
rect 1454 18672 13266 18728
rect 13322 18672 15658 18728
rect 15714 18672 15719 18728
rect 1393 18670 15719 18672
rect 1393 18667 1459 18670
rect 13261 18667 13327 18670
rect 15653 18667 15719 18670
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1577 18322 1643 18325
rect 0 18320 1643 18322
rect 0 18264 1582 18320
rect 1638 18264 1643 18320
rect 0 18262 1643 18264
rect 0 18232 480 18262
rect 1577 18259 1643 18262
rect 1025 18186 1091 18189
rect 8937 18186 9003 18189
rect 1025 18184 9003 18186
rect 1025 18128 1030 18184
rect 1086 18128 8942 18184
rect 8998 18128 9003 18184
rect 1025 18126 9003 18128
rect 1025 18123 1091 18126
rect 8937 18123 9003 18126
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1761 17914 1827 17917
rect 0 17912 1827 17914
rect 0 17856 1766 17912
rect 1822 17856 1827 17912
rect 0 17854 1827 17856
rect 0 17824 480 17854
rect 1761 17851 1827 17854
rect 2681 17778 2747 17781
rect 8477 17778 8543 17781
rect 2681 17776 8543 17778
rect 2681 17720 2686 17776
rect 2742 17720 8482 17776
rect 8538 17720 8543 17776
rect 2681 17718 8543 17720
rect 2681 17715 2747 17718
rect 8477 17715 8543 17718
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 2865 17370 2931 17373
rect 0 17368 2931 17370
rect 0 17312 2870 17368
rect 2926 17312 2931 17368
rect 0 17310 2931 17312
rect 0 17280 480 17310
rect 2865 17307 2931 17310
rect 0 16962 480 16992
rect 1669 16962 1735 16965
rect 0 16960 1735 16962
rect 0 16904 1674 16960
rect 1730 16904 1735 16960
rect 0 16902 1735 16904
rect 0 16872 480 16902
rect 1669 16899 1735 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 480 16494
rect 1945 16491 2011 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1669 16010 1735 16013
rect 0 16008 1735 16010
rect 0 15952 1674 16008
rect 1730 15952 1735 16008
rect 0 15950 1735 15952
rect 0 15920 480 15950
rect 1669 15947 1735 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 2865 15602 2931 15605
rect 0 15600 2931 15602
rect 0 15544 2870 15600
rect 2926 15544 2931 15600
rect 0 15542 2931 15544
rect 0 15512 480 15542
rect 2865 15539 2931 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 2957 15058 3023 15061
rect 0 15056 3023 15058
rect 0 15000 2962 15056
rect 3018 15000 3023 15056
rect 0 14998 3023 15000
rect 0 14968 480 14998
rect 2957 14995 3023 14998
rect 12893 15058 12959 15061
rect 16205 15058 16271 15061
rect 12893 15056 16271 15058
rect 12893 15000 12898 15056
rect 12954 15000 16210 15056
rect 16266 15000 16271 15056
rect 12893 14998 16271 15000
rect 12893 14995 12959 14998
rect 16205 14995 16271 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 2497 14650 2563 14653
rect 0 14648 2563 14650
rect 0 14592 2502 14648
rect 2558 14592 2563 14648
rect 0 14590 2563 14592
rect 0 14560 480 14590
rect 2497 14587 2563 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1853 14106 1919 14109
rect 0 14104 1919 14106
rect 0 14048 1858 14104
rect 1914 14048 1919 14104
rect 0 14046 1919 14048
rect 0 14016 480 14046
rect 1853 14043 1919 14046
rect 12341 14106 12407 14109
rect 12709 14106 12775 14109
rect 12341 14104 12775 14106
rect 12341 14048 12346 14104
rect 12402 14048 12714 14104
rect 12770 14048 12775 14104
rect 12341 14046 12775 14048
rect 12341 14043 12407 14046
rect 12709 14043 12775 14046
rect 0 13698 480 13728
rect 1945 13698 2011 13701
rect 0 13696 2011 13698
rect 0 13640 1950 13696
rect 2006 13640 2011 13696
rect 0 13638 2011 13640
rect 0 13608 480 13638
rect 1945 13635 2011 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 4061 13290 4127 13293
rect 0 13288 4127 13290
rect 0 13232 4066 13288
rect 4122 13232 4127 13288
rect 0 13230 4127 13232
rect 0 13200 480 13230
rect 4061 13227 4127 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 480 12686
rect 4061 12683 4127 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 3693 12338 3759 12341
rect 0 12336 3759 12338
rect 0 12280 3698 12336
rect 3754 12280 3759 12336
rect 0 12278 3759 12280
rect 0 12248 480 12278
rect 3693 12275 3759 12278
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 480 11734
rect 4061 11731 4127 11734
rect 19977 11522 20043 11525
rect 22320 11522 22800 11552
rect 19977 11520 22800 11522
rect 19977 11464 19982 11520
rect 20038 11464 22800 11520
rect 19977 11462 22800 11464
rect 19977 11459 20043 11462
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 22320 11432 22800 11462
rect 14672 11391 14992 11392
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 480 11326
rect 3969 11323 4035 11326
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 0 10782 4170 10842
rect 0 10752 480 10782
rect 4110 10706 4170 10782
rect 8661 10706 8727 10709
rect 4110 10704 8727 10706
rect 4110 10648 8666 10704
rect 8722 10648 8727 10704
rect 4110 10646 8727 10648
rect 8661 10643 8727 10646
rect 9305 10706 9371 10709
rect 9581 10706 9647 10709
rect 9305 10704 9647 10706
rect 9305 10648 9310 10704
rect 9366 10648 9586 10704
rect 9642 10648 9647 10704
rect 9305 10646 9647 10648
rect 9305 10643 9371 10646
rect 9581 10643 9647 10646
rect 9581 10570 9647 10573
rect 4846 10568 9647 10570
rect 4846 10512 9586 10568
rect 9642 10512 9647 10568
rect 4846 10510 9647 10512
rect 0 10434 480 10464
rect 4846 10434 4906 10510
rect 9581 10507 9647 10510
rect 0 10374 4906 10434
rect 0 10344 480 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 4061 10162 4127 10165
rect 5809 10162 5875 10165
rect 4061 10160 5875 10162
rect 4061 10104 4066 10160
rect 4122 10104 5814 10160
rect 5870 10104 5875 10160
rect 4061 10102 5875 10104
rect 4061 10099 4127 10102
rect 5809 10099 5875 10102
rect 0 10026 480 10056
rect 3601 10026 3667 10029
rect 0 10024 3667 10026
rect 0 9968 3606 10024
rect 3662 9968 3667 10024
rect 0 9966 3667 9968
rect 0 9936 480 9966
rect 3601 9963 3667 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 11053 9754 11119 9757
rect 11053 9752 11162 9754
rect 11053 9696 11058 9752
rect 11114 9696 11162 9752
rect 11053 9691 11162 9696
rect 0 9482 480 9512
rect 3141 9482 3207 9485
rect 0 9480 3207 9482
rect 0 9424 3146 9480
rect 3202 9424 3207 9480
rect 0 9422 3207 9424
rect 0 9392 480 9422
rect 3141 9419 3207 9422
rect 9949 9482 10015 9485
rect 11102 9482 11162 9691
rect 9949 9480 11162 9482
rect 9949 9424 9954 9480
rect 10010 9424 11162 9480
rect 9949 9422 11162 9424
rect 9949 9419 10015 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 0 9014 4906 9074
rect 0 8984 480 9014
rect 4846 8802 4906 9014
rect 9581 8802 9647 8805
rect 4846 8800 9647 8802
rect 4846 8744 9586 8800
rect 9642 8744 9647 8800
rect 4846 8742 9647 8744
rect 9581 8739 9647 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 3877 8530 3943 8533
rect 0 8528 3943 8530
rect 0 8472 3882 8528
rect 3938 8472 3943 8528
rect 0 8470 3943 8472
rect 0 8440 480 8470
rect 3877 8467 3943 8470
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 3325 8122 3391 8125
rect 0 8120 3391 8122
rect 0 8064 3330 8120
rect 3386 8064 3391 8120
rect 0 8062 3391 8064
rect 0 8032 480 8062
rect 3325 8059 3391 8062
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3969 7578 4035 7581
rect 0 7576 4035 7578
rect 0 7520 3974 7576
rect 4030 7520 4035 7576
rect 0 7518 4035 7520
rect 0 7488 480 7518
rect 3969 7515 4035 7518
rect 0 7170 480 7200
rect 3877 7170 3943 7173
rect 0 7168 3943 7170
rect 0 7112 3882 7168
rect 3938 7112 3943 7168
rect 0 7110 3943 7112
rect 0 7080 480 7110
rect 3877 7107 3943 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 8753 6762 8819 6765
rect 0 6760 8819 6762
rect 0 6704 8758 6760
rect 8814 6704 8819 6760
rect 0 6702 8819 6704
rect 0 6672 480 6702
rect 8753 6699 8819 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 480 6248
rect 7189 6218 7255 6221
rect 0 6216 7255 6218
rect 0 6160 7194 6216
rect 7250 6160 7255 6216
rect 0 6158 7255 6160
rect 0 6128 480 6158
rect 7189 6155 7255 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 3969 5266 4035 5269
rect 0 5264 4035 5266
rect 0 5208 3974 5264
rect 4030 5208 4035 5264
rect 0 5206 4035 5208
rect 0 5176 480 5206
rect 3969 5203 4035 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 480 4798
rect 4061 4795 4127 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 2865 4314 2931 4317
rect 0 4312 2931 4314
rect 0 4256 2870 4312
rect 2926 4256 2931 4312
rect 0 4254 2931 4256
rect 0 4224 480 4254
rect 2865 4251 2931 4254
rect 0 3906 480 3936
rect 3417 3906 3483 3909
rect 0 3904 3483 3906
rect 0 3848 3422 3904
rect 3478 3848 3483 3904
rect 0 3846 3483 3848
rect 0 3816 480 3846
rect 3417 3843 3483 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 0 3498 480 3528
rect 3877 3498 3943 3501
rect 0 3496 3943 3498
rect 0 3440 3882 3496
rect 3938 3440 3943 3496
rect 0 3438 3943 3440
rect 0 3408 480 3438
rect 3877 3435 3943 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 480 2984
rect 3969 2954 4035 2957
rect 0 2952 4035 2954
rect 0 2896 3974 2952
rect 4030 2896 4035 2952
rect 0 2894 4035 2896
rect 0 2864 480 2894
rect 3969 2891 4035 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 5257 2546 5323 2549
rect 0 2544 5323 2546
rect 0 2488 5262 2544
rect 5318 2488 5323 2544
rect 0 2486 5323 2488
rect 0 2456 480 2486
rect 5257 2483 5323 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 4061 2002 4127 2005
rect 0 2000 4127 2002
rect 0 1944 4066 2000
rect 4122 1944 4127 2000
rect 0 1942 4127 1944
rect 0 1912 480 1942
rect 4061 1939 4127 1942
rect 0 1594 480 1624
rect 3693 1594 3759 1597
rect 0 1592 3759 1594
rect 0 1536 3698 1592
rect 3754 1536 3759 1592
rect 0 1534 3759 1536
rect 0 1504 480 1534
rect 3693 1531 3759 1534
rect 0 1050 480 1080
rect 3233 1050 3299 1053
rect 0 1048 3299 1050
rect 0 992 3238 1048
rect 3294 992 3299 1048
rect 0 990 3299 992
rect 0 960 480 990
rect 3233 987 3299 990
rect 0 642 480 672
rect 3601 642 3667 645
rect 0 640 3667 642
rect 0 584 3606 640
rect 3662 584 3667 640
rect 0 582 3667 584
rect 0 552 480 582
rect 3601 579 3667 582
rect 0 234 480 264
rect 4705 234 4771 237
rect 0 232 4771 234
rect 0 176 4710 232
rect 4766 176 4771 232
rect 0 174 4771 176
rect 0 144 480 174
rect 4705 171 4771 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606821651
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606821651
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606821651
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606821651
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606821651
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606821651
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606821651
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606821651
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606821651
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606821651
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1606821651
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606821651
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1606821651
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1606821651
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606821651
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606821651
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1606821651
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606821651
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1606821651
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1606821651
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606821651
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606821651
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606821651
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606821651
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606821651
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1606821651
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1606821651
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1606821651
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1606821651
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606821651
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1606821651
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1606821651
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1606821651
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606821651
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606821651
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606821651
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606821651
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606821651
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606821651
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1606821651
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606821651
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1606821651
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1606821651
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1606821651
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606821651
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606821651
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606821651
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606821651
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606821651
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606821651
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606821651
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606821651
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1606821651
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1606821651
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1606821651
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1606821651
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1606821651
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1606821651
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606821651
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606821651
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606821651
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606821651
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1606821651
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1606821651
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1606821651
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1606821651
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1606821651
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1606821651
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp 1606821651
transform 1 0 20240 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1606821651
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606821651
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606821651
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606821651
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606821651
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606821651
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606821651
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606821651
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606821651
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606821651
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606821651
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1606821651
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1606821651
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1606821651
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1606821651
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1606821651
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1606821651
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1606821651
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1606821651
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1606821651
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1606821651
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1606821651
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1606821651
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1606821651
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1606821651
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606821651
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606821651
transform 1 0 19872 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1606821651
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_202
timestamp 1606821651
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1606821651
transform 1 0 19136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606821651
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606821651
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606821651
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1606821651
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _067_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_46
timestamp 1606821651
transform 1 0 5336 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_58
timestamp 1606821651
transform 1 0 6440 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8188 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7084 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1606821651
transform 1 0 6992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_74
timestamp 1606821651
transform 1 0 7912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_86
timestamp 1606821651
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1606821651
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1606821651
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1606821651
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1606821651
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1606821651
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1606821651
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606821651
transform 1 0 19412 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_190
timestamp 1606821651
transform 1 0 18584 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_198
timestamp 1606821651
transform 1 0 19320 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_203
timestamp 1606821651
transform 1 0 19780 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1606821651
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606821651
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2944 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1606821651
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1606821651
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4600 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1606821651
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_54
timestamp 1606821651
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606821651
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 8280 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7268 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1606821651
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1606821651
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_87
timestamp 1606821651
transform 1 0 9108 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1606821651
transform 1 0 10212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_111
timestamp 1606821651
transform 1 0 11316 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1606821651
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1606821651
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1606821651
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1606821651
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1606821651
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606821651
transform 1 0 18952 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_192
timestamp 1606821651
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_198
timestamp 1606821651
transform 1 0 19320 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_210
timestamp 1606821651
transform 1 0 20424 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_218
timestamp 1606821651
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2024 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1606821651
transform 1 0 1932 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_16
timestamp 1606821651
transform 1 0 2576 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1606821651
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1606821651
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5060 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6716 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1606821651
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8372 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 1606821651
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1606821651
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1606821651
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1606821651
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1606821651
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1606821651
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1606821651
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_178
timestamp 1606821651
transform 1 0 17480 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1606821651
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606821651
transform 1 0 18400 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_192
timestamp 1606821651
transform 1 0 18768 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1606821651
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1606821651
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606821651
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2116 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1606821651
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1606821651
transform 1 0 3588 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 1606821651
transform 1 0 3956 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1606821651
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1606821651
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1606821651
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7084 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8740 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1606821651
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_92
timestamp 1606821651
transform 1 0 9568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_104
timestamp 1606821651
transform 1 0 10672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_116
timestamp 1606821651
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1606821651
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1606821651
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1606821651
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1606821651
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606821651
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606821651
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606821651
transform 1 0 2300 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606821651
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1606821651
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_17
timestamp 1606821651
transform 1 0 2668 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4692 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606821651
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1606821651
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606821651
transform 1 0 6348 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_48
timestamp 1606821651
transform 1 0 5520 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1606821651
transform 1 0 6256 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_60
timestamp 1606821651
transform 1 0 6624 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7912 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1606821651
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_114
timestamp 1606821651
transform 1 0 11592 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_126
timestamp 1606821651
transform 1 0 12696 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_138
timestamp 1606821651
transform 1 0 13800 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1606821651
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1606821651
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1606821651
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1606821651
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1606821651
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606821651
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_15
timestamp 1606821651
transform 1 0 2484 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606821651
transform 1 0 3404 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1606821651
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_41
timestamp 1606821651
transform 1 0 4876 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1606821651
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1606821651
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5704 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_49
timestamp 1606821651
transform 1 0 5612 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1606821651
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_71
timestamp 1606821651
transform 1 0 7636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_66
timestamp 1606821651
transform 1 0 7176 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_74
timestamp 1606821651
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1606821651
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1606821651
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10948 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12604 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1606821651
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_105
timestamp 1606821651
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1606821651
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1606821651
transform 1 0 13524 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_139
timestamp 1606821651
transform 1 0 13892 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1606821651
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16376 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1606821651
transform 1 0 14812 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1606821651
transform 1 0 15916 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_164
timestamp 1606821651
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16560 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1606821651
transform 1 0 16468 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_177
timestamp 1606821651
transform 1 0 17388 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_182
timestamp 1606821651
transform 1 0 17848 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1606821651
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1606821651
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_194
timestamp 1606821651
transform 1 0 18952 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1606821651
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606821651
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1606821651
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1606821651
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1606821651
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_41
timestamp 1606821651
transform 1 0 4876 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5796 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1606821651
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_54
timestamp 1606821651
transform 1 0 6072 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1606821651
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1606821651
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10028 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 9476 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1606821651
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_94
timestamp 1606821651
transform 1 0 9752 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1606821651
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1606821651
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13156 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_126
timestamp 1606821651
transform 1 0 12696 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_130
timestamp 1606821651
transform 1 0 13064 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606821651
transform 1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15732 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_147
timestamp 1606821651
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_152
timestamp 1606821651
transform 1 0 15088 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_158
timestamp 1606821651
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606821651
transform 1 0 17388 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1606821651
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1606821651
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_200
timestamp 1606821651
transform 1 0 19504 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1606821651
transform 1 0 20608 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2852 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1932 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1606821651
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1606821651
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606821651
transform 1 0 4508 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1606821651
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1606821651
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_40
timestamp 1606821651
transform 1 0 4784 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_52
timestamp 1606821651
transform 1 0 5888 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7452 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1606821651
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606821651
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1606821651
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10764 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11868 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_114
timestamp 1606821651
transform 1 0 11592 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_126
timestamp 1606821651
transform 1 0 12696 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1606821651
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_163
timestamp 1606821651
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_175
timestamp 1606821651
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_187
timestamp 1606821651
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_199
timestamp 1606821651
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1606821651
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2760 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1748 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1606821651
transform 1 0 2300 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_17
timestamp 1606821651
transform 1 0 2668 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4416 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1606821651
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_45
timestamp 1606821651
transform 1 0 5244 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1606821651
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7912 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_71
timestamp 1606821651
transform 1 0 7636 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606821651
transform 1 0 9660 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10120 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_90
timestamp 1606821651
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1606821651
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_114
timestamp 1606821651
transform 1 0 11592 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_118
timestamp 1606821651
transform 1 0 11960 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14168 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13432 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1606821651
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1606821651
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15824 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1606821651
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606821651
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1606821651
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606821651
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19688 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_195
timestamp 1606821651
transform 1 0 19044 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_201
timestamp 1606821651
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1606821651
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2760 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1606821651
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1606821651
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_24
timestamp 1606821651
transform 1 0 3312 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1606821651
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5704 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1606821651
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7452 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_66
timestamp 1606821651
transform 1 0 7176 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_78
timestamp 1606821651
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10120 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606821651
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1606821651
transform 1 0 10028 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11408 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1606821651
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_111
timestamp 1606821651
transform 1 0 11316 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13708 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_128
timestamp 1606821651
transform 1 0 12880 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_136
timestamp 1606821651
transform 1 0 13616 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15456 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1606821651
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1606821651
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1606821651
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606821651
transform 1 0 16468 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17296 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 16928 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1606821651
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_175
timestamp 1606821651
transform 1 0 17204 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18952 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1606821651
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_203
timestamp 1606821651
transform 1 0 19780 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1606821651
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606821651
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1606821651
transform 1 0 1932 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1606821651
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1606821651
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606821651
transform 1 0 2300 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606821651
transform 1 0 2852 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_16
timestamp 1606821651
transform 1 0 2576 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4692 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_23
timestamp 1606821651
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_36
timestamp 1606821651
transform 1 0 4416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1606821651
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_40
timestamp 1606821651
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4968 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_55
timestamp 1606821651
transform 1 0 6164 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp 1606821651
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_62
timestamp 1606821651
transform 1 0 6808 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1606821651
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8096 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8188 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 7268 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1606821651
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_70
timestamp 1606821651
transform 1 0 7544 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1606821651
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1606821651
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606821651
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_86
timestamp 1606821651
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_92
timestamp 1606821651
transform 1 0 9568 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1606821651
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_100
timestamp 1606821651
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10580 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12604 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10764 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1606821651
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13156 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13800 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1606821651
transform 1 0 12696 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1606821651
transform 1 0 13064 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_134
timestamp 1606821651
transform 1 0 13432 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606821651
transform 1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15548 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_147
timestamp 1606821651
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1606821651
transform 1 0 15088 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_156
timestamp 1606821651
transform 1 0 15456 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_147
timestamp 1606821651
transform 1 0 14628 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1606821651
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16836 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_173
timestamp 1606821651
transform 1 0 17020 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606821651
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_187
timestamp 1606821651
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1606821651
transform 1 0 18860 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1606821651
transform 1 0 19964 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_199
timestamp 1606821651
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1606821651
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1606821651
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1932 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1606821651
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_15
timestamp 1606821651
transform 1 0 2484 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606821651
transform 1 0 3128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_21
timestamp 1606821651
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1606821651
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_36
timestamp 1606821651
transform 1 0 4416 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4968 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1606821651
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8372 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_71
timestamp 1606821651
transform 1 0 7636 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_95
timestamp 1606821651
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12512 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1606821651
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1606821651
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13892 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_133
timestamp 1606821651
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_138
timestamp 1606821651
transform 1 0 13800 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16008 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_148
timestamp 1606821651
transform 1 0 14720 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1606821651
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1606821651
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1606821651
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1606821651
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1606821651
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606821651
transform 1 0 1564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_9
timestamp 1606821651
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_17
timestamp 1606821651
transform 1 0 2668 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1606821651
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606821651
transform 1 0 6164 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6624 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_48
timestamp 1606821651
transform 1 0 5520 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_54
timestamp 1606821651
transform 1 0 6072 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1606821651
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8280 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1606821651
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10580 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1606821651
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1606821651
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_96
timestamp 1606821651
transform 1 0 9936 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_102
timestamp 1606821651
transform 1 0 10488 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12236 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_119
timestamp 1606821651
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 13432 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_130
timestamp 1606821651
transform 1 0 13064 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15824 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_150
timestamp 1606821651
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606821651
transform 1 0 17848 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_169
timestamp 1606821651
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_180
timestamp 1606821651
transform 1 0 17664 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_185
timestamp 1606821651
transform 1 0 18124 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18400 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_204
timestamp 1606821651
transform 1 0 19872 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1606821651
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606821651
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2760 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1932 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1606821651
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_15
timestamp 1606821651
transform 1 0 2484 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_34
timestamp 1606821651
transform 1 0 4232 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5612 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_46
timestamp 1606821651
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1606821651
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8740 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_78
timestamp 1606821651
transform 1 0 8280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_82
timestamp 1606821651
transform 1 0 8648 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_99
timestamp 1606821651
transform 1 0 10212 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606821651
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 14352 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13340 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1606821651
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_142
timestamp 1606821651
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15548 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1606821651
transform 1 0 15180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1606821651
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18308 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16560 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_177
timestamp 1606821651
transform 1 0 17388 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_203
timestamp 1606821651
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606821651
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606821651
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1932 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1606821651
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_15
timestamp 1606821651
transform 1 0 2484 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606821651
transform 1 0 3220 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4784 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_26
timestamp 1606821651
transform 1 0 3496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1606821651
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 6440 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1606821651
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_61
timestamp 1606821651
transform 1 0 6716 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 7820 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1606821651
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_76
timestamp 1606821651
transform 1 0 8096 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_80
timestamp 1606821651
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606821651
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1606821651
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10948 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_106
timestamp 1606821651
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_123
timestamp 1606821651
transform 1 0 12420 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13984 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1606821651
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15732 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 15456 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1606821651
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606821651
transform 1 0 17388 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1606821651
transform 1 0 17940 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_175
timestamp 1606821651
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_180
timestamp 1606821651
transform 1 0 17664 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606821651
transform 1 0 18952 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1606821651
transform 1 0 18768 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1606821651
transform 1 0 19228 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1606821651
transform 1 0 20332 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1606821651
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606821651
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2576 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1606821651
transform 1 0 2116 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1606821651
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4232 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_32
timestamp 1606821651
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1606821651
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5244 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1606821651
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1606821651
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_62
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7452 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_68
timestamp 1606821651
transform 1 0 7360 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_78
timestamp 1606821651
transform 1 0 8280 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9016 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_102
timestamp 1606821651
transform 1 0 10488 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 12604 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_114
timestamp 1606821651
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606821651
transform 1 0 12880 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13340 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1606821651
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16284 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14996 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1606821651
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_160
timestamp 1606821651
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1606821651
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1606821651
transform 1 0 18860 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1606821651
transform 1 0 19964 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_217
timestamp 1606821651
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1606821651
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_8
timestamp 1606821651
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1932 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606821651
transform 1 0 1472 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 1606821651
transform 1 0 2852 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1606821651
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_16
timestamp 1606821651
transform 1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2852 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2944 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_28
timestamp 1606821651
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1606821651
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_36
timestamp 1606821651
transform 1 0 4416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606821651
transform 1 0 6624 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4968 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5612 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_58
timestamp 1606821651
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_48
timestamp 1606821651
transform 1 0 5520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1606821651
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_62
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7452 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7084 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_63
timestamp 1606821651
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1606821651
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_68
timestamp 1606821651
transform 1 0 7360 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606821651
transform 1 0 9200 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1606821651
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1606821651
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_85
timestamp 1606821651
transform 1 0 8924 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1606821651
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10856 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12512 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_122
timestamp 1606821651
transform 1 0 12328 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_109
timestamp 1606821651
transform 1 0 11132 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1606821651
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606821651
transform 1 0 13432 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13524 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1606821651
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_144
timestamp 1606821651
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1606821651
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1606821651
transform 1 0 13708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1606821651
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1606821651
transform 1 0 14812 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_161
timestamp 1606821651
transform 1 0 15916 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17848 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_170
timestamp 1606821651
transform 1 0 16744 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1606821651
transform 1 0 16652 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1606821651
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_198
timestamp 1606821651
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_200
timestamp 1606821651
transform 1 0 19504 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1606821651
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_212
timestamp 1606821651
transform 1 0 20608 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606821651
transform 1 0 2668 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1932 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1606821651
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1606821651
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606821651
transform 1 0 3312 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1606821651
transform 1 0 3036 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1606821651
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5336 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_44
timestamp 1606821651
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_62
timestamp 1606821651
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6992 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_70
timestamp 1606821651
transform 1 0 7544 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_82
timestamp 1606821651
transform 1 0 8648 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606821651
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1606821651
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1606821651
transform 1 0 11592 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1606821651
transform 1 0 11960 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1606821651
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_146
timestamp 1606821651
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1606821651
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_163
timestamp 1606821651
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1606821651
transform 1 0 17388 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1606821651
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1606821651
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606821651
transform 1 0 18400 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_191
timestamp 1606821651
transform 1 0 18676 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_203
timestamp 1606821651
transform 1 0 19780 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1606821651
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606821651
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606821651
transform 1 0 1564 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2944 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1606821651
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_17
timestamp 1606821651
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_36
timestamp 1606821651
transform 1 0 4416 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606821651
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5244 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_44
timestamp 1606821651
transform 1 0 5152 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1606821651
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606821651
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 7084 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_71
timestamp 1606821651
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9844 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_86
timestamp 1606821651
transform 1 0 9016 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_94
timestamp 1606821651
transform 1 0 9752 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_111
timestamp 1606821651
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1606821651
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14260 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1606821651
transform 1 0 13892 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_152
timestamp 1606821651
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606821651
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_170
timestamp 1606821651
transform 1 0 16744 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_176
timestamp 1606821651
transform 1 0 17296 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606821651
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_190
timestamp 1606821651
transform 1 0 18584 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_202
timestamp 1606821651
transform 1 0 19688 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_214
timestamp 1606821651
transform 1 0 20792 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1932 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1606821651
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1606821651
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_19
timestamp 1606821651
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606821651
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_41
timestamp 1606821651
transform 1 0 4876 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5428 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606821651
transform 1 0 7176 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8648 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7636 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_63
timestamp 1606821651
transform 1 0 6900 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_69
timestamp 1606821651
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1606821651
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10028 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1606821651
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11868 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_113
timestamp 1606821651
transform 1 0 11500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_123
timestamp 1606821651
transform 1 0 12420 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13984 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1606821651
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16376 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15364 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_146
timestamp 1606821651
transform 1 0 14536 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1606821651
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_154
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_164
timestamp 1606821651
transform 1 0 16192 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18216 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17480 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_172
timestamp 1606821651
transform 1 0 16928 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1606821651
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_192
timestamp 1606821651
transform 1 0 18768 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1606821651
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1606821651
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606821651
transform 1 0 1656 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_10
timestamp 1606821651
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1606821651
transform 1 0 2760 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3220 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_22
timestamp 1606821651
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_39
timestamp 1606821651
transform 1 0 4692 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5060 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606821651
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_62
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7636 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_70
timestamp 1606821651
transform 1 0 7544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606821651
transform 1 0 9384 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9844 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_87
timestamp 1606821651
transform 1 0 9108 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1606821651
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606821651
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12604 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_111
timestamp 1606821651
transform 1 0 11316 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_115
timestamp 1606821651
transform 1 0 11684 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606821651
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606821651
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13340 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_131
timestamp 1606821651
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606821651
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1606821651
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606821651
transform 1 0 16284 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14628 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15548 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1606821651
transform 1 0 15180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1606821651
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17204 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1606821651
transform 1 0 16652 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1606821651
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606821651
transform 1 0 19320 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606821651
transform 1 0 18768 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 19964 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_190
timestamp 1606821651
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1606821651
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_202
timestamp 1606821651
transform 1 0 19688 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_217
timestamp 1606821651
transform 1 0 21068 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606821651
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606821651
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1606821651
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1606821651
transform 1 0 2668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606821651
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_25
timestamp 1606821651
transform 1 0 3404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1606821651
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_41
timestamp 1606821651
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5152 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1606821651
transform 1 0 5980 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1606821651
transform 1 0 6716 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8648 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_75
timestamp 1606821651
transform 1 0 8004 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_81
timestamp 1606821651
transform 1 0 8556 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1606821651
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_103
timestamp 1606821651
transform 1 0 10580 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_115
timestamp 1606821651
transform 1 0 11684 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_123
timestamp 1606821651
transform 1 0 12420 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606821651
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606821651
transform 1 0 13800 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13064 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1606821651
transform 1 0 12972 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1606821651
transform 1 0 13616 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_142
timestamp 1606821651
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606821651
transform 1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_148
timestamp 1606821651
transform 1 0 14720 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1606821651
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1606821651
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_166
timestamp 1606821651
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606821651
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606821651
transform 1 0 17112 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606821651
transform 1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_172
timestamp 1606821651
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1606821651
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1606821651
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_191
timestamp 1606821651
transform 1 0 18676 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_203
timestamp 1606821651
transform 1 0 19780 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606821651
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal3 s 22320 11432 22800 11552 6 ccff_head
port 0 nsew default input
rlabel metal2 s 11426 0 11482 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 3790 22320 3846 22800 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 8390 22320 8446 22800 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 8850 22320 8906 22800 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 9310 22320 9366 22800 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 9770 22320 9826 22800 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10230 22320 10286 22800 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 10690 22320 10746 22800 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 12438 22320 12494 22800 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 4250 22320 4306 22800 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 5170 22320 5226 22800 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 5630 22320 5686 22800 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 6090 22320 6146 22800 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 6550 22320 6606 22800 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 7010 22320 7066 22800 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 7470 22320 7526 22800 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 7930 22320 7986 22800 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 12898 22320 12954 22800 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 17958 22320 18014 22800 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18418 22320 18474 22800 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 18878 22320 18934 22800 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19338 22320 19394 22800 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 19798 22320 19854 22800 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20258 22320 20314 22800 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 20718 22320 20774 22800 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 21178 22320 21234 22800 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 21638 22320 21694 22800 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 13358 22320 13414 22800 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 13818 22320 13874 22800 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 14278 22320 14334 22800 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 14738 22320 14794 22800 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 15198 22320 15254 22800 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 15658 22320 15714 22800 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 16118 22320 16174 22800 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 16578 22320 16634 22800 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 17038 22320 17094 22800 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_11_
port 82 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_13_
port 83 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_15_
port 84 nsew default input
rlabel metal3 s 0 3816 480 3936 6 left_bottom_grid_pin_17_
port 85 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 86 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 87 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_5_
port 88 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_7_
port 89 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_9_
port 90 nsew default input
rlabel metal2 s 22098 22320 22154 22800 6 prog_clk_0_N_in
port 91 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 92 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_43_
port 93 nsew default input
rlabel metal2 s 1030 22320 1086 22800 6 top_left_grid_pin_44_
port 94 nsew default input
rlabel metal2 s 1490 22320 1546 22800 6 top_left_grid_pin_45_
port 95 nsew default input
rlabel metal2 s 1950 22320 2006 22800 6 top_left_grid_pin_46_
port 96 nsew default input
rlabel metal2 s 2410 22320 2466 22800 6 top_left_grid_pin_47_
port 97 nsew default input
rlabel metal2 s 2870 22320 2926 22800 6 top_left_grid_pin_48_
port 98 nsew default input
rlabel metal2 s 3330 22320 3386 22800 6 top_left_grid_pin_49_
port 99 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 top_right_grid_pin_1_
port 100 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 101 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 102 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
