magic
tech EFS8A
magscale 1 2
timestamp 1602252528
<< locali >>
rect 4439 6953 4445 6987
rect 4439 6885 4473 6953
rect 3335 3927 3369 3995
rect 3335 3893 3341 3927
rect 4439 3689 4445 3723
rect 4439 3621 4473 3689
rect 4531 2839 4565 2907
rect 4531 2805 4537 2839
rect 4439 2601 4445 2635
rect 4439 2533 4473 2601
rect 3249 2363 3283 2533
<< viali >>
rect 2605 8313 2639 8347
rect 1777 8245 1811 8279
rect 2329 8245 2363 8279
rect 2145 8041 2179 8075
rect 2558 7973 2592 8007
rect 2237 7837 2271 7871
rect 1685 7701 1719 7735
rect 4261 7701 4295 7735
rect 3801 7497 3835 7531
rect 1685 7293 1719 7327
rect 2145 7293 2179 7327
rect 2513 7293 2547 7327
rect 2881 7293 2915 7327
rect 3985 7293 4019 7327
rect 3433 7225 3467 7259
rect 4306 7225 4340 7259
rect 1961 7157 1995 7191
rect 4445 6953 4479 6987
rect 3157 6885 3191 6919
rect 1961 6817 1995 6851
rect 2145 6817 2179 6851
rect 2513 6817 2547 6851
rect 2881 6817 2915 6851
rect 3433 6749 3467 6783
rect 4077 6749 4111 6783
rect 3801 6613 3835 6647
rect 1777 6409 1811 6443
rect 4169 6409 4203 6443
rect 2145 6341 2179 6375
rect 3709 6273 3743 6307
rect 2237 6205 2271 6239
rect 2697 6205 2731 6239
rect 3065 6205 3099 6239
rect 3617 6205 3651 6239
rect 4445 6069 4479 6103
rect 4813 6069 4847 6103
rect 2513 5865 2547 5899
rect 2789 5865 2823 5899
rect 3525 5865 3559 5899
rect 4261 5865 4295 5899
rect 2145 5797 2179 5831
rect 2053 5729 2087 5763
rect 3157 5729 3191 5763
rect 2605 5321 2639 5355
rect 2881 5321 2915 5355
rect 1501 5185 1535 5219
rect 3801 5185 3835 5219
rect 4629 5185 4663 5219
rect 1685 5117 1719 5151
rect 3157 5117 3191 5151
rect 4537 5117 4571 5151
rect 4721 5117 4755 5151
rect 1869 5049 1903 5083
rect 2237 5049 2271 5083
rect 1777 4981 1811 5015
rect 4077 4981 4111 5015
rect 1685 4777 1719 4811
rect 2145 4777 2179 4811
rect 3433 4777 3467 4811
rect 3709 4777 3743 4811
rect 2237 4709 2271 4743
rect 2329 4709 2363 4743
rect 3065 4709 3099 4743
rect 1961 4641 1995 4675
rect 2697 4573 2731 4607
rect 4353 4437 4387 4471
rect 2421 4233 2455 4267
rect 2789 4233 2823 4267
rect 1409 4097 1443 4131
rect 4169 4097 4203 4131
rect 1593 4029 1627 4063
rect 2973 4029 3007 4063
rect 4905 4029 4939 4063
rect 1777 3961 1811 3995
rect 2145 3961 2179 3995
rect 1685 3893 1719 3927
rect 3341 3893 3375 3927
rect 4629 3893 4663 3927
rect 1593 3689 1627 3723
rect 2605 3689 2639 3723
rect 3709 3689 3743 3723
rect 4445 3689 4479 3723
rect 1961 3621 1995 3655
rect 2329 3621 2363 3655
rect 2697 3621 2731 3655
rect 2513 3553 2547 3587
rect 3341 3553 3375 3587
rect 3065 3485 3099 3519
rect 4077 3485 4111 3519
rect 5273 3485 5307 3519
rect 1685 3145 1719 3179
rect 4077 3145 4111 3179
rect 5733 3145 5767 3179
rect 3249 3077 3283 3111
rect 3617 3009 3651 3043
rect 4169 3009 4203 3043
rect 6101 3009 6135 3043
rect 1869 2941 1903 2975
rect 2605 2941 2639 2975
rect 2789 2941 2823 2975
rect 3065 2941 3099 2975
rect 4537 2805 4571 2839
rect 5365 2805 5399 2839
rect 1961 2601 1995 2635
rect 4445 2601 4479 2635
rect 5273 2601 5307 2635
rect 2599 2533 2633 2567
rect 3249 2533 3283 2567
rect 2237 2397 2271 2431
rect 4077 2465 4111 2499
rect 5641 2465 5675 2499
rect 6009 2397 6043 2431
rect 3249 2329 3283 2363
rect 3525 2329 3559 2363
rect 3801 2329 3835 2363
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1946 8304 1952 8356
rect 2004 8344 2010 8356
rect 2593 8347 2651 8353
rect 2593 8344 2605 8347
rect 2004 8316 2605 8344
rect 2004 8304 2010 8316
rect 2593 8313 2605 8316
rect 2639 8313 2651 8347
rect 2593 8307 2651 8313
rect 1762 8276 1768 8288
rect 1723 8248 1768 8276
rect 1762 8236 1768 8248
rect 1820 8236 1826 8288
rect 2314 8276 2320 8288
rect 2275 8248 2320 8276
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2866 8072 2872 8084
rect 2179 8044 2872 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 2314 7964 2320 8016
rect 2372 8004 2378 8016
rect 2546 8007 2604 8013
rect 2546 8004 2558 8007
rect 2372 7976 2558 8004
rect 2372 7964 2378 7976
rect 2546 7973 2558 7976
rect 2592 7973 2604 8007
rect 2546 7967 2604 7973
rect 1946 7828 1952 7880
rect 2004 7868 2010 7880
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 2004 7840 2237 7868
rect 2004 7828 2010 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 4212 7704 4261 7732
rect 4212 7692 4218 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 3789 7531 3847 7537
rect 3789 7528 3801 7531
rect 2372 7500 3801 7528
rect 2372 7488 2378 7500
rect 3789 7497 3801 7500
rect 3835 7497 3847 7531
rect 3789 7491 3847 7497
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 1762 7284 1768 7336
rect 1820 7324 1826 7336
rect 2130 7324 2136 7336
rect 1820 7296 2136 7324
rect 1820 7284 1826 7296
rect 2130 7284 2136 7296
rect 2188 7284 2194 7336
rect 2498 7324 2504 7336
rect 2459 7296 2504 7324
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 2866 7324 2872 7336
rect 2827 7296 2872 7324
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 2516 7256 2544 7284
rect 3421 7259 3479 7265
rect 3421 7256 3433 7259
rect 2516 7228 3433 7256
rect 3421 7225 3433 7228
rect 3467 7225 3479 7259
rect 3804 7256 3832 7491
rect 3970 7324 3976 7336
rect 3931 7296 3976 7324
rect 3970 7284 3976 7296
rect 4028 7324 4034 7336
rect 4154 7324 4160 7336
rect 4028 7296 4160 7324
rect 4028 7284 4034 7296
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4294 7259 4352 7265
rect 4294 7256 4306 7259
rect 3804 7228 4306 7256
rect 3421 7219 3479 7225
rect 4294 7225 4306 7228
rect 4340 7256 4352 7259
rect 4430 7256 4436 7268
rect 4340 7228 4436 7256
rect 4340 7225 4352 7228
rect 4294 7219 4352 7225
rect 4430 7216 4436 7228
rect 4488 7216 4494 7268
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 4430 6984 4436 6996
rect 4391 6956 4436 6984
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 3145 6919 3203 6925
rect 3145 6885 3157 6919
rect 3191 6916 3203 6919
rect 3970 6916 3976 6928
rect 3191 6888 3976 6916
rect 3191 6885 3203 6888
rect 3145 6879 3203 6885
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 1946 6848 1952 6860
rect 1907 6820 1952 6848
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2130 6848 2136 6860
rect 2091 6820 2136 6848
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 2498 6848 2504 6860
rect 2459 6820 2504 6848
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2866 6848 2872 6860
rect 2827 6820 2872 6848
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 1964 6780 1992 6808
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 1964 6752 3433 6780
rect 3421 6749 3433 6752
rect 3467 6780 3479 6783
rect 3510 6780 3516 6792
rect 3467 6752 3516 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 4062 6780 4068 6792
rect 4023 6752 4068 6780
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 2866 6440 2872 6452
rect 1811 6412 2872 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4430 6440 4436 6452
rect 4203 6412 4436 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 2133 6375 2191 6381
rect 2133 6341 2145 6375
rect 2179 6372 2191 6375
rect 2498 6372 2504 6384
rect 2179 6344 2504 6372
rect 2179 6341 2191 6344
rect 2133 6335 2191 6341
rect 2498 6332 2504 6344
rect 2556 6332 2562 6384
rect 2516 6304 2544 6332
rect 3697 6307 3755 6313
rect 2516 6276 3096 6304
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 3068 6245 3096 6276
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 4062 6304 4068 6316
rect 3743 6276 4068 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 2225 6239 2283 6245
rect 2225 6236 2237 6239
rect 2004 6208 2237 6236
rect 2004 6196 2010 6208
rect 2225 6205 2237 6208
rect 2271 6205 2283 6239
rect 2225 6199 2283 6205
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6236 3663 6239
rect 3786 6236 3792 6248
rect 3651 6208 3792 6236
rect 3651 6205 3663 6208
rect 3605 6199 3663 6205
rect 2130 6128 2136 6180
rect 2188 6168 2194 6180
rect 2700 6168 2728 6199
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 2188 6140 2728 6168
rect 2188 6128 2194 6140
rect 2700 6100 2728 6140
rect 4126 6140 4384 6168
rect 4126 6100 4154 6140
rect 4356 6112 4384 6140
rect 2700 6072 4154 6100
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 4396 6072 4445 6100
rect 4396 6060 4402 6072
rect 4433 6069 4445 6072
rect 4479 6100 4491 6103
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4479 6072 4813 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 2498 5896 2504 5908
rect 1544 5868 2504 5896
rect 1544 5856 1550 5868
rect 2498 5856 2504 5868
rect 2556 5896 2562 5908
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 2556 5868 2789 5896
rect 2556 5856 2562 5868
rect 2777 5865 2789 5868
rect 2823 5865 2835 5899
rect 3510 5896 3516 5908
rect 3471 5868 3516 5896
rect 2777 5859 2835 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4120 5868 4261 5896
rect 4120 5856 4126 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4249 5859 4307 5865
rect 2130 5828 2136 5840
rect 2091 5800 2136 5828
rect 2130 5788 2136 5800
rect 2188 5788 2194 5840
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 1912 5732 2053 5760
rect 1912 5720 1918 5732
rect 2041 5729 2053 5732
rect 2087 5760 2099 5763
rect 3145 5763 3203 5769
rect 3145 5760 3157 5763
rect 2087 5732 3157 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 3145 5729 3157 5732
rect 3191 5729 3203 5763
rect 3145 5723 3203 5729
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 1688 5324 2605 5352
rect 1486 5216 1492 5228
rect 1447 5188 1492 5216
rect 1486 5176 1492 5188
rect 1544 5176 1550 5228
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 1688 5157 1716 5324
rect 2593 5321 2605 5324
rect 2639 5352 2651 5355
rect 2866 5352 2872 5364
rect 2639 5324 2872 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 1762 5244 1768 5296
rect 1820 5284 1826 5296
rect 1820 5256 4752 5284
rect 1820 5244 1826 5256
rect 3786 5216 3792 5228
rect 3747 5188 3792 5216
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4120 5188 4629 5216
rect 4120 5176 4126 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 1673 5151 1731 5157
rect 1673 5148 1685 5151
rect 1636 5120 1685 5148
rect 1636 5108 1642 5120
rect 1673 5117 1685 5120
rect 1719 5117 1731 5151
rect 1673 5111 1731 5117
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 2924 5120 3157 5148
rect 2924 5108 2930 5120
rect 3145 5117 3157 5120
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 1854 5080 1860 5092
rect 1815 5052 1860 5080
rect 1854 5040 1860 5052
rect 1912 5040 1918 5092
rect 2222 5080 2228 5092
rect 2183 5052 2228 5080
rect 2222 5040 2228 5052
rect 2280 5040 2286 5092
rect 3804 5080 3832 5176
rect 4724 5157 4752 5256
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4709 5151 4767 5157
rect 4709 5148 4721 5151
rect 4571 5120 4721 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 4709 5117 4721 5120
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 4614 5080 4620 5092
rect 3804 5052 4620 5080
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 106 4972 112 5024
rect 164 5012 170 5024
rect 1670 5012 1676 5024
rect 164 4984 1676 5012
rect 164 4972 170 4984
rect 1670 4972 1676 4984
rect 1728 5012 1734 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 1728 4984 1777 5012
rect 1728 4972 1734 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 1765 4975 1823 4981
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 3476 4984 4077 5012
rect 3476 4972 3482 4984
rect 4065 4981 4077 4984
rect 4111 4981 4123 5015
rect 4065 4975 4123 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 1854 4768 1860 4820
rect 1912 4808 1918 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1912 4780 2145 4808
rect 1912 4768 1918 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 3418 4808 3424 4820
rect 3379 4780 3424 4808
rect 2133 4771 2191 4777
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3697 4811 3755 4817
rect 3697 4808 3709 4811
rect 3568 4780 3709 4808
rect 3568 4768 3574 4780
rect 3697 4777 3709 4780
rect 3743 4808 3755 4811
rect 4062 4808 4068 4820
rect 3743 4780 4068 4808
rect 3743 4777 3755 4780
rect 3697 4771 3755 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 1486 4700 1492 4752
rect 1544 4740 1550 4752
rect 2225 4743 2283 4749
rect 2225 4740 2237 4743
rect 1544 4712 2237 4740
rect 1544 4700 1550 4712
rect 2225 4709 2237 4712
rect 2271 4709 2283 4743
rect 2225 4703 2283 4709
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 2406 4740 2412 4752
rect 2363 4712 2412 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 1949 4675 2007 4681
rect 1949 4672 1961 4675
rect 1728 4644 1961 4672
rect 1728 4632 1734 4644
rect 1949 4641 1961 4644
rect 1995 4641 2007 4675
rect 2240 4672 2268 4703
rect 2406 4700 2412 4712
rect 2464 4700 2470 4752
rect 3053 4743 3111 4749
rect 3053 4709 3065 4743
rect 3099 4740 3111 4743
rect 3234 4740 3240 4752
rect 3099 4712 3240 4740
rect 3099 4709 3111 4712
rect 3053 4703 3111 4709
rect 3234 4700 3240 4712
rect 3292 4740 3298 4752
rect 4430 4740 4436 4752
rect 3292 4712 4436 4740
rect 3292 4700 3298 4712
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 2774 4672 2780 4684
rect 2240 4644 2780 4672
rect 1949 4635 2007 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 4154 4604 4160 4616
rect 2731 4576 4160 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 4341 4471 4399 4477
rect 4341 4437 4353 4471
rect 4387 4468 4399 4471
rect 4614 4468 4620 4480
rect 4387 4440 4620 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 2409 4267 2467 4273
rect 2409 4264 2421 4267
rect 1728 4236 2421 4264
rect 1728 4224 1734 4236
rect 2409 4233 2421 4236
rect 2455 4233 2467 4267
rect 2774 4264 2780 4276
rect 2735 4236 2780 4264
rect 2409 4227 2467 4233
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 1486 4128 1492 4140
rect 1443 4100 1492 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 3326 4088 3332 4140
rect 3384 4128 3390 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 3384 4100 4169 4128
rect 3384 4088 3390 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 1578 4060 1584 4072
rect 1539 4032 1584 4060
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 2958 4060 2964 4072
rect 2919 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4060 3022 4072
rect 4893 4063 4951 4069
rect 4893 4060 4905 4063
rect 3016 4032 4905 4060
rect 3016 4020 3022 4032
rect 4893 4029 4905 4032
rect 4939 4029 4951 4063
rect 4893 4023 4951 4029
rect 1762 3992 1768 4004
rect 1723 3964 1768 3992
rect 1762 3952 1768 3964
rect 1820 3952 1826 4004
rect 2130 3992 2136 4004
rect 2091 3964 2136 3992
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 1673 3927 1731 3933
rect 1673 3893 1685 3927
rect 1719 3924 1731 3927
rect 1946 3924 1952 3936
rect 1719 3896 1952 3924
rect 1719 3893 1731 3896
rect 1673 3887 1731 3893
rect 1946 3884 1952 3896
rect 2004 3924 2010 3936
rect 2314 3924 2320 3936
rect 2004 3896 2320 3924
rect 2004 3884 2010 3896
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 3329 3927 3387 3933
rect 3329 3924 3341 3927
rect 3292 3896 3341 3924
rect 3292 3884 3298 3896
rect 3329 3893 3341 3896
rect 3375 3893 3387 3927
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 3329 3887 3387 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 2593 3723 2651 3729
rect 2593 3720 2605 3723
rect 1964 3692 2605 3720
rect 1486 3612 1492 3664
rect 1544 3652 1550 3664
rect 1964 3661 1992 3692
rect 2593 3689 2605 3692
rect 2639 3720 2651 3723
rect 2774 3720 2780 3732
rect 2639 3692 2780 3720
rect 2639 3689 2651 3692
rect 2593 3683 2651 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 3697 3723 3755 3729
rect 3697 3720 3709 3723
rect 3568 3692 3709 3720
rect 3568 3680 3574 3692
rect 3697 3689 3709 3692
rect 3743 3689 3755 3723
rect 4430 3720 4436 3732
rect 4391 3692 4436 3720
rect 3697 3683 3755 3689
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 1949 3655 2007 3661
rect 1949 3652 1961 3655
rect 1544 3624 1961 3652
rect 1544 3612 1550 3624
rect 1949 3621 1961 3624
rect 1995 3621 2007 3655
rect 2314 3652 2320 3664
rect 2275 3624 2320 3652
rect 1949 3615 2007 3621
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 2406 3612 2412 3664
rect 2464 3652 2470 3664
rect 2685 3655 2743 3661
rect 2685 3652 2697 3655
rect 2464 3624 2697 3652
rect 2464 3612 2470 3624
rect 2685 3621 2697 3624
rect 2731 3652 2743 3655
rect 3050 3652 3056 3664
rect 2731 3624 3056 3652
rect 2731 3621 2743 3624
rect 2685 3615 2743 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 2501 3587 2559 3593
rect 2501 3584 2513 3587
rect 1820 3556 2513 3584
rect 1820 3544 1826 3556
rect 2501 3553 2513 3556
rect 2547 3584 2559 3587
rect 3326 3584 3332 3596
rect 2547 3556 3332 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3099 3488 4077 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 4065 3485 4077 3488
rect 4111 3516 4123 3519
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 4111 3488 5273 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 4430 3176 4436 3188
rect 4111 3148 4436 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 4672 3148 5733 3176
rect 4672 3136 4678 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 2958 3068 2964 3120
rect 3016 3108 3022 3120
rect 3237 3111 3295 3117
rect 3237 3108 3249 3111
rect 3016 3080 3249 3108
rect 3016 3068 3022 3080
rect 3237 3077 3249 3080
rect 3283 3077 3295 3111
rect 3237 3071 3295 3077
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 2792 3012 3617 3040
rect 2792 2984 2820 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 6089 3043 6147 3049
rect 6089 3040 6101 3043
rect 4212 3012 6101 3040
rect 4212 3000 4218 3012
rect 6089 3009 6101 3012
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1728 2944 1869 2972
rect 1728 2932 1734 2944
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2941 2651 2975
rect 2774 2972 2780 2984
rect 2735 2944 2780 2972
rect 2593 2935 2651 2941
rect 2608 2904 2636 2935
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 3050 2972 3056 2984
rect 3011 2944 3056 2972
rect 3050 2932 3056 2944
rect 3108 2972 3114 2984
rect 4614 2972 4620 2984
rect 3108 2944 4620 2972
rect 3108 2932 3114 2944
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 4338 2904 4344 2916
rect 2608 2876 4344 2904
rect 4338 2864 4344 2876
rect 4396 2904 4402 2916
rect 5258 2904 5264 2916
rect 4396 2876 5264 2904
rect 4396 2864 4402 2876
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 4430 2796 4436 2848
rect 4488 2836 4494 2848
rect 4525 2839 4583 2845
rect 4525 2836 4537 2839
rect 4488 2808 4537 2836
rect 4488 2796 4494 2808
rect 4525 2805 4537 2808
rect 4571 2836 4583 2839
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 4571 2808 5365 2836
rect 4571 2805 4583 2808
rect 4525 2799 4583 2805
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 5353 2799 5411 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2774 2632 2780 2644
rect 1995 2604 2780 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4522 2632 4528 2644
rect 4479 2604 4528 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 5258 2632 5264 2644
rect 5219 2604 5264 2632
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 2587 2567 2645 2573
rect 2587 2533 2599 2567
rect 2633 2564 2645 2567
rect 3237 2567 3295 2573
rect 3237 2564 3249 2567
rect 2633 2536 3249 2564
rect 2633 2533 2645 2536
rect 2587 2527 2645 2533
rect 3237 2533 3249 2536
rect 3283 2533 3295 2567
rect 3237 2527 3295 2533
rect 2130 2456 2136 2508
rect 2188 2496 2194 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 2188 2468 4077 2496
rect 2188 2456 2194 2468
rect 4065 2465 4077 2468
rect 4111 2496 4123 2499
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 4111 2468 5641 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5629 2465 5641 2468
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 2222 2388 2228 2400
rect 2280 2428 2286 2440
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 2280 2400 6009 2428
rect 2280 2388 2286 2400
rect 5997 2397 6009 2400
rect 6043 2397 6055 2431
rect 5997 2391 6055 2397
rect 3237 2363 3295 2369
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 3513 2363 3571 2369
rect 3513 2360 3525 2363
rect 3283 2332 3525 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 3513 2329 3525 2332
rect 3559 2360 3571 2363
rect 3789 2363 3847 2369
rect 3789 2360 3801 2363
rect 3559 2332 3801 2360
rect 3559 2329 3571 2332
rect 3513 2323 3571 2329
rect 3789 2329 3801 2332
rect 3835 2360 3847 2363
rect 4062 2360 4068 2372
rect 3835 2332 4068 2360
rect 3835 2329 3847 2332
rect 3789 2323 3847 2329
rect 4062 2320 4068 2332
rect 4120 2360 4126 2372
rect 4430 2360 4436 2372
rect 4120 2332 4436 2360
rect 4120 2320 4126 2332
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1952 8304 2004 8356
rect 1768 8279 1820 8288
rect 1768 8245 1777 8279
rect 1777 8245 1811 8279
rect 1811 8245 1820 8279
rect 1768 8236 1820 8245
rect 2320 8279 2372 8288
rect 2320 8245 2329 8279
rect 2329 8245 2363 8279
rect 2363 8245 2372 8279
rect 2320 8236 2372 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2872 8032 2924 8084
rect 2320 7964 2372 8016
rect 1952 7828 2004 7880
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 4160 7692 4212 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2320 7488 2372 7540
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 1768 7284 1820 7336
rect 2136 7327 2188 7336
rect 2136 7293 2145 7327
rect 2145 7293 2179 7327
rect 2179 7293 2188 7327
rect 2136 7284 2188 7293
rect 2504 7327 2556 7336
rect 2504 7293 2513 7327
rect 2513 7293 2547 7327
rect 2547 7293 2556 7327
rect 2504 7284 2556 7293
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 4160 7284 4212 7336
rect 4436 7216 4488 7268
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 4436 6987 4488 6996
rect 4436 6953 4445 6987
rect 4445 6953 4479 6987
rect 4479 6953 4488 6987
rect 4436 6944 4488 6953
rect 3976 6876 4028 6928
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 2136 6851 2188 6860
rect 2136 6817 2145 6851
rect 2145 6817 2179 6851
rect 2179 6817 2188 6851
rect 2136 6808 2188 6817
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 3516 6740 3568 6792
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2872 6400 2924 6452
rect 4436 6400 4488 6452
rect 2504 6332 2556 6384
rect 1952 6196 2004 6248
rect 4068 6264 4120 6316
rect 2136 6128 2188 6180
rect 3792 6196 3844 6248
rect 4344 6060 4396 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1492 5856 1544 5908
rect 2504 5899 2556 5908
rect 2504 5865 2513 5899
rect 2513 5865 2547 5899
rect 2547 5865 2556 5899
rect 2504 5856 2556 5865
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 4068 5856 4120 5908
rect 2136 5831 2188 5840
rect 2136 5797 2145 5831
rect 2145 5797 2179 5831
rect 2179 5797 2188 5831
rect 2136 5788 2188 5797
rect 1860 5720 1912 5772
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1492 5219 1544 5228
rect 1492 5185 1501 5219
rect 1501 5185 1535 5219
rect 1535 5185 1544 5219
rect 1492 5176 1544 5185
rect 1584 5108 1636 5160
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 1768 5244 1820 5296
rect 3792 5219 3844 5228
rect 3792 5185 3801 5219
rect 3801 5185 3835 5219
rect 3835 5185 3844 5219
rect 3792 5176 3844 5185
rect 4068 5176 4120 5228
rect 2872 5108 2924 5160
rect 1860 5083 1912 5092
rect 1860 5049 1869 5083
rect 1869 5049 1903 5083
rect 1903 5049 1912 5083
rect 1860 5040 1912 5049
rect 2228 5083 2280 5092
rect 2228 5049 2237 5083
rect 2237 5049 2271 5083
rect 2271 5049 2280 5083
rect 2228 5040 2280 5049
rect 4620 5040 4672 5092
rect 112 4972 164 5024
rect 1676 4972 1728 5024
rect 3424 4972 3476 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 1860 4768 1912 4820
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 3516 4768 3568 4820
rect 4068 4768 4120 4820
rect 1492 4700 1544 4752
rect 1676 4632 1728 4684
rect 2412 4700 2464 4752
rect 3240 4700 3292 4752
rect 4436 4700 4488 4752
rect 2780 4632 2832 4684
rect 4160 4564 4212 4616
rect 4620 4428 4672 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1676 4224 1728 4276
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 1492 4088 1544 4140
rect 3332 4088 3384 4140
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 1768 3995 1820 4004
rect 1768 3961 1777 3995
rect 1777 3961 1811 3995
rect 1811 3961 1820 3995
rect 1768 3952 1820 3961
rect 2136 3995 2188 4004
rect 2136 3961 2145 3995
rect 2145 3961 2179 3995
rect 2179 3961 2188 3995
rect 2136 3952 2188 3961
rect 1952 3884 2004 3936
rect 2320 3884 2372 3936
rect 3240 3884 3292 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 1492 3612 1544 3664
rect 2780 3680 2832 3732
rect 3516 3680 3568 3732
rect 4436 3723 4488 3732
rect 4436 3689 4445 3723
rect 4445 3689 4479 3723
rect 4479 3689 4488 3723
rect 4436 3680 4488 3689
rect 2320 3655 2372 3664
rect 2320 3621 2329 3655
rect 2329 3621 2363 3655
rect 2363 3621 2372 3655
rect 2320 3612 2372 3621
rect 2412 3612 2464 3664
rect 3056 3612 3108 3664
rect 1768 3544 1820 3596
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 4436 3136 4488 3188
rect 4620 3136 4672 3188
rect 2964 3068 3016 3120
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 1676 2932 1728 2984
rect 2780 2975 2832 2984
rect 2780 2941 2789 2975
rect 2789 2941 2823 2975
rect 2823 2941 2832 2975
rect 2780 2932 2832 2941
rect 3056 2975 3108 2984
rect 3056 2941 3065 2975
rect 3065 2941 3099 2975
rect 3099 2941 3108 2975
rect 3056 2932 3108 2941
rect 4620 2932 4672 2984
rect 4344 2864 4396 2916
rect 5264 2864 5316 2916
rect 4436 2796 4488 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2780 2592 2832 2644
rect 4528 2592 4580 2644
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 2136 2456 2188 2508
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 4068 2320 4120 2372
rect 4436 2320 4488 2372
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 2778 27554 2834 28000
rect 2778 27526 2912 27554
rect 2778 27520 2834 27526
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1688 7342 1716 7686
rect 1780 7342 1808 8230
rect 1964 7886 1992 8298
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 8022 2360 8230
rect 2502 8120 2558 8129
rect 2884 8090 2912 27526
rect 8298 27520 8354 28000
rect 13910 27520 13966 28000
rect 19522 27520 19578 28000
rect 25134 27520 25190 28000
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 2502 8055 2558 8064
rect 2872 8084 2924 8090
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1504 5234 1532 5850
rect 1688 5250 1716 7278
rect 1964 7206 1992 7822
rect 2332 7546 2360 7958
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2516 7342 2544 8055
rect 2872 8026 2924 8032
rect 2884 7342 2912 8026
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7342 4200 7686
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 2148 6866 2176 7278
rect 2516 6866 2544 7278
rect 2884 6866 2912 7278
rect 3988 6934 4016 7278
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4448 7002 4476 7210
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 1964 6254 1992 6802
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1768 5296 1820 5302
rect 1688 5244 1768 5250
rect 1688 5238 1820 5244
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1688 5222 1808 5238
rect 110 5128 166 5137
rect 110 5063 166 5072
rect 124 5030 152 5063
rect 112 5024 164 5030
rect 112 4966 164 4972
rect 1504 4758 1532 5170
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1492 4752 1544 4758
rect 1492 4694 1544 4700
rect 1504 4146 1532 4694
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1504 3670 1532 4082
rect 1596 4078 1624 5102
rect 1688 5030 1716 5222
rect 1872 5098 1900 5714
rect 1860 5092 1912 5098
rect 1860 5034 1912 5040
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4826 1716 4966
rect 1872 4826 1900 5034
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1688 4690 1716 4762
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4282 1716 4626
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1596 3738 1624 4014
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1492 3664 1544 3670
rect 1492 3606 1544 3612
rect 1688 3194 1716 4218
rect 1872 4154 1900 4762
rect 1780 4126 1900 4154
rect 1780 4010 1808 4126
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 1780 3602 1808 3946
rect 1964 3942 1992 6190
rect 2148 6186 2176 6802
rect 2516 6390 2544 6802
rect 2884 6458 2912 6802
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 2148 5846 2176 6122
rect 2516 5914 2544 6326
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 2884 5370 2912 6394
rect 3528 5914 3556 6734
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6254 3832 6598
rect 4080 6322 4108 6734
rect 4448 6458 4476 6938
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2884 5166 2912 5306
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1688 2990 1716 3130
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1398 82 1454 480
rect 1780 82 1808 3538
rect 2148 2514 2176 3946
rect 2136 2508 2188 2514
rect 2136 2450 2188 2456
rect 2240 2446 2268 5034
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3436 4826 3464 4966
rect 3528 4826 3556 5850
rect 3804 5234 3832 6190
rect 4080 5914 4108 6258
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4080 4826 4108 5170
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 3670 2360 3878
rect 2424 3670 2452 4694
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2792 4282 2820 4626
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2792 2990 2820 3674
rect 2976 3126 3004 4014
rect 3252 3942 3280 4694
rect 3436 4154 3464 4762
rect 3344 4146 3464 4154
rect 3332 4140 3464 4146
rect 3384 4126 3464 4140
rect 3332 4082 3384 4088
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 3068 2990 3096 3606
rect 3344 3602 3372 4082
rect 3528 3738 3556 4762
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 4172 3058 4200 4558
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2792 2650 2820 2926
rect 4356 2922 4384 6054
rect 4448 4758 4476 6394
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4448 3738 4476 4694
rect 4632 4486 4660 5034
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 3942 4660 4422
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4448 3194 4476 3674
rect 4632 3194 4660 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4448 2854 4476 3130
rect 4632 2990 4660 3130
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 4448 2632 4476 2790
rect 5276 2650 5304 2858
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 4528 2644 4580 2650
rect 4448 2604 4528 2632
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 4448 2378 4476 2604
rect 4528 2586 4580 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 1398 54 1808 82
rect 4080 82 4108 2314
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 4158 82 4214 480
rect 4080 54 4214 82
rect 1398 0 1454 54
rect 4158 0 4214 54
rect 6918 0 6974 480
rect 9770 0 9826 480
rect 12530 0 12586 480
rect 15382 0 15438 480
rect 18142 0 18198 480
rect 20902 0 20958 480
rect 23754 0 23810 480
rect 26514 0 26570 480
<< via2 >>
rect 2502 8064 2558 8120
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 110 5072 166 5128
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
<< metal3 >>
rect 0 26120 480 26240
rect 27520 25848 28000 25968
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22584 480 22704
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 27520 21904 28000 22024
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19048 480 19168
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 27520 17824 28000 17944
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 10277 15808 10597 15809
rect 0 15648 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 27520 13880 28000 14000
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 0 12112 480 12232
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9920
rect 24277 9759 24597 9760
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 5610 8736 5930 8737
rect 0 8576 480 8696
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 62 8122 122 8576
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 2497 8122 2563 8125
rect 62 8120 2563 8122
rect 62 8064 2502 8120
rect 2558 8064 2563 8120
rect 62 8062 2563 8064
rect 2497 8059 2563 8062
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 27520 5856 28000 5976
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5128 480 5160
rect 0 5072 110 5128
rect 166 5072 480 5128
rect 0 5040 480 5072
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 27520 1912 28000 2032
rect 0 1640 480 1760
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__11__C tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 1050 592
use scs8hd_nor4_4  _11_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__C
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_44
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__11__B
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_52
timestamp 1586364061
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_51
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__D
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_61
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_56
timestamp 1586364061
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_60
timestamp 1586364061
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_and4_4  _09_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__07__B
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_11
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__B
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 3680 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_22
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_59
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_and4_4  _07_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__08__C
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__D
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__11__D
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_and4_4  _08_
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__06__C
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__08__B
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__07__C
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__08__D
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_72
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_and4_4  _06_
timestamp 1586364061
transform 1 0 1472 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__06__B
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_13
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _04_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _03_
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__03__A
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_8
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__12__D
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_12
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__C
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__C
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _10_
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 1602 592
use scs8hd_inv_8  _05_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__06__D
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_29
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_28
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__B
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__B
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_54
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_nor4_4  _12_
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 1602 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__10__D
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_67
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_nor4_4  _13_
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 1602 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__13__C
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_54
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__D
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_8
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_48
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__13__B
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_8
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_30
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_54
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 1640 480 1760 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 5040 480 5160 6 address[1]
port 1 nsew default input
rlabel metal2 s 2778 27520 2834 28000 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 8576 480 8696 6 address[3]
port 3 nsew default input
rlabel metal2 s 4158 0 4214 480 6 data_in
port 4 nsew default input
rlabel metal2 s 1398 0 1454 480 6 enable
port 5 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 gfpga_pad_GPIO_PAD[0]
port 6 nsew default bidirectional
rlabel metal2 s 8298 27520 8354 28000 6 gfpga_pad_GPIO_PAD[1]
port 7 nsew default bidirectional
rlabel metal3 s 27520 5856 28000 5976 6 gfpga_pad_GPIO_PAD[2]
port 8 nsew default bidirectional
rlabel metal2 s 6918 0 6974 480 6 gfpga_pad_GPIO_PAD[3]
port 9 nsew default bidirectional
rlabel metal3 s 27520 9800 28000 9920 6 gfpga_pad_GPIO_PAD[4]
port 10 nsew default bidirectional
rlabel metal3 s 0 12112 480 12232 6 gfpga_pad_GPIO_PAD[5]
port 11 nsew default bidirectional
rlabel metal2 s 9770 0 9826 480 6 gfpga_pad_GPIO_PAD[6]
port 12 nsew default bidirectional
rlabel metal2 s 12530 0 12586 480 6 gfpga_pad_GPIO_PAD[7]
port 13 nsew default bidirectional
rlabel metal2 s 15382 0 15438 480 6 right_width_0_height_0__pin_0_
port 14 nsew default input
rlabel metal3 s 0 22584 480 22704 6 right_width_0_height_0__pin_10_
port 15 nsew default input
rlabel metal2 s 19522 27520 19578 28000 6 right_width_0_height_0__pin_11_
port 16 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 right_width_0_height_0__pin_12_
port 17 nsew default input
rlabel metal3 s 0 26120 480 26240 6 right_width_0_height_0__pin_13_
port 18 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 right_width_0_height_0__pin_14_
port 19 nsew default input
rlabel metal2 s 25134 27520 25190 28000 6 right_width_0_height_0__pin_15_
port 20 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 right_width_0_height_0__pin_1_
port 21 nsew default tristate
rlabel metal3 s 27520 13880 28000 14000 6 right_width_0_height_0__pin_2_
port 22 nsew default input
rlabel metal3 s 0 15648 480 15768 6 right_width_0_height_0__pin_3_
port 23 nsew default tristate
rlabel metal2 s 13910 27520 13966 28000 6 right_width_0_height_0__pin_4_
port 24 nsew default input
rlabel metal3 s 0 19048 480 19168 6 right_width_0_height_0__pin_5_
port 25 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 right_width_0_height_0__pin_6_
port 26 nsew default input
rlabel metal2 s 20902 0 20958 480 6 right_width_0_height_0__pin_7_
port 27 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 right_width_0_height_0__pin_8_
port 28 nsew default input
rlabel metal3 s 27520 21904 28000 22024 6 right_width_0_height_0__pin_9_
port 29 nsew default tristate
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 30 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 31 nsew default input
<< end >>
