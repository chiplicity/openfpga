VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_3__3_
  CLASS BLOCK ;
  FOREIGN sb_3__3_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 137.935 BY 137.320 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 2.400 ;
    END
  END address[5]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN bottom_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 2.400 ;
    END
  END bottom_right_grid_pin_13_
  PIN bottom_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END bottom_right_grid_pin_15_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.400 ;
    END
  END bottom_right_grid_pin_1_
  PIN bottom_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END bottom_right_grid_pin_3_
  PIN bottom_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END bottom_right_grid_pin_5_
  PIN bottom_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 2.400 ;
    END
  END bottom_right_grid_pin_7_
  PIN bottom_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 2.400 ;
    END
  END bottom_right_grid_pin_9_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_left_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 2.400 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END left_top_grid_pin_11_
  PIN left_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 2.400 131.880 ;
    END
  END left_top_grid_pin_13_
  PIN left_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 2.400 137.320 ;
    END
  END left_top_grid_pin_15_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END left_top_grid_pin_1_
  PIN left_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END left_top_grid_pin_3_
  PIN left_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END left_top_grid_pin_5_
  PIN left_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END left_top_grid_pin_7_
  PIN left_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END left_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 1.910 2.760 134.320 128.080 ;
      LAYER met2 ;
        RECT 1.940 2.680 137.910 137.205 ;
        RECT 2.490 2.195 5.330 2.680 ;
        RECT 6.170 2.195 9.470 2.680 ;
        RECT 10.310 2.195 13.610 2.680 ;
        RECT 14.450 2.195 17.290 2.680 ;
        RECT 18.130 2.195 21.430 2.680 ;
        RECT 22.270 2.195 25.570 2.680 ;
        RECT 26.410 2.195 29.250 2.680 ;
        RECT 30.090 2.195 33.390 2.680 ;
        RECT 34.230 2.195 37.530 2.680 ;
        RECT 38.370 2.195 41.210 2.680 ;
        RECT 42.050 2.195 45.350 2.680 ;
        RECT 46.190 2.195 49.490 2.680 ;
        RECT 50.330 2.195 53.170 2.680 ;
        RECT 54.010 2.195 57.310 2.680 ;
        RECT 58.150 2.195 61.450 2.680 ;
        RECT 62.290 2.195 65.130 2.680 ;
        RECT 65.970 2.195 69.270 2.680 ;
        RECT 70.110 2.195 73.410 2.680 ;
        RECT 74.250 2.195 77.550 2.680 ;
        RECT 78.390 2.195 81.230 2.680 ;
        RECT 82.070 2.195 85.370 2.680 ;
        RECT 86.210 2.195 89.510 2.680 ;
        RECT 90.350 2.195 93.190 2.680 ;
        RECT 94.030 2.195 97.330 2.680 ;
        RECT 98.170 2.195 101.470 2.680 ;
        RECT 102.310 2.195 105.150 2.680 ;
        RECT 105.990 2.195 109.290 2.680 ;
        RECT 110.130 2.195 113.430 2.680 ;
        RECT 114.270 2.195 117.110 2.680 ;
        RECT 117.950 2.195 121.250 2.680 ;
        RECT 122.090 2.195 125.390 2.680 ;
        RECT 126.230 2.195 129.070 2.680 ;
        RECT 129.910 2.195 133.210 2.680 ;
        RECT 134.050 2.195 137.350 2.680 ;
      LAYER met3 ;
        RECT 2.800 136.320 137.935 137.185 ;
        RECT 2.400 132.280 137.935 136.320 ;
        RECT 2.800 130.880 137.935 132.280 ;
        RECT 2.400 127.520 137.935 130.880 ;
        RECT 2.800 126.120 137.935 127.520 ;
        RECT 2.400 122.080 137.935 126.120 ;
        RECT 2.800 120.680 137.935 122.080 ;
        RECT 2.400 116.640 137.935 120.680 ;
        RECT 2.800 115.240 137.935 116.640 ;
        RECT 2.400 111.880 137.935 115.240 ;
        RECT 2.800 110.480 137.935 111.880 ;
        RECT 2.400 106.440 137.935 110.480 ;
        RECT 2.800 105.040 137.935 106.440 ;
        RECT 2.400 101.000 137.935 105.040 ;
        RECT 2.800 99.600 137.935 101.000 ;
        RECT 2.400 96.240 137.935 99.600 ;
        RECT 2.800 94.840 137.935 96.240 ;
        RECT 2.400 90.800 137.935 94.840 ;
        RECT 2.800 89.400 137.935 90.800 ;
        RECT 2.400 86.040 137.935 89.400 ;
        RECT 2.800 84.640 137.935 86.040 ;
        RECT 2.400 80.600 137.935 84.640 ;
        RECT 2.800 79.200 137.935 80.600 ;
        RECT 2.400 75.160 137.935 79.200 ;
        RECT 2.800 73.760 137.935 75.160 ;
        RECT 2.400 70.400 137.935 73.760 ;
        RECT 2.800 69.000 137.935 70.400 ;
        RECT 2.400 64.960 137.935 69.000 ;
        RECT 2.800 63.560 137.935 64.960 ;
        RECT 2.400 59.520 137.935 63.560 ;
        RECT 2.800 58.120 137.935 59.520 ;
        RECT 2.400 54.760 137.935 58.120 ;
        RECT 2.800 53.360 137.935 54.760 ;
        RECT 2.400 49.320 137.935 53.360 ;
        RECT 2.800 47.920 137.935 49.320 ;
        RECT 2.400 44.560 137.935 47.920 ;
        RECT 2.800 43.160 137.935 44.560 ;
        RECT 2.400 39.120 137.935 43.160 ;
        RECT 2.800 37.720 137.935 39.120 ;
        RECT 2.400 33.680 137.935 37.720 ;
        RECT 2.800 32.280 137.935 33.680 ;
        RECT 2.400 28.920 137.935 32.280 ;
        RECT 2.800 27.520 137.935 28.920 ;
        RECT 2.400 23.480 137.935 27.520 ;
        RECT 2.800 22.080 137.935 23.480 ;
        RECT 2.400 18.040 137.935 22.080 ;
        RECT 2.800 16.640 137.935 18.040 ;
        RECT 2.400 13.280 137.935 16.640 ;
        RECT 2.800 11.880 137.935 13.280 ;
        RECT 2.400 7.840 137.935 11.880 ;
        RECT 2.800 6.440 137.935 7.840 ;
        RECT 2.400 3.080 137.935 6.440 ;
        RECT 2.800 2.215 137.935 3.080 ;
      LAYER met4 ;
        RECT 7.655 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
      LAYER met5 ;
        RECT 30.020 17.900 113.500 19.500 ;
  END
END sb_3__3_
END LIBRARY

