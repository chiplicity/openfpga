magic
tech EFS8A
magscale 1 2
timestamp 1604399453
<< locali >>
rect 13093 12631 13127 12869
rect 16037 12631 16071 12937
rect 23121 11067 23155 11305
rect 11621 9367 11655 9537
rect 24501 9367 24535 9537
rect 14657 8279 14691 8381
rect 7849 6103 7883 6205
rect 24041 5151 24075 5253
rect 12817 3927 12851 4233
rect 15945 3995 15979 4233
rect 20453 3927 20487 4029
rect 6193 3383 6227 3553
rect 14473 2975 14507 3145
<< viali >>
rect 1593 23273 1627 23307
rect 24777 23273 24811 23307
rect 1409 23137 1443 23171
rect 24593 23137 24627 23171
rect 23857 22729 23891 22763
rect 24685 22729 24719 22763
rect 23673 22525 23707 22559
rect 24133 22525 24167 22559
rect 1685 22389 1719 22423
rect 24593 22049 24627 22083
rect 24777 21913 24811 21947
rect 24593 21301 24627 21335
rect 24777 21097 24811 21131
rect 24593 20961 24627 20995
rect 1593 20553 1627 20587
rect 2697 20553 2731 20587
rect 13369 20417 13403 20451
rect 1409 20349 1443 20383
rect 2513 20349 2547 20383
rect 13461 20349 13495 20383
rect 13728 20349 13762 20383
rect 2053 20213 2087 20247
rect 3065 20213 3099 20247
rect 14841 20213 14875 20247
rect 24593 20213 24627 20247
rect 1593 20009 1627 20043
rect 2697 20009 2731 20043
rect 1409 19873 1443 19907
rect 2513 19873 2547 19907
rect 13461 19669 13495 19703
rect 1409 19261 1443 19295
rect 13461 19261 13495 19295
rect 13728 19193 13762 19227
rect 1593 19125 1627 19159
rect 2053 19125 2087 19159
rect 2605 19125 2639 19159
rect 13369 19125 13403 19159
rect 14841 19125 14875 19159
rect 12357 18921 12391 18955
rect 12265 18785 12299 18819
rect 12725 18785 12759 18819
rect 1685 18717 1719 18751
rect 12817 18717 12851 18751
rect 13001 18717 13035 18751
rect 13921 18717 13955 18751
rect 10425 18581 10459 18615
rect 13553 18581 13587 18615
rect 1593 18377 1627 18411
rect 11529 18377 11563 18411
rect 10333 18309 10367 18343
rect 12265 18309 12299 18343
rect 10977 18241 11011 18275
rect 1409 18173 1443 18207
rect 12449 18173 12483 18207
rect 10793 18105 10827 18139
rect 12716 18105 12750 18139
rect 2053 18037 2087 18071
rect 10149 18037 10183 18071
rect 10701 18037 10735 18071
rect 11805 18037 11839 18071
rect 13829 18037 13863 18071
rect 1593 17833 1627 17867
rect 9321 17833 9355 17867
rect 12449 17833 12483 17867
rect 13553 17833 13587 17867
rect 14657 17833 14691 17867
rect 24777 17833 24811 17867
rect 13001 17765 13035 17799
rect 1409 17697 1443 17731
rect 11325 17697 11359 17731
rect 13921 17697 13955 17731
rect 24593 17697 24627 17731
rect 11069 17629 11103 17663
rect 14013 17629 14047 17663
rect 14105 17629 14139 17663
rect 10333 17493 10367 17527
rect 10885 17493 10919 17527
rect 13369 17493 13403 17527
rect 1593 17289 1627 17323
rect 2329 17289 2363 17323
rect 10333 17289 10367 17323
rect 12449 17289 12483 17323
rect 24777 17289 24811 17323
rect 11897 17221 11931 17255
rect 9137 17153 9171 17187
rect 9781 17153 9815 17187
rect 11345 17153 11379 17187
rect 13001 17153 13035 17187
rect 14657 17153 14691 17187
rect 1409 17085 1443 17119
rect 9597 17085 9631 17119
rect 11161 17085 11195 17119
rect 13553 17085 13587 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 10609 17017 10643 17051
rect 11253 17017 11287 17051
rect 12817 17017 12851 17051
rect 13921 17017 13955 17051
rect 14473 17017 14507 17051
rect 15577 17017 15611 17051
rect 2053 16949 2087 16983
rect 9229 16949 9263 16983
rect 9689 16949 9723 16983
rect 10793 16949 10827 16983
rect 12173 16949 12207 16983
rect 12909 16949 12943 16983
rect 14013 16949 14047 16983
rect 14381 16949 14415 16983
rect 15117 16949 15151 16983
rect 24409 16949 24443 16983
rect 1593 16745 1627 16779
rect 9321 16745 9355 16779
rect 10425 16745 10459 16779
rect 11897 16745 11931 16779
rect 12541 16745 12575 16779
rect 13553 16745 13587 16779
rect 14105 16745 14139 16779
rect 15025 16745 15059 16779
rect 23765 16745 23799 16779
rect 24777 16745 24811 16779
rect 10762 16677 10796 16711
rect 12909 16677 12943 16711
rect 14013 16677 14047 16711
rect 15546 16677 15580 16711
rect 1409 16609 1443 16643
rect 10517 16609 10551 16643
rect 23581 16609 23615 16643
rect 24593 16609 24627 16643
rect 14289 16541 14323 16575
rect 15301 16541 15335 16575
rect 8861 16405 8895 16439
rect 13645 16405 13679 16439
rect 16681 16405 16715 16439
rect 2697 16201 2731 16235
rect 8769 16201 8803 16235
rect 10149 16201 10183 16235
rect 11437 16201 11471 16235
rect 13277 16201 13311 16235
rect 14381 16201 14415 16235
rect 24685 16201 24719 16235
rect 1593 16133 1627 16167
rect 23857 16133 23891 16167
rect 8309 16065 8343 16099
rect 9321 16065 9355 16099
rect 10885 16065 10919 16099
rect 13829 16065 13863 16099
rect 14013 16065 14047 16099
rect 1409 15997 1443 16031
rect 2505 15997 2539 16031
rect 9229 15997 9263 16031
rect 9873 15997 9907 16031
rect 10793 15997 10827 16031
rect 12265 15997 12299 16031
rect 13737 15997 13771 16031
rect 14933 15997 14967 16031
rect 15200 15997 15234 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 2329 15929 2363 15963
rect 3065 15929 3099 15963
rect 10701 15929 10735 15963
rect 11713 15929 11747 15963
rect 12909 15929 12943 15963
rect 16865 15929 16899 15963
rect 1961 15861 1995 15895
rect 8585 15861 8619 15895
rect 9137 15861 9171 15895
rect 10333 15861 10367 15895
rect 13369 15861 13403 15895
rect 14749 15861 14783 15895
rect 16313 15861 16347 15895
rect 18245 15861 18279 15895
rect 22569 15861 22603 15895
rect 24225 15861 24259 15895
rect 1593 15657 1627 15691
rect 8493 15657 8527 15691
rect 10609 15657 10643 15691
rect 13093 15657 13127 15691
rect 14105 15657 14139 15691
rect 15301 15657 15335 15691
rect 15669 15657 15703 15691
rect 24777 15657 24811 15691
rect 14013 15589 14047 15623
rect 15761 15589 15795 15623
rect 1409 15521 1443 15555
rect 2605 15521 2639 15555
rect 6837 15521 6871 15555
rect 8401 15521 8435 15555
rect 10793 15521 10827 15555
rect 11060 15521 11094 15555
rect 13461 15521 13495 15555
rect 14749 15521 14783 15555
rect 16865 15521 16899 15555
rect 18429 15521 18463 15555
rect 19441 15521 19475 15555
rect 23581 15521 23615 15555
rect 24593 15521 24627 15555
rect 6929 15453 6963 15487
rect 7113 15453 7147 15487
rect 8585 15453 8619 15487
rect 14289 15453 14323 15487
rect 15025 15453 15059 15487
rect 15853 15453 15887 15487
rect 22569 15453 22603 15487
rect 6469 15385 6503 15419
rect 13645 15385 13679 15419
rect 2789 15317 2823 15351
rect 4261 15317 4295 15351
rect 8033 15317 8067 15351
rect 12173 15317 12207 15351
rect 16405 15317 16439 15351
rect 16773 15317 16807 15351
rect 17049 15317 17083 15351
rect 18613 15317 18647 15351
rect 19625 15317 19659 15351
rect 23765 15317 23799 15351
rect 2053 15113 2087 15147
rect 2513 15113 2547 15147
rect 2789 15113 2823 15147
rect 3893 15113 3927 15147
rect 7113 15113 7147 15147
rect 10333 15113 10367 15147
rect 10793 15113 10827 15147
rect 13001 15113 13035 15147
rect 13369 15113 13403 15147
rect 15853 15113 15887 15147
rect 24777 15113 24811 15147
rect 22293 15045 22327 15079
rect 3801 14977 3835 15011
rect 4445 14977 4479 15011
rect 6561 14977 6595 15011
rect 11345 14977 11379 15011
rect 16865 14977 16899 15011
rect 19993 14977 20027 15011
rect 1869 14909 1903 14943
rect 4261 14909 4295 14943
rect 7941 14909 7975 14943
rect 13829 14909 13863 14943
rect 16773 14909 16807 14943
rect 19165 14909 19199 14943
rect 19625 14909 19659 14943
rect 20177 14909 20211 14943
rect 22109 14909 22143 14943
rect 24409 14909 24443 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 4353 14841 4387 14875
rect 6193 14841 6227 14875
rect 7757 14841 7791 14875
rect 8186 14841 8220 14875
rect 9965 14841 9999 14875
rect 11161 14841 11195 14875
rect 12449 14841 12483 14875
rect 14096 14841 14130 14875
rect 16221 14841 16255 14875
rect 16681 14841 16715 14875
rect 20637 14841 20671 14875
rect 1685 14773 1719 14807
rect 3341 14773 3375 14807
rect 7389 14773 7423 14807
rect 9321 14773 9355 14807
rect 10701 14773 10735 14807
rect 11253 14773 11287 14807
rect 11805 14773 11839 14807
rect 13645 14773 13679 14807
rect 15209 14773 15243 14807
rect 16313 14773 16347 14807
rect 17325 14773 17359 14807
rect 18061 14773 18095 14807
rect 18521 14773 18555 14807
rect 19349 14773 19383 14807
rect 20361 14773 20395 14807
rect 22661 14773 22695 14807
rect 23857 14773 23891 14807
rect 1593 14569 1627 14603
rect 2697 14569 2731 14603
rect 4077 14569 4111 14603
rect 8033 14569 8067 14603
rect 8401 14569 8435 14603
rect 8677 14569 8711 14603
rect 11621 14569 11655 14603
rect 13553 14569 13587 14603
rect 13921 14569 13955 14603
rect 15301 14569 15335 14603
rect 18613 14569 18647 14603
rect 23765 14569 23799 14603
rect 24777 14569 24811 14603
rect 3893 14501 3927 14535
rect 4537 14501 4571 14535
rect 5886 14501 5920 14535
rect 15669 14501 15703 14535
rect 15761 14501 15795 14535
rect 16313 14501 16347 14535
rect 1409 14433 1443 14467
rect 2513 14433 2547 14467
rect 4445 14433 4479 14467
rect 9689 14433 9723 14467
rect 9956 14433 9990 14467
rect 12541 14433 12575 14467
rect 14197 14433 14231 14467
rect 17233 14433 17267 14467
rect 18429 14433 18463 14467
rect 19533 14433 19567 14467
rect 20913 14433 20947 14467
rect 22569 14433 22603 14467
rect 23581 14433 23615 14467
rect 24593 14433 24627 14467
rect 3065 14365 3099 14399
rect 4629 14365 4663 14399
rect 5089 14365 5123 14399
rect 5641 14365 5675 14399
rect 12633 14365 12667 14399
rect 12817 14365 12851 14399
rect 15945 14365 15979 14399
rect 17325 14365 17359 14399
rect 17417 14365 17451 14399
rect 15117 14297 15151 14331
rect 16865 14297 16899 14331
rect 3433 14229 3467 14263
rect 7021 14229 7055 14263
rect 11069 14229 11103 14263
rect 12173 14229 12207 14263
rect 14381 14229 14415 14263
rect 14749 14229 14783 14263
rect 16681 14229 16715 14263
rect 18153 14229 18187 14263
rect 19717 14229 19751 14263
rect 21097 14229 21131 14263
rect 22753 14229 22787 14263
rect 1593 14025 1627 14059
rect 2421 14025 2455 14059
rect 3801 14025 3835 14059
rect 5641 14025 5675 14059
rect 6561 14025 6595 14059
rect 8677 14025 8711 14059
rect 9781 14025 9815 14059
rect 10609 14025 10643 14059
rect 11713 14025 11747 14059
rect 13001 14025 13035 14059
rect 15577 14025 15611 14059
rect 17325 14025 17359 14059
rect 19073 14025 19107 14059
rect 19809 14025 19843 14059
rect 23397 14025 23431 14059
rect 2697 13957 2731 13991
rect 4169 13957 4203 13991
rect 6193 13957 6227 13991
rect 7113 13957 7147 13991
rect 10517 13957 10551 13991
rect 16129 13957 16163 13991
rect 16313 13957 16347 13991
rect 21097 13957 21131 13991
rect 24777 13957 24811 13991
rect 3157 13889 3191 13923
rect 4261 13889 4295 13923
rect 7297 13889 7331 13923
rect 11161 13889 11195 13923
rect 16773 13889 16807 13923
rect 16957 13889 16991 13923
rect 18521 13889 18555 13923
rect 18613 13889 18647 13923
rect 20085 13889 20119 13923
rect 1409 13821 1443 13855
rect 2053 13821 2087 13855
rect 2519 13821 2553 13855
rect 4517 13821 4551 13855
rect 10057 13821 10091 13855
rect 10977 13821 11011 13855
rect 12173 13821 12207 13855
rect 13553 13821 13587 13855
rect 13820 13821 13854 13855
rect 17785 13821 17819 13855
rect 19625 13821 19659 13855
rect 20453 13821 20487 13855
rect 20913 13821 20947 13855
rect 21741 13821 21775 13855
rect 22569 13821 22603 13855
rect 23121 13821 23155 13855
rect 23949 13821 23983 13855
rect 24593 13821 24627 13855
rect 25145 13821 25179 13855
rect 7542 13753 7576 13787
rect 11069 13753 11103 13787
rect 16681 13753 16715 13787
rect 12633 13685 12667 13719
rect 13461 13685 13495 13719
rect 14933 13685 14967 13719
rect 18061 13685 18095 13719
rect 18429 13685 18463 13719
rect 21465 13685 21499 13719
rect 22753 13685 22787 13719
rect 24409 13685 24443 13719
rect 1593 13481 1627 13515
rect 2697 13481 2731 13515
rect 5641 13481 5675 13515
rect 7573 13481 7607 13515
rect 8585 13481 8619 13515
rect 10701 13481 10735 13515
rect 10793 13481 10827 13515
rect 11253 13481 11287 13515
rect 13645 13481 13679 13515
rect 15117 13481 15151 13515
rect 15577 13481 15611 13515
rect 18153 13481 18187 13515
rect 18705 13481 18739 13515
rect 20085 13481 20119 13515
rect 23765 13481 23799 13515
rect 24777 13481 24811 13515
rect 7389 13413 7423 13447
rect 8033 13413 8067 13447
rect 13553 13413 13587 13447
rect 14657 13413 14691 13447
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 3065 13345 3099 13379
rect 4261 13345 4295 13379
rect 4528 13345 4562 13379
rect 7021 13345 7055 13379
rect 7941 13345 7975 13379
rect 11161 13345 11195 13379
rect 12633 13345 12667 13379
rect 14013 13345 14047 13379
rect 14105 13345 14139 13379
rect 16488 13345 16522 13379
rect 19073 13345 19107 13379
rect 19717 13345 19751 13379
rect 23581 13345 23615 13379
rect 24593 13345 24627 13379
rect 2421 13277 2455 13311
rect 8125 13277 8159 13311
rect 9689 13277 9723 13311
rect 11437 13277 11471 13311
rect 14289 13277 14323 13311
rect 16221 13277 16255 13311
rect 19165 13277 19199 13311
rect 19257 13277 19291 13311
rect 20913 13277 20947 13311
rect 22569 13277 22603 13311
rect 1961 13209 1995 13243
rect 3525 13141 3559 13175
rect 3801 13141 3835 13175
rect 12817 13141 12851 13175
rect 13093 13141 13127 13175
rect 16129 13141 16163 13175
rect 17601 13141 17635 13175
rect 18521 13141 18555 13175
rect 1593 12937 1627 12971
rect 1961 12937 1995 12971
rect 3157 12937 3191 12971
rect 4261 12937 4295 12971
rect 6653 12937 6687 12971
rect 8217 12937 8251 12971
rect 11253 12937 11287 12971
rect 11805 12937 11839 12971
rect 13829 12937 13863 12971
rect 16037 12937 16071 12971
rect 16129 12937 16163 12971
rect 16313 12937 16347 12971
rect 23857 12937 23891 12971
rect 24777 12937 24811 12971
rect 4721 12869 4755 12903
rect 7389 12869 7423 12903
rect 10793 12869 10827 12903
rect 13093 12869 13127 12903
rect 3617 12801 3651 12835
rect 3709 12801 3743 12835
rect 5273 12801 5307 12835
rect 5733 12801 5767 12835
rect 8769 12801 8803 12835
rect 10333 12801 10367 12835
rect 1409 12733 1443 12767
rect 3065 12733 3099 12767
rect 4629 12733 4663 12767
rect 5089 12733 5123 12767
rect 7757 12733 7791 12767
rect 8585 12733 8619 12767
rect 9321 12733 9355 12767
rect 11345 12733 11379 12767
rect 12817 12733 12851 12767
rect 3525 12665 3559 12699
rect 5181 12665 5215 12699
rect 8125 12665 8159 12699
rect 8677 12665 8711 12699
rect 9689 12665 9723 12699
rect 10149 12665 10183 12699
rect 12725 12665 12759 12699
rect 14381 12801 14415 12835
rect 14933 12801 14967 12835
rect 15485 12801 15519 12835
rect 13737 12733 13771 12767
rect 14197 12733 14231 12767
rect 18061 12869 18095 12903
rect 19625 12869 19659 12903
rect 22753 12869 22787 12903
rect 24409 12869 24443 12903
rect 16957 12801 16991 12835
rect 17325 12801 17359 12835
rect 18613 12801 18647 12835
rect 19073 12801 19107 12835
rect 20085 12801 20119 12835
rect 20177 12801 20211 12835
rect 16681 12733 16715 12767
rect 19993 12733 20027 12767
rect 22561 12733 22595 12767
rect 24593 12733 24627 12767
rect 25145 12733 25179 12767
rect 17785 12665 17819 12699
rect 18429 12665 18463 12699
rect 18521 12665 18555 12699
rect 19533 12665 19567 12699
rect 23029 12665 23063 12699
rect 2513 12597 2547 12631
rect 9781 12597 9815 12631
rect 10241 12597 10275 12631
rect 11529 12597 11563 12631
rect 12265 12597 12299 12631
rect 13001 12597 13035 12631
rect 13093 12597 13127 12631
rect 13277 12597 13311 12631
rect 14289 12597 14323 12631
rect 15853 12597 15887 12631
rect 16037 12597 16071 12631
rect 16773 12597 16807 12631
rect 20729 12597 20763 12631
rect 21189 12597 21223 12631
rect 1593 12393 1627 12427
rect 2421 12393 2455 12427
rect 4261 12393 4295 12427
rect 7757 12393 7791 12427
rect 14197 12393 14231 12427
rect 15301 12393 15335 12427
rect 16129 12393 16163 12427
rect 16589 12393 16623 12427
rect 19625 12393 19659 12427
rect 20269 12393 20303 12427
rect 24777 12393 24811 12427
rect 2789 12325 2823 12359
rect 5641 12325 5675 12359
rect 14933 12325 14967 12359
rect 1409 12257 1443 12291
rect 5733 12257 5767 12291
rect 7297 12257 7331 12291
rect 8125 12257 8159 12291
rect 10517 12257 10551 12291
rect 10773 12257 10807 12291
rect 13553 12257 13587 12291
rect 17040 12257 17074 12291
rect 19073 12257 19107 12291
rect 19717 12257 19751 12291
rect 21925 12257 21959 12291
rect 22181 12257 22215 12291
rect 24593 12257 24627 12291
rect 2881 12189 2915 12223
rect 2973 12189 3007 12223
rect 5089 12189 5123 12223
rect 5825 12189 5859 12223
rect 7665 12189 7699 12223
rect 8217 12189 8251 12223
rect 8401 12189 8435 12223
rect 13645 12189 13679 12223
rect 13829 12189 13863 12223
rect 14565 12189 14599 12223
rect 16773 12189 16807 12223
rect 19809 12189 19843 12223
rect 20913 12189 20947 12223
rect 3801 12121 3835 12155
rect 5273 12121 5307 12155
rect 9873 12121 9907 12155
rect 11897 12121 11931 12155
rect 13001 12121 13035 12155
rect 1869 12053 1903 12087
rect 2329 12053 2363 12087
rect 3433 12053 3467 12087
rect 4813 12053 4847 12087
rect 6285 12053 6319 12087
rect 6653 12053 6687 12087
rect 13185 12053 13219 12087
rect 18153 12053 18187 12087
rect 18705 12053 18739 12087
rect 19257 12053 19291 12087
rect 21373 12053 21407 12087
rect 21833 12053 21867 12087
rect 23305 12053 23339 12087
rect 23949 12053 23983 12087
rect 1777 11849 1811 11883
rect 3341 11849 3375 11883
rect 5181 11849 5215 11883
rect 6469 11849 6503 11883
rect 7113 11849 7147 11883
rect 9229 11849 9263 11883
rect 9689 11849 9723 11883
rect 10793 11849 10827 11883
rect 11897 11849 11931 11883
rect 13277 11849 13311 11883
rect 16129 11849 16163 11883
rect 17509 11849 17543 11883
rect 22845 11849 22879 11883
rect 23397 11849 23431 11883
rect 18797 11781 18831 11815
rect 2789 11713 2823 11747
rect 7297 11713 7331 11747
rect 11437 11713 11471 11747
rect 16589 11713 16623 11747
rect 16773 11713 16807 11747
rect 22385 11713 22419 11747
rect 3709 11645 3743 11679
rect 3801 11645 3835 11679
rect 7564 11645 7598 11679
rect 9781 11645 9815 11679
rect 12449 11645 12483 11679
rect 13645 11645 13679 11679
rect 13912 11645 13946 11679
rect 15669 11645 15703 11679
rect 19165 11645 19199 11679
rect 19349 11645 19383 11679
rect 22201 11645 22235 11679
rect 23673 11645 23707 11679
rect 2697 11577 2731 11611
rect 4046 11577 4080 11611
rect 5825 11577 5859 11611
rect 10701 11577 10735 11611
rect 11161 11577 11195 11611
rect 19594 11577 19628 11611
rect 21649 11577 21683 11611
rect 23940 11577 23974 11611
rect 2053 11509 2087 11543
rect 2237 11509 2271 11543
rect 2605 11509 2639 11543
rect 6193 11509 6227 11543
rect 8677 11509 8711 11543
rect 9965 11509 9999 11543
rect 10241 11509 10275 11543
rect 11253 11509 11287 11543
rect 15025 11509 15059 11543
rect 16037 11509 16071 11543
rect 16497 11509 16531 11543
rect 17233 11509 17267 11543
rect 18061 11509 18095 11543
rect 20729 11509 20763 11543
rect 21281 11509 21315 11543
rect 21833 11509 21867 11543
rect 22293 11509 22327 11543
rect 25053 11509 25087 11543
rect 1593 11305 1627 11339
rect 2421 11305 2455 11339
rect 4077 11305 4111 11339
rect 4445 11305 4479 11339
rect 7389 11305 7423 11339
rect 7941 11305 7975 11339
rect 12081 11305 12115 11339
rect 13093 11305 13127 11339
rect 13185 11305 13219 11339
rect 14657 11305 14691 11339
rect 16681 11305 16715 11339
rect 18705 11305 18739 11339
rect 19257 11305 19291 11339
rect 20729 11305 20763 11339
rect 22845 11305 22879 11339
rect 23121 11305 23155 11339
rect 23857 11305 23891 11339
rect 25145 11305 25179 11339
rect 4537 11237 4571 11271
rect 7665 11237 7699 11271
rect 8309 11237 8343 11271
rect 13645 11237 13679 11271
rect 1409 11169 1443 11203
rect 1961 11169 1995 11203
rect 2789 11169 2823 11203
rect 6009 11169 6043 11203
rect 10609 11169 10643 11203
rect 10701 11169 10735 11203
rect 10968 11169 11002 11203
rect 13553 11169 13587 11203
rect 15568 11169 15602 11203
rect 19625 11169 19659 11203
rect 19717 11169 19751 11203
rect 21169 11169 21203 11203
rect 2881 11101 2915 11135
rect 2973 11101 3007 11135
rect 4629 11101 4663 11135
rect 6101 11101 6135 11135
rect 6285 11101 6319 11135
rect 8401 11101 8435 11135
rect 8493 11101 8527 11135
rect 9689 11101 9723 11135
rect 13829 11101 13863 11135
rect 14289 11101 14323 11135
rect 15301 11101 15335 11135
rect 18153 11101 18187 11135
rect 19901 11101 19935 11135
rect 20913 11101 20947 11135
rect 23765 11169 23799 11203
rect 24961 11169 24995 11203
rect 23949 11101 23983 11135
rect 2237 11033 2271 11067
rect 3433 11033 3467 11067
rect 3893 11033 3927 11067
rect 5641 11033 5675 11067
rect 6653 11033 6687 11067
rect 10149 11033 10183 11067
rect 20361 11033 20395 11067
rect 22293 11033 22327 11067
rect 23121 11033 23155 11067
rect 23213 11033 23247 11067
rect 24593 11033 24627 11067
rect 5089 10965 5123 10999
rect 5457 10965 5491 10999
rect 12725 10965 12759 10999
rect 18061 10965 18095 10999
rect 19165 10965 19199 10999
rect 23397 10965 23431 10999
rect 1593 10761 1627 10795
rect 3985 10761 4019 10795
rect 4629 10761 4663 10795
rect 5089 10761 5123 10795
rect 7573 10761 7607 10795
rect 11437 10761 11471 10795
rect 13461 10761 13495 10795
rect 14197 10761 14231 10795
rect 15025 10761 15059 10795
rect 15393 10761 15427 10795
rect 16865 10761 16899 10795
rect 20085 10761 20119 10795
rect 20637 10761 20671 10795
rect 22661 10761 22695 10795
rect 24961 10761 24995 10795
rect 25421 10761 25455 10795
rect 7205 10693 7239 10727
rect 10333 10693 10367 10727
rect 12449 10693 12483 10727
rect 20545 10693 20579 10727
rect 23489 10693 23523 10727
rect 5549 10625 5583 10659
rect 5733 10625 5767 10659
rect 7665 10625 7699 10659
rect 10241 10625 10275 10659
rect 10885 10625 10919 10659
rect 12265 10625 12299 10659
rect 13001 10625 13035 10659
rect 15485 10625 15519 10659
rect 21097 10625 21131 10659
rect 21189 10625 21223 10659
rect 24317 10625 24351 10659
rect 1409 10557 1443 10591
rect 2513 10557 2547 10591
rect 2605 10557 2639 10591
rect 7932 10557 7966 10591
rect 12817 10557 12851 10591
rect 15752 10557 15786 10591
rect 18153 10557 18187 10591
rect 21005 10557 21039 10591
rect 22477 10557 22511 10591
rect 23029 10557 23063 10591
rect 24041 10557 24075 10591
rect 24133 10557 24167 10591
rect 25237 10557 25271 10591
rect 25789 10557 25823 10591
rect 2872 10489 2906 10523
rect 4997 10489 5031 10523
rect 5457 10489 5491 10523
rect 6193 10489 6227 10523
rect 10793 10489 10827 10523
rect 11805 10489 11839 10523
rect 18398 10489 18432 10523
rect 21649 10489 21683 10523
rect 1961 10421 1995 10455
rect 6561 10421 6595 10455
rect 9045 10421 9079 10455
rect 9781 10421 9815 10455
rect 10701 10421 10735 10455
rect 12909 10421 12943 10455
rect 13921 10421 13955 10455
rect 14473 10421 14507 10455
rect 17417 10421 17451 10455
rect 17877 10421 17911 10455
rect 19533 10421 19567 10455
rect 22017 10421 22051 10455
rect 23673 10421 23707 10455
rect 1593 10217 1627 10251
rect 1961 10217 1995 10251
rect 2421 10217 2455 10251
rect 2789 10217 2823 10251
rect 7573 10217 7607 10251
rect 8585 10217 8619 10251
rect 9505 10217 9539 10251
rect 10057 10217 10091 10251
rect 10977 10217 11011 10251
rect 11621 10217 11655 10251
rect 12725 10217 12759 10251
rect 13185 10217 13219 10251
rect 15761 10217 15795 10251
rect 16129 10217 16163 10251
rect 17141 10217 17175 10251
rect 18245 10217 18279 10251
rect 18613 10217 18647 10251
rect 20545 10217 20579 10251
rect 20913 10217 20947 10251
rect 21281 10217 21315 10251
rect 22109 10217 22143 10251
rect 25145 10217 25179 10251
rect 13093 10149 13127 10183
rect 22753 10149 22787 10183
rect 23121 10149 23155 10183
rect 1409 10081 1443 10115
rect 4804 10081 4838 10115
rect 7941 10081 7975 10115
rect 8033 10081 8067 10115
rect 10149 10081 10183 10115
rect 11529 10081 11563 10115
rect 17049 10081 17083 10115
rect 19349 10081 19383 10115
rect 19809 10081 19843 10115
rect 23213 10081 23247 10115
rect 23480 10081 23514 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 4537 10013 4571 10047
rect 8217 10013 8251 10047
rect 11713 10013 11747 10047
rect 13369 10013 13403 10047
rect 15301 10013 15335 10047
rect 17325 10013 17359 10047
rect 17785 10013 17819 10047
rect 18705 10013 18739 10047
rect 18889 10013 18923 10047
rect 21373 10013 21407 10047
rect 21465 10013 21499 10047
rect 3525 9945 3559 9979
rect 7113 9945 7147 9979
rect 7481 9945 7515 9979
rect 8953 9945 8987 9979
rect 10333 9945 10367 9979
rect 11161 9945 11195 9979
rect 16681 9945 16715 9979
rect 19993 9945 20027 9979
rect 2329 9877 2363 9911
rect 3893 9877 3927 9911
rect 4445 9877 4479 9911
rect 5917 9877 5951 9911
rect 6469 9877 6503 9911
rect 10609 9877 10643 9911
rect 12541 9877 12575 9911
rect 13829 9877 13863 9911
rect 14105 9877 14139 9911
rect 14565 9877 14599 9911
rect 16589 9877 16623 9911
rect 18153 9877 18187 9911
rect 19717 9877 19751 9911
rect 24593 9877 24627 9911
rect 1593 9673 1627 9707
rect 10425 9673 10459 9707
rect 17417 9673 17451 9707
rect 17877 9673 17911 9707
rect 19993 9673 20027 9707
rect 20361 9673 20395 9707
rect 21097 9673 21131 9707
rect 21465 9673 21499 9707
rect 23305 9673 23339 9707
rect 2789 9605 2823 9639
rect 3893 9605 3927 9639
rect 4353 9605 4387 9639
rect 6561 9605 6595 9639
rect 9321 9605 9355 9639
rect 11805 9605 11839 9639
rect 12449 9605 12483 9639
rect 13461 9605 13495 9639
rect 13829 9605 13863 9639
rect 14473 9605 14507 9639
rect 16037 9605 16071 9639
rect 23673 9605 23707 9639
rect 25421 9605 25455 9639
rect 2697 9537 2731 9571
rect 3433 9537 3467 9571
rect 4997 9537 5031 9571
rect 10977 9537 11011 9571
rect 11621 9537 11655 9571
rect 13093 9537 13127 9571
rect 15025 9537 15059 9571
rect 16589 9537 16623 9571
rect 22477 9537 22511 9571
rect 22661 9537 22695 9571
rect 24317 9537 24351 9571
rect 24501 9537 24535 9571
rect 1409 9469 1443 9503
rect 3249 9469 3283 9503
rect 4813 9469 4847 9503
rect 7941 9469 7975 9503
rect 8197 9469 8231 9503
rect 10333 9469 10367 9503
rect 10793 9469 10827 9503
rect 4261 9401 4295 9435
rect 4721 9401 4755 9435
rect 6837 9401 6871 9435
rect 12173 9469 12207 9503
rect 12909 9469 12943 9503
rect 14841 9469 14875 9503
rect 16405 9469 16439 9503
rect 18061 9469 18095 9503
rect 18317 9469 18351 9503
rect 20545 9469 20579 9503
rect 21925 9469 21959 9503
rect 22385 9469 22419 9503
rect 24041 9469 24075 9503
rect 12817 9401 12851 9435
rect 14933 9401 14967 9435
rect 15577 9401 15611 9435
rect 24133 9401 24167 9435
rect 25237 9469 25271 9503
rect 25789 9469 25823 9503
rect 25053 9401 25087 9435
rect 2053 9333 2087 9367
rect 3157 9333 3191 9367
rect 5365 9333 5399 9367
rect 5825 9333 5859 9367
rect 6193 9333 6227 9367
rect 7573 9333 7607 9367
rect 9965 9333 9999 9367
rect 10885 9333 10919 9367
rect 11529 9333 11563 9367
rect 11621 9333 11655 9367
rect 14289 9333 14323 9367
rect 15945 9333 15979 9367
rect 16497 9333 16531 9367
rect 17049 9333 17083 9367
rect 19441 9333 19475 9367
rect 20729 9333 20763 9367
rect 22017 9333 22051 9367
rect 24501 9333 24535 9367
rect 24777 9333 24811 9367
rect 2421 9129 2455 9163
rect 2789 9129 2823 9163
rect 7113 9129 7147 9163
rect 7205 9129 7239 9163
rect 7573 9129 7607 9163
rect 9321 9129 9355 9163
rect 11713 9129 11747 9163
rect 14565 9129 14599 9163
rect 15025 9129 15059 9163
rect 16681 9129 16715 9163
rect 17325 9129 17359 9163
rect 17601 9129 17635 9163
rect 18153 9129 18187 9163
rect 21373 9129 21407 9163
rect 22385 9129 22419 9163
rect 22845 9129 22879 9163
rect 23213 9129 23247 9163
rect 23673 9129 23707 9163
rect 1961 9061 1995 9095
rect 15546 9061 15580 9095
rect 18521 9061 18555 9095
rect 21281 9061 21315 9095
rect 22109 9061 22143 9095
rect 24032 9061 24066 9095
rect 2881 8993 2915 9027
rect 4077 8993 4111 9027
rect 4344 8993 4378 9027
rect 9045 8993 9079 9027
rect 10600 8993 10634 9027
rect 13185 8993 13219 9027
rect 13277 8993 13311 9027
rect 19717 8993 19751 9027
rect 20269 8993 20303 9027
rect 22661 8993 22695 9027
rect 23765 8993 23799 9027
rect 1409 8925 1443 8959
rect 3065 8925 3099 8959
rect 7665 8925 7699 8959
rect 7757 8925 7791 8959
rect 10333 8925 10367 8959
rect 13369 8925 13403 8959
rect 15301 8925 15335 8959
rect 18613 8925 18647 8959
rect 18797 8925 18831 8959
rect 21465 8925 21499 8959
rect 3525 8857 3559 8891
rect 19349 8857 19383 8891
rect 20913 8857 20947 8891
rect 2329 8789 2363 8823
rect 3893 8789 3927 8823
rect 5457 8789 5491 8823
rect 6101 8789 6135 8823
rect 6745 8789 6779 8823
rect 8309 8789 8343 8823
rect 8585 8789 8619 8823
rect 10241 8789 10275 8823
rect 12449 8789 12483 8823
rect 12817 8789 12851 8823
rect 13829 8789 13863 8823
rect 18061 8789 18095 8823
rect 19901 8789 19935 8823
rect 20729 8789 20763 8823
rect 25145 8789 25179 8823
rect 3617 8585 3651 8619
rect 4537 8585 4571 8619
rect 7113 8585 7147 8619
rect 10057 8585 10091 8619
rect 10977 8585 11011 8619
rect 13829 8585 13863 8619
rect 17877 8585 17911 8619
rect 19441 8585 19475 8619
rect 20177 8585 20211 8619
rect 20545 8585 20579 8619
rect 24961 8585 24995 8619
rect 25329 8585 25363 8619
rect 25697 8585 25731 8619
rect 5181 8517 5215 8551
rect 16313 8517 16347 8551
rect 22017 8517 22051 8551
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 7665 8449 7699 8483
rect 10609 8449 10643 8483
rect 11345 8449 11379 8483
rect 11897 8449 11931 8483
rect 23121 8449 23155 8483
rect 24409 8449 24443 8483
rect 24593 8449 24627 8483
rect 2145 8381 2179 8415
rect 2237 8381 2271 8415
rect 5549 8381 5583 8415
rect 8677 8381 8711 8415
rect 8944 8381 8978 8415
rect 12449 8381 12483 8415
rect 12705 8381 12739 8415
rect 14657 8381 14691 8415
rect 14933 8381 14967 8415
rect 17509 8381 17543 8415
rect 18061 8381 18095 8415
rect 20637 8381 20671 8415
rect 25513 8381 25547 8415
rect 26065 8381 26099 8415
rect 2482 8313 2516 8347
rect 4261 8313 4295 8347
rect 5089 8313 5123 8347
rect 5641 8313 5675 8347
rect 6561 8313 6595 8347
rect 7573 8313 7607 8347
rect 8493 8313 8527 8347
rect 12173 8313 12207 8347
rect 14473 8313 14507 8347
rect 15200 8313 15234 8347
rect 17049 8313 17083 8347
rect 18328 8313 18362 8347
rect 20882 8313 20916 8347
rect 22661 8313 22695 8347
rect 23489 8313 23523 8347
rect 24317 8313 24351 8347
rect 1777 8245 1811 8279
rect 7481 8245 7515 8279
rect 8125 8245 8159 8279
rect 14657 8245 14691 8279
rect 14749 8245 14783 8279
rect 23949 8245 23983 8279
rect 2237 8041 2271 8075
rect 3249 8041 3283 8075
rect 4537 8041 4571 8075
rect 5273 8041 5307 8075
rect 5825 8041 5859 8075
rect 7573 8041 7607 8075
rect 10701 8041 10735 8075
rect 11069 8041 11103 8075
rect 12541 8041 12575 8075
rect 13185 8041 13219 8075
rect 13645 8041 13679 8075
rect 14013 8041 14047 8075
rect 15485 8041 15519 8075
rect 16129 8041 16163 8075
rect 17141 8041 17175 8075
rect 17693 8041 17727 8075
rect 18153 8041 18187 8075
rect 18705 8041 18739 8075
rect 19257 8041 19291 8075
rect 19625 8041 19659 8075
rect 20729 8041 20763 8075
rect 22293 8041 22327 8075
rect 23489 8041 23523 8075
rect 2145 7973 2179 8007
rect 10149 7973 10183 8007
rect 11428 7973 11462 8007
rect 24216 7973 24250 8007
rect 2605 7905 2639 7939
rect 4445 7905 4479 7939
rect 6193 7905 6227 7939
rect 6285 7905 6319 7939
rect 8033 7905 8067 7939
rect 14105 7905 14139 7939
rect 16497 7905 16531 7939
rect 16589 7905 16623 7939
rect 18061 7905 18095 7939
rect 19165 7905 19199 7939
rect 20361 7905 20395 7939
rect 21180 7905 21214 7939
rect 2697 7837 2731 7871
rect 2789 7837 2823 7871
rect 4629 7837 4663 7871
rect 6377 7837 6411 7871
rect 8125 7837 8159 7871
rect 8309 7837 8343 7871
rect 11161 7837 11195 7871
rect 14197 7837 14231 7871
rect 16773 7837 16807 7871
rect 17601 7837 17635 7871
rect 18245 7837 18279 7871
rect 19717 7837 19751 7871
rect 19809 7837 19843 7871
rect 20913 7837 20947 7871
rect 23949 7837 23983 7871
rect 4077 7769 4111 7803
rect 5733 7769 5767 7803
rect 8769 7769 8803 7803
rect 9321 7769 9355 7803
rect 16037 7769 16071 7803
rect 1593 7701 1627 7735
rect 3801 7701 3835 7735
rect 7113 7701 7147 7735
rect 7665 7701 7699 7735
rect 9873 7701 9907 7735
rect 13461 7701 13495 7735
rect 14657 7701 14691 7735
rect 15025 7701 15059 7735
rect 22845 7701 22879 7735
rect 23765 7701 23799 7735
rect 25329 7701 25363 7735
rect 2053 7497 2087 7531
rect 4537 7497 4571 7531
rect 8217 7497 8251 7531
rect 10701 7497 10735 7531
rect 11989 7497 12023 7531
rect 13369 7497 13403 7531
rect 16313 7497 16347 7531
rect 17325 7497 17359 7531
rect 17785 7497 17819 7531
rect 20729 7497 20763 7531
rect 21741 7497 21775 7531
rect 23673 7497 23707 7531
rect 25145 7497 25179 7531
rect 5181 7429 5215 7463
rect 6285 7429 6319 7463
rect 8769 7429 8803 7463
rect 9321 7429 9355 7463
rect 11621 7429 11655 7463
rect 13645 7429 13679 7463
rect 15209 7429 15243 7463
rect 19349 7429 19383 7463
rect 23489 7429 23523 7463
rect 2145 7361 2179 7395
rect 4169 7361 4203 7395
rect 5825 7361 5859 7395
rect 9965 7361 9999 7395
rect 11161 7361 11195 7395
rect 13829 7361 13863 7395
rect 16957 7361 16991 7395
rect 18521 7361 18555 7395
rect 18705 7361 18739 7395
rect 21373 7361 21407 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 5549 7293 5583 7327
rect 5641 7293 5675 7327
rect 6837 7293 6871 7327
rect 7093 7293 7127 7327
rect 10333 7293 10367 7327
rect 14096 7293 14130 7327
rect 15853 7293 15887 7327
rect 16681 7293 16715 7327
rect 18429 7293 18463 7327
rect 19625 7293 19659 7327
rect 20177 7293 20211 7327
rect 22109 7293 22143 7327
rect 22477 7293 22511 7327
rect 23121 7293 23155 7327
rect 25237 7293 25271 7327
rect 25789 7293 25823 7327
rect 1685 7225 1719 7259
rect 2390 7225 2424 7259
rect 5089 7225 5123 7259
rect 9781 7225 9815 7259
rect 12725 7225 12759 7259
rect 16129 7225 16163 7259
rect 16773 7225 16807 7259
rect 20545 7225 20579 7259
rect 21097 7225 21131 7259
rect 21189 7225 21223 7259
rect 24041 7225 24075 7259
rect 3525 7157 3559 7191
rect 6561 7157 6595 7191
rect 9137 7157 9171 7191
rect 9689 7157 9723 7191
rect 12817 7157 12851 7191
rect 18061 7157 18095 7191
rect 19809 7157 19843 7191
rect 22661 7157 22695 7191
rect 24685 7157 24719 7191
rect 25421 7157 25455 7191
rect 2329 6953 2363 6987
rect 2421 6953 2455 6987
rect 12173 6953 12207 6987
rect 18061 6953 18095 6987
rect 18889 6953 18923 6987
rect 20269 6953 20303 6987
rect 20729 6953 20763 6987
rect 22293 6953 22327 6987
rect 23213 6953 23247 6987
rect 5724 6885 5758 6919
rect 8309 6885 8343 6919
rect 13185 6885 13219 6919
rect 13737 6885 13771 6919
rect 24032 6885 24066 6919
rect 1409 6817 1443 6851
rect 2789 6817 2823 6851
rect 4077 6817 4111 6851
rect 5273 6817 5307 6851
rect 8401 6817 8435 6851
rect 9781 6817 9815 6851
rect 11060 6817 11094 6851
rect 15025 6817 15059 6851
rect 15577 6817 15611 6851
rect 16293 6817 16327 6851
rect 19993 6817 20027 6851
rect 21169 6817 21203 6851
rect 1961 6749 1995 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 5457 6749 5491 6783
rect 8493 6749 8527 6783
rect 10793 6749 10827 6783
rect 13829 6749 13863 6783
rect 13921 6749 13955 6783
rect 16037 6749 16071 6783
rect 18981 6749 19015 6783
rect 19073 6749 19107 6783
rect 20913 6749 20947 6783
rect 23765 6749 23799 6783
rect 1593 6681 1627 6715
rect 7941 6681 7975 6715
rect 12909 6681 12943 6715
rect 3433 6613 3467 6647
rect 3893 6613 3927 6647
rect 4629 6613 4663 6647
rect 6837 6613 6871 6647
rect 7665 6613 7699 6647
rect 8953 6613 8987 6647
rect 9321 6613 9355 6647
rect 10241 6613 10275 6647
rect 10609 6613 10643 6647
rect 13369 6613 13403 6647
rect 14381 6613 14415 6647
rect 15945 6613 15979 6647
rect 17417 6613 17451 6647
rect 18521 6613 18555 6647
rect 19533 6613 19567 6647
rect 22937 6613 22971 6647
rect 23673 6613 23707 6647
rect 25145 6613 25179 6647
rect 2145 6409 2179 6443
rect 2789 6409 2823 6443
rect 4445 6409 4479 6443
rect 5825 6409 5859 6443
rect 6653 6409 6687 6443
rect 9505 6409 9539 6443
rect 13369 6409 13403 6443
rect 15117 6409 15151 6443
rect 17509 6409 17543 6443
rect 17877 6409 17911 6443
rect 21189 6409 21223 6443
rect 23121 6409 23155 6443
rect 2513 6341 2547 6375
rect 5457 6341 5491 6375
rect 10517 6341 10551 6375
rect 12173 6341 12207 6375
rect 18797 6341 18831 6375
rect 3249 6273 3283 6307
rect 3433 6273 3467 6307
rect 5089 6273 5123 6307
rect 6837 6273 6871 6307
rect 11161 6273 11195 6307
rect 17049 6273 17083 6307
rect 22661 6273 22695 6307
rect 3157 6205 3191 6239
rect 3985 6205 4019 6239
rect 4813 6205 4847 6239
rect 7849 6205 7883 6239
rect 8125 6205 8159 6239
rect 10977 6205 11011 6239
rect 12633 6205 12667 6239
rect 13737 6205 13771 6239
rect 14004 6205 14038 6239
rect 16865 6205 16899 6239
rect 18153 6205 18187 6239
rect 19257 6205 19291 6239
rect 23489 6205 23523 6239
rect 23949 6205 23983 6239
rect 24133 6205 24167 6239
rect 24400 6205 24434 6239
rect 4353 6137 4387 6171
rect 7665 6137 7699 6171
rect 8392 6137 8426 6171
rect 11069 6137 11103 6171
rect 11621 6137 11655 6171
rect 15853 6137 15887 6171
rect 16313 6137 16347 6171
rect 16773 6137 16807 6171
rect 19073 6137 19107 6171
rect 19524 6137 19558 6171
rect 22385 6137 22419 6171
rect 1409 6069 1443 6103
rect 4905 6069 4939 6103
rect 6193 6069 6227 6103
rect 7849 6069 7883 6103
rect 7941 6069 7975 6103
rect 10149 6069 10183 6103
rect 10609 6069 10643 6103
rect 12817 6069 12851 6103
rect 16405 6069 16439 6103
rect 18337 6069 18371 6103
rect 20637 6069 20671 6103
rect 21833 6069 21867 6103
rect 22017 6069 22051 6103
rect 22477 6069 22511 6103
rect 25513 6069 25547 6103
rect 1593 5865 1627 5899
rect 2789 5865 2823 5899
rect 3433 5865 3467 5899
rect 4537 5865 4571 5899
rect 5641 5865 5675 5899
rect 7481 5865 7515 5899
rect 8033 5865 8067 5899
rect 8493 5865 8527 5899
rect 9689 5865 9723 5899
rect 10885 5865 10919 5899
rect 11253 5865 11287 5899
rect 12541 5865 12575 5899
rect 14105 5865 14139 5899
rect 14657 5865 14691 5899
rect 15025 5865 15059 5899
rect 16129 5865 16163 5899
rect 16497 5865 16531 5899
rect 18797 5865 18831 5899
rect 19717 5865 19751 5899
rect 21649 5865 21683 5899
rect 24409 5865 24443 5899
rect 25053 5865 25087 5899
rect 12992 5797 13026 5831
rect 17040 5797 17074 5831
rect 22109 5797 22143 5831
rect 2697 5729 2731 5763
rect 4445 5729 4479 5763
rect 6009 5729 6043 5763
rect 8401 5729 8435 5763
rect 10057 5729 10091 5763
rect 12725 5729 12759 5763
rect 15301 5729 15335 5763
rect 16773 5729 16807 5763
rect 19625 5729 19659 5763
rect 21097 5729 21131 5763
rect 22201 5729 22235 5763
rect 22468 5729 22502 5763
rect 2881 5661 2915 5695
rect 4721 5661 4755 5695
rect 6101 5661 6135 5695
rect 6193 5661 6227 5695
rect 8677 5661 8711 5695
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 11713 5661 11747 5695
rect 19901 5661 19935 5695
rect 25145 5661 25179 5695
rect 25329 5661 25363 5695
rect 4077 5593 4111 5627
rect 7941 5593 7975 5627
rect 19165 5593 19199 5627
rect 24685 5593 24719 5627
rect 2053 5525 2087 5559
rect 2329 5525 2363 5559
rect 3801 5525 3835 5559
rect 5089 5525 5123 5559
rect 5549 5525 5583 5559
rect 6929 5525 6963 5559
rect 9413 5525 9447 5559
rect 11529 5525 11563 5559
rect 15485 5525 15519 5559
rect 18153 5525 18187 5559
rect 19257 5525 19291 5559
rect 20637 5525 20671 5559
rect 21281 5525 21315 5559
rect 23581 5525 23615 5559
rect 1409 5321 1443 5355
rect 2789 5321 2823 5355
rect 3801 5321 3835 5355
rect 4169 5321 4203 5355
rect 9137 5321 9171 5355
rect 11345 5321 11379 5355
rect 11805 5321 11839 5355
rect 13001 5321 13035 5355
rect 13553 5321 13587 5355
rect 14933 5321 14967 5355
rect 17049 5321 17083 5355
rect 17785 5321 17819 5355
rect 20085 5321 20119 5355
rect 21649 5321 21683 5355
rect 24317 5321 24351 5355
rect 25697 5321 25731 5355
rect 8769 5253 8803 5287
rect 10701 5253 10735 5287
rect 12173 5253 12207 5287
rect 16497 5253 16531 5287
rect 19441 5253 19475 5287
rect 24041 5253 24075 5287
rect 24133 5253 24167 5287
rect 25329 5253 25363 5287
rect 2053 5185 2087 5219
rect 3249 5185 3283 5219
rect 6193 5185 6227 5219
rect 13461 5185 13495 5219
rect 14197 5185 14231 5219
rect 15117 5185 15151 5219
rect 18061 5185 18095 5219
rect 21097 5185 21131 5219
rect 23489 5185 23523 5219
rect 24869 5185 24903 5219
rect 1777 5117 1811 5151
rect 4261 5117 4295 5151
rect 6561 5117 6595 5151
rect 6837 5117 6871 5151
rect 7093 5117 7127 5151
rect 9321 5117 9355 5151
rect 12449 5117 12483 5151
rect 13921 5117 13955 5151
rect 14013 5117 14047 5151
rect 18317 5117 18351 5151
rect 20913 5117 20947 5151
rect 22477 5117 22511 5151
rect 24041 5117 24075 5151
rect 24685 5117 24719 5151
rect 4528 5049 4562 5083
rect 9566 5049 9600 5083
rect 14657 5049 14691 5083
rect 15362 5049 15396 5083
rect 17509 5049 17543 5083
rect 21005 5049 21039 5083
rect 23121 5049 23155 5083
rect 1869 4981 1903 5015
rect 2421 4981 2455 5015
rect 5641 4981 5675 5015
rect 8217 4981 8251 5015
rect 12633 4981 12667 5015
rect 20361 4981 20395 5015
rect 20545 4981 20579 5015
rect 22293 4981 22327 5015
rect 22661 4981 22695 5015
rect 24777 4981 24811 5015
rect 1593 4777 1627 4811
rect 1961 4777 1995 4811
rect 2421 4777 2455 4811
rect 3709 4777 3743 4811
rect 4813 4777 4847 4811
rect 5181 4777 5215 4811
rect 5273 4777 5307 4811
rect 6377 4777 6411 4811
rect 6837 4777 6871 4811
rect 8401 4777 8435 4811
rect 9045 4777 9079 4811
rect 9965 4777 9999 4811
rect 12541 4777 12575 4811
rect 13553 4777 13587 4811
rect 15301 4777 15335 4811
rect 16865 4777 16899 4811
rect 17233 4777 17267 4811
rect 19073 4777 19107 4811
rect 19257 4777 19291 4811
rect 19625 4777 19659 4811
rect 19717 4777 19751 4811
rect 21465 4777 21499 4811
rect 22017 4777 22051 4811
rect 22477 4777 22511 4811
rect 24777 4777 24811 4811
rect 11428 4709 11462 4743
rect 17325 4709 17359 4743
rect 21373 4709 21407 4743
rect 2329 4641 2363 4675
rect 6745 4641 6779 4675
rect 8309 4641 8343 4675
rect 10057 4641 10091 4675
rect 11161 4641 11195 4675
rect 14013 4641 14047 4675
rect 15669 4641 15703 4675
rect 16773 4641 16807 4675
rect 20545 4641 20579 4675
rect 22836 4641 22870 4675
rect 25053 4641 25087 4675
rect 2605 4573 2639 4607
rect 3341 4573 3375 4607
rect 5457 4573 5491 4607
rect 6929 4573 6963 4607
rect 8493 4573 8527 4607
rect 14105 4573 14139 4607
rect 14197 4573 14231 4607
rect 15761 4573 15795 4607
rect 15945 4573 15979 4607
rect 16313 4573 16347 4607
rect 17509 4573 17543 4607
rect 19809 4573 19843 4607
rect 21649 4573 21683 4607
rect 22569 4573 22603 4607
rect 4721 4505 4755 4539
rect 7665 4505 7699 4539
rect 9321 4505 9355 4539
rect 10241 4505 10275 4539
rect 13645 4505 13679 4539
rect 15025 4505 15059 4539
rect 18337 4505 18371 4539
rect 21005 4505 21039 4539
rect 2973 4437 3007 4471
rect 4261 4437 4295 4471
rect 5825 4437 5859 4471
rect 6285 4437 6319 4471
rect 7941 4437 7975 4471
rect 10701 4437 10735 4471
rect 11069 4437 11103 4471
rect 13185 4437 13219 4471
rect 14749 4437 14783 4471
rect 17969 4437 18003 4471
rect 18705 4437 18739 4471
rect 23949 4437 23983 4471
rect 25237 4437 25271 4471
rect 5181 4233 5215 4267
rect 6469 4233 6503 4267
rect 11161 4233 11195 4267
rect 11621 4233 11655 4267
rect 12817 4233 12851 4267
rect 14105 4233 14139 4267
rect 15669 4233 15703 4267
rect 15945 4233 15979 4267
rect 16221 4233 16255 4267
rect 17325 4233 17359 4267
rect 18245 4233 18279 4267
rect 19349 4233 19383 4267
rect 21741 4233 21775 4267
rect 23397 4233 23431 4267
rect 25881 4233 25915 4267
rect 4537 4165 4571 4199
rect 4905 4165 4939 4199
rect 5733 4097 5767 4131
rect 7481 4097 7515 4131
rect 7665 4097 7699 4131
rect 10701 4097 10735 4131
rect 12173 4097 12207 4131
rect 2053 4029 2087 4063
rect 2320 4029 2354 4063
rect 5549 4029 5583 4063
rect 5641 4029 5675 4063
rect 10517 4029 10551 4063
rect 7205 3961 7239 3995
rect 7932 3961 7966 3995
rect 9689 3961 9723 3995
rect 13645 4097 13679 4131
rect 15209 4097 15243 4131
rect 12909 4029 12943 4063
rect 14565 4029 14599 4063
rect 15117 4029 15151 4063
rect 17785 4165 17819 4199
rect 16773 4097 16807 4131
rect 18797 4097 18831 4131
rect 19901 4097 19935 4131
rect 21281 4097 21315 4131
rect 24685 4097 24719 4131
rect 25145 4097 25179 4131
rect 16129 4029 16163 4063
rect 16589 4029 16623 4063
rect 18613 4029 18647 4063
rect 20453 4029 20487 4063
rect 21097 4029 21131 4063
rect 22477 4029 22511 4063
rect 24501 4029 24535 4063
rect 13461 3961 13495 3995
rect 15945 3961 15979 3995
rect 16681 3961 16715 3995
rect 20269 3961 20303 3995
rect 22201 3961 22235 3995
rect 24593 3961 24627 3995
rect 25513 3961 25547 3995
rect 1869 3893 1903 3927
rect 3433 3893 3467 3927
rect 4077 3893 4111 3927
rect 9045 3893 9079 3927
rect 9965 3893 9999 3927
rect 10149 3893 10183 3927
rect 10609 3893 10643 3927
rect 12817 3893 12851 3927
rect 13093 3893 13127 3927
rect 13553 3893 13587 3927
rect 14657 3893 14691 3927
rect 15025 3893 15059 3927
rect 18705 3893 18739 3927
rect 20453 3893 20487 3927
rect 20545 3893 20579 3927
rect 20729 3893 20763 3927
rect 21189 3893 21223 3927
rect 22661 3893 22695 3927
rect 23121 3893 23155 3927
rect 23949 3893 23983 3927
rect 24133 3893 24167 3927
rect 2053 3689 2087 3723
rect 2513 3689 2547 3723
rect 3065 3689 3099 3723
rect 3433 3689 3467 3723
rect 6561 3689 6595 3723
rect 8401 3689 8435 3723
rect 8585 3689 8619 3723
rect 10333 3689 10367 3723
rect 10793 3689 10827 3723
rect 12265 3689 12299 3723
rect 13093 3689 13127 3723
rect 13369 3689 13403 3723
rect 13737 3689 13771 3723
rect 15025 3689 15059 3723
rect 15301 3689 15335 3723
rect 15669 3689 15703 3723
rect 16405 3689 16439 3723
rect 16773 3689 16807 3723
rect 17417 3689 17451 3723
rect 18521 3689 18555 3723
rect 19073 3689 19107 3723
rect 20269 3689 20303 3723
rect 20913 3689 20947 3723
rect 21281 3689 21315 3723
rect 21925 3689 21959 3723
rect 22293 3689 22327 3723
rect 23029 3689 23063 3723
rect 4322 3621 4356 3655
rect 7021 3621 7055 3655
rect 9045 3621 9079 3655
rect 15761 3621 15795 3655
rect 18429 3621 18463 3655
rect 19533 3621 19567 3655
rect 20729 3621 20763 3655
rect 23848 3621 23882 3655
rect 2421 3553 2455 3587
rect 6193 3553 6227 3587
rect 6929 3553 6963 3587
rect 7941 3553 7975 3587
rect 9781 3553 9815 3587
rect 10885 3553 10919 3587
rect 11152 3553 11186 3587
rect 16865 3553 16899 3587
rect 19717 3553 19751 3587
rect 22477 3553 22511 3587
rect 2697 3485 2731 3519
rect 4077 3485 4111 3519
rect 5457 3417 5491 3451
rect 7205 3485 7239 3519
rect 13829 3485 13863 3519
rect 13921 3485 13955 3519
rect 15853 3485 15887 3519
rect 18613 3485 18647 3519
rect 21373 3485 21407 3519
rect 21465 3485 21499 3519
rect 23581 3485 23615 3519
rect 6469 3417 6503 3451
rect 9413 3417 9447 3451
rect 17969 3417 18003 3451
rect 22661 3417 22695 3451
rect 1685 3349 1719 3383
rect 3893 3349 3927 3383
rect 6101 3349 6135 3383
rect 6193 3349 6227 3383
rect 7573 3349 7607 3383
rect 9965 3349 9999 3383
rect 14657 3349 14691 3383
rect 17049 3349 17083 3383
rect 18061 3349 18095 3383
rect 19901 3349 19935 3383
rect 23489 3349 23523 3383
rect 24961 3349 24995 3383
rect 2973 3145 3007 3179
rect 6837 3145 6871 3179
rect 7849 3145 7883 3179
rect 8677 3145 8711 3179
rect 10977 3145 11011 3179
rect 12449 3145 12483 3179
rect 13553 3145 13587 3179
rect 14473 3145 14507 3179
rect 14565 3145 14599 3179
rect 16129 3145 16163 3179
rect 17049 3145 17083 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 19441 3145 19475 3179
rect 20177 3145 20211 3179
rect 23121 3145 23155 3179
rect 25513 3145 25547 3179
rect 11897 3077 11931 3111
rect 6285 3009 6319 3043
rect 7297 3009 7331 3043
rect 7389 3009 7423 3043
rect 8861 3009 8895 3043
rect 11345 3009 11379 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 14289 3009 14323 3043
rect 26065 3077 26099 3111
rect 18061 3009 18095 3043
rect 1593 2941 1627 2975
rect 3709 2941 3743 2975
rect 4077 2941 4111 2975
rect 4261 2941 4295 2975
rect 4517 2941 4551 2975
rect 7205 2941 7239 2975
rect 9117 2941 9151 2975
rect 12173 2941 12207 2975
rect 12817 2941 12851 2975
rect 14473 2941 14507 2975
rect 14749 2941 14783 2975
rect 15005 2941 15039 2975
rect 16681 2941 16715 2975
rect 18317 2941 18351 2975
rect 20545 2941 20579 2975
rect 20637 2941 20671 2975
rect 20904 2941 20938 2975
rect 23397 2941 23431 2975
rect 23949 2941 23983 2975
rect 24133 2941 24167 2975
rect 24400 2941 24434 2975
rect 1860 2873 1894 2907
rect 8309 2873 8343 2907
rect 5641 2805 5675 2839
rect 6561 2805 6595 2839
rect 10241 2805 10275 2839
rect 13829 2805 13863 2839
rect 22017 2805 22051 2839
rect 22569 2805 22603 2839
rect 1593 2601 1627 2635
rect 1869 2601 1903 2635
rect 2329 2601 2363 2635
rect 2881 2601 2915 2635
rect 3893 2601 3927 2635
rect 5733 2601 5767 2635
rect 6929 2601 6963 2635
rect 8493 2601 8527 2635
rect 9781 2601 9815 2635
rect 14013 2601 14047 2635
rect 15209 2601 15243 2635
rect 16865 2601 16899 2635
rect 18061 2601 18095 2635
rect 19717 2601 19751 2635
rect 21005 2601 21039 2635
rect 22569 2601 22603 2635
rect 24225 2601 24259 2635
rect 2237 2533 2271 2567
rect 10977 2533 11011 2567
rect 12081 2533 12115 2567
rect 12878 2533 12912 2567
rect 18604 2533 18638 2567
rect 20637 2533 20671 2567
rect 21456 2533 21490 2567
rect 4353 2465 4387 2499
rect 4620 2465 4654 2499
rect 6377 2465 6411 2499
rect 7297 2465 7331 2499
rect 8585 2465 8619 2499
rect 9597 2465 9631 2499
rect 10149 2465 10183 2499
rect 11253 2465 11287 2499
rect 11437 2465 11471 2499
rect 15485 2465 15519 2499
rect 15741 2465 15775 2499
rect 17693 2465 17727 2499
rect 18337 2465 18371 2499
rect 21189 2465 21223 2499
rect 24593 2465 24627 2499
rect 2513 2397 2547 2431
rect 3525 2397 3559 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 7941 2397 7975 2431
rect 10241 2397 10275 2431
rect 10425 2397 10459 2431
rect 12357 2397 12391 2431
rect 12633 2397 12667 2431
rect 14933 2397 14967 2431
rect 23489 2397 23523 2431
rect 24685 2397 24719 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 9137 2329 9171 2363
rect 8769 2261 8803 2295
rect 11621 2261 11655 2295
rect 23765 2261 23799 2295
<< metal1 >>
rect 14090 26256 14096 26308
rect 14148 26296 14154 26308
rect 24762 26296 24768 26308
rect 14148 26268 24768 26296
rect 14148 26256 14154 26268
rect 24762 26256 24768 26268
rect 24820 26256 24826 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 23845 22763 23903 22769
rect 23845 22729 23857 22763
rect 23891 22760 23903 22763
rect 24670 22760 24676 22772
rect 23891 22732 24676 22760
rect 23891 22729 23903 22732
rect 23845 22723 23903 22729
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 23658 22556 23664 22568
rect 23619 22528 23664 22556
rect 23658 22516 23664 22528
rect 23716 22556 23722 22568
rect 24121 22559 24179 22565
rect 24121 22556 24133 22559
rect 23716 22528 24133 22556
rect 23716 22516 23722 22528
rect 24121 22525 24133 22528
rect 24167 22525 24179 22559
rect 24121 22519 24179 22525
rect 1394 22380 1400 22432
rect 1452 22420 1458 22432
rect 1673 22423 1731 22429
rect 1673 22420 1685 22423
rect 1452 22392 1685 22420
rect 1452 22380 1458 22392
rect 1673 22389 1685 22392
rect 1719 22420 1731 22423
rect 2682 22420 2688 22432
rect 1719 22392 2688 22420
rect 1719 22389 1731 22392
rect 1673 22383 1731 22389
rect 2682 22380 2688 22392
rect 2740 22380 2746 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 24581 22083 24639 22089
rect 24581 22049 24593 22083
rect 24627 22080 24639 22083
rect 24627 22052 24716 22080
rect 24627 22049 24639 22052
rect 24581 22043 24639 22049
rect 24688 22024 24716 22052
rect 24670 21972 24676 22024
rect 24728 21972 24734 22024
rect 24762 21944 24768 21956
rect 24723 21916 24768 21944
rect 24762 21904 24768 21916
rect 24820 21904 24826 21956
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 24578 21332 24584 21344
rect 24539 21304 24584 21332
rect 24578 21292 24584 21304
rect 24636 21292 24642 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 24762 21128 24768 21140
rect 24723 21100 24768 21128
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 24210 20952 24216 21004
rect 24268 20992 24274 21004
rect 24581 20995 24639 21001
rect 24581 20992 24593 20995
rect 24268 20964 24593 20992
rect 24268 20952 24274 20964
rect 24581 20961 24593 20964
rect 24627 20961 24639 20995
rect 24581 20955 24639 20961
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 2682 20584 2688 20596
rect 2643 20556 2688 20584
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20448 13415 20451
rect 13403 20420 13584 20448
rect 13403 20417 13415 20420
rect 13357 20411 13415 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 2501 20383 2559 20389
rect 1443 20352 2084 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2056 20256 2084 20352
rect 2501 20349 2513 20383
rect 2547 20380 2559 20383
rect 13446 20380 13452 20392
rect 2547 20352 3096 20380
rect 13407 20352 13452 20380
rect 2547 20349 2559 20352
rect 2501 20343 2559 20349
rect 3068 20256 3096 20352
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 13556 20380 13584 20420
rect 13722 20389 13728 20392
rect 13716 20380 13728 20389
rect 13556 20352 13728 20380
rect 13716 20343 13728 20352
rect 13722 20340 13728 20343
rect 13780 20340 13786 20392
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 3050 20204 3056 20256
rect 3108 20244 3114 20256
rect 3108 20216 3153 20244
rect 3108 20204 3114 20216
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 14700 20216 14841 20244
rect 14700 20204 14706 20216
rect 14829 20213 14841 20216
rect 14875 20213 14887 20247
rect 14829 20207 14887 20213
rect 24210 20204 24216 20256
rect 24268 20244 24274 20256
rect 24581 20247 24639 20253
rect 24581 20244 24593 20247
rect 24268 20216 24593 20244
rect 24268 20204 24274 20216
rect 24581 20213 24593 20216
rect 24627 20213 24639 20247
rect 24581 20207 24639 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1486 20000 1492 20052
rect 1544 20040 1550 20052
rect 1581 20043 1639 20049
rect 1581 20040 1593 20043
rect 1544 20012 1593 20040
rect 1544 20000 1550 20012
rect 1581 20009 1593 20012
rect 1627 20009 1639 20043
rect 1581 20003 1639 20009
rect 2038 20000 2044 20052
rect 2096 20040 2102 20052
rect 2685 20043 2743 20049
rect 2685 20040 2697 20043
rect 2096 20012 2697 20040
rect 2096 20000 2102 20012
rect 2685 20009 2697 20012
rect 2731 20009 2743 20043
rect 2685 20003 2743 20009
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2406 19904 2412 19916
rect 1443 19876 2412 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19904 2559 19907
rect 2590 19904 2596 19916
rect 2547 19876 2596 19904
rect 2547 19873 2559 19876
rect 2501 19867 2559 19873
rect 2590 19864 2596 19876
rect 2648 19864 2654 19916
rect 13446 19700 13452 19712
rect 13407 19672 13452 19700
rect 13446 19660 13452 19672
rect 13504 19660 13510 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1854 19320 1860 19372
rect 1912 19360 1918 19372
rect 3326 19360 3332 19372
rect 1912 19332 3332 19360
rect 1912 19320 1918 19332
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1670 19292 1676 19304
rect 1443 19264 1676 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 13464 19168 13492 19255
rect 13716 19227 13774 19233
rect 13716 19193 13728 19227
rect 13762 19224 13774 19227
rect 13814 19224 13820 19236
rect 13762 19196 13820 19224
rect 13762 19193 13774 19196
rect 13716 19187 13774 19193
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 1394 19116 1400 19168
rect 1452 19156 1458 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 1452 19128 1593 19156
rect 1452 19116 1458 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 1581 19119 1639 19125
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2406 19156 2412 19168
rect 2087 19128 2412 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 2590 19156 2596 19168
rect 2551 19128 2596 19156
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 13357 19159 13415 19165
rect 13357 19125 13369 19159
rect 13403 19156 13415 19159
rect 13446 19156 13452 19168
rect 13403 19128 13452 19156
rect 13403 19125 13415 19128
rect 13357 19119 13415 19125
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 14826 19156 14832 19168
rect 14787 19128 14832 19156
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 12342 18952 12348 18964
rect 12303 18924 12348 18952
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18816 12311 18819
rect 12713 18819 12771 18825
rect 12713 18816 12725 18819
rect 12299 18788 12725 18816
rect 12299 18785 12311 18788
rect 12253 18779 12311 18785
rect 12713 18785 12725 18788
rect 12759 18816 12771 18819
rect 12894 18816 12900 18828
rect 12759 18788 12900 18816
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 14826 18816 14832 18828
rect 13004 18788 14832 18816
rect 1670 18748 1676 18760
rect 1631 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 13004 18757 13032 18788
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12492 18720 12817 18748
rect 12492 18708 12498 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 12989 18751 13047 18757
rect 12989 18717 13001 18751
rect 13035 18717 13047 18751
rect 13906 18748 13912 18760
rect 13867 18720 13912 18748
rect 12989 18711 13047 18717
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 13004 18680 13032 18711
rect 13906 18708 13912 18720
rect 13964 18708 13970 18760
rect 12308 18652 13032 18680
rect 12308 18640 12314 18652
rect 10413 18615 10471 18621
rect 10413 18581 10425 18615
rect 10459 18612 10471 18615
rect 10962 18612 10968 18624
rect 10459 18584 10968 18612
rect 10459 18581 10471 18584
rect 10413 18575 10471 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 13541 18615 13599 18621
rect 13541 18581 13553 18615
rect 13587 18612 13599 18615
rect 13814 18612 13820 18624
rect 13587 18584 13820 18612
rect 13587 18581 13599 18584
rect 13541 18575 13599 18581
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 11517 18411 11575 18417
rect 11517 18377 11529 18411
rect 11563 18408 11575 18411
rect 12434 18408 12440 18420
rect 11563 18380 12440 18408
rect 11563 18377 11575 18380
rect 11517 18371 11575 18377
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 10321 18343 10379 18349
rect 10321 18340 10333 18343
rect 9732 18312 10333 18340
rect 9732 18300 9738 18312
rect 10321 18309 10333 18312
rect 10367 18309 10379 18343
rect 12250 18340 12256 18352
rect 12211 18312 12256 18340
rect 10321 18303 10379 18309
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 10962 18272 10968 18284
rect 10923 18244 10968 18272
rect 10962 18232 10968 18244
rect 11020 18232 11026 18284
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 1443 18176 2084 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2056 18080 2084 18176
rect 11808 18176 12449 18204
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 10781 18139 10839 18145
rect 10781 18136 10793 18139
rect 10100 18108 10793 18136
rect 10100 18096 10106 18108
rect 10781 18105 10793 18108
rect 10827 18105 10839 18139
rect 10781 18099 10839 18105
rect 2038 18068 2044 18080
rect 1999 18040 2044 18068
rect 2038 18028 2044 18040
rect 2096 18028 2102 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10137 18071 10195 18077
rect 10137 18068 10149 18071
rect 9824 18040 10149 18068
rect 9824 18028 9830 18040
rect 10137 18037 10149 18040
rect 10183 18068 10195 18071
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10183 18040 10701 18068
rect 10183 18037 10195 18040
rect 10137 18031 10195 18037
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 10689 18031 10747 18037
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11808 18077 11836 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12710 18145 12716 18148
rect 12704 18136 12716 18145
rect 12671 18108 12716 18136
rect 12704 18099 12716 18108
rect 12710 18096 12716 18099
rect 12768 18096 12774 18148
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11480 18040 11805 18068
rect 11480 18028 11486 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 11793 18031 11851 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 1762 17864 1768 17876
rect 1627 17836 1768 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 1762 17824 1768 17836
rect 1820 17824 1826 17876
rect 9309 17867 9367 17873
rect 9309 17833 9321 17867
rect 9355 17864 9367 17867
rect 9582 17864 9588 17876
rect 9355 17836 9588 17864
rect 9355 17833 9367 17836
rect 9309 17827 9367 17833
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 11330 17824 11336 17876
rect 11388 17864 11394 17876
rect 12437 17867 12495 17873
rect 12437 17864 12449 17867
rect 11388 17836 12449 17864
rect 11388 17824 11394 17836
rect 12437 17833 12449 17836
rect 12483 17833 12495 17867
rect 12437 17827 12495 17833
rect 12452 17796 12480 17827
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 13541 17867 13599 17873
rect 13541 17864 13553 17867
rect 12952 17836 13553 17864
rect 12952 17824 12958 17836
rect 13541 17833 13553 17836
rect 13587 17833 13599 17867
rect 14642 17864 14648 17876
rect 14603 17836 14648 17864
rect 13541 17827 13599 17833
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 12710 17796 12716 17808
rect 12452 17768 12716 17796
rect 12710 17756 12716 17768
rect 12768 17796 12774 17808
rect 12989 17799 13047 17805
rect 12989 17796 13001 17799
rect 12768 17768 13001 17796
rect 12768 17756 12774 17768
rect 12989 17765 13001 17768
rect 13035 17765 13047 17799
rect 12989 17759 13047 17765
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 2314 17728 2320 17740
rect 1443 17700 2320 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 10318 17688 10324 17740
rect 10376 17728 10382 17740
rect 11313 17731 11371 17737
rect 11313 17728 11325 17731
rect 10376 17700 11325 17728
rect 10376 17688 10382 17700
rect 11313 17697 11325 17700
rect 11359 17728 11371 17731
rect 11882 17728 11888 17740
rect 11359 17700 11888 17728
rect 11359 17697 11371 17700
rect 11313 17691 11371 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 13538 17688 13544 17740
rect 13596 17728 13602 17740
rect 13906 17728 13912 17740
rect 13596 17700 13912 17728
rect 13596 17688 13602 17700
rect 13906 17688 13912 17700
rect 13964 17688 13970 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 11057 17663 11115 17669
rect 11057 17629 11069 17663
rect 11103 17629 11115 17663
rect 13998 17660 14004 17672
rect 13959 17632 14004 17660
rect 11057 17623 11115 17629
rect 10042 17484 10048 17536
rect 10100 17524 10106 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 10100 17496 10333 17524
rect 10100 17484 10106 17496
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10870 17524 10876 17536
rect 10831 17496 10876 17524
rect 10321 17487 10379 17493
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11072 17524 11100 17623
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 13814 17592 13820 17604
rect 13372 17564 13820 17592
rect 13372 17536 13400 17564
rect 13814 17552 13820 17564
rect 13872 17592 13878 17604
rect 14108 17592 14136 17623
rect 13872 17564 14136 17592
rect 13872 17552 13878 17564
rect 24578 17552 24584 17604
rect 24636 17592 24642 17604
rect 24762 17592 24768 17604
rect 24636 17564 24768 17592
rect 24636 17552 24642 17564
rect 24762 17552 24768 17564
rect 24820 17552 24826 17604
rect 11422 17524 11428 17536
rect 11072 17496 11428 17524
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 13354 17524 13360 17536
rect 13315 17496 13360 17524
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1486 17280 1492 17332
rect 1544 17320 1550 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1544 17292 1593 17320
rect 1544 17280 1550 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 2314 17320 2320 17332
rect 2275 17292 2320 17320
rect 1581 17283 1639 17289
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 10318 17320 10324 17332
rect 10279 17292 10324 17320
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 24762 17320 24768 17332
rect 12492 17292 12537 17320
rect 24723 17292 24768 17320
rect 12492 17280 12498 17292
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 11885 17255 11943 17261
rect 11885 17252 11897 17255
rect 11480 17224 11897 17252
rect 11480 17212 11486 17224
rect 11885 17221 11897 17224
rect 11931 17252 11943 17255
rect 13446 17252 13452 17264
rect 11931 17224 13452 17252
rect 11931 17221 11943 17224
rect 11885 17215 11943 17221
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 8352 17156 9137 17184
rect 8352 17144 8358 17156
rect 9125 17153 9137 17156
rect 9171 17184 9183 17187
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9171 17156 9781 17184
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 11330 17184 11336 17196
rect 11291 17156 11336 17184
rect 9769 17147 9827 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12584 17156 13001 17184
rect 12584 17144 12590 17156
rect 12989 17153 13001 17156
rect 13035 17184 13047 17187
rect 13354 17184 13360 17196
rect 13035 17156 13360 17184
rect 13035 17153 13047 17156
rect 12989 17147 13047 17153
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 14642 17184 14648 17196
rect 14603 17156 14648 17184
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 9582 17116 9588 17128
rect 1443 17088 2084 17116
rect 9543 17088 9588 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2056 16992 2084 17088
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 10928 17088 11161 17116
rect 10928 17076 10934 17088
rect 11149 17085 11161 17088
rect 11195 17116 11207 17119
rect 13078 17116 13084 17128
rect 11195 17088 13084 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 13998 17116 14004 17128
rect 13587 17088 14004 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 13998 17076 14004 17088
rect 14056 17116 14062 17128
rect 14056 17088 14596 17116
rect 14056 17076 14062 17088
rect 10594 17048 10600 17060
rect 10555 17020 10600 17048
rect 10594 17008 10600 17020
rect 10652 17048 10658 17060
rect 11238 17048 11244 17060
rect 10652 17020 11244 17048
rect 10652 17008 10658 17020
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 12805 17051 12863 17057
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 13909 17051 13967 17057
rect 13909 17048 13921 17051
rect 12851 17020 13921 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 13909 17017 13921 17020
rect 13955 17048 13967 17051
rect 14461 17051 14519 17057
rect 14461 17048 14473 17051
rect 13955 17020 14473 17048
rect 13955 17017 13967 17020
rect 13909 17011 13967 17017
rect 14461 17017 14473 17020
rect 14507 17017 14519 17051
rect 14461 17011 14519 17017
rect 2038 16980 2044 16992
rect 1999 16952 2044 16980
rect 2038 16940 2044 16952
rect 2096 16940 2102 16992
rect 9214 16980 9220 16992
rect 9175 16952 9220 16980
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 9306 16940 9312 16992
rect 9364 16980 9370 16992
rect 9677 16983 9735 16989
rect 9677 16980 9689 16983
rect 9364 16952 9689 16980
rect 9364 16940 9370 16952
rect 9677 16949 9689 16952
rect 9723 16949 9735 16983
rect 9677 16943 9735 16949
rect 10781 16983 10839 16989
rect 10781 16949 10793 16983
rect 10827 16980 10839 16983
rect 10870 16980 10876 16992
rect 10827 16952 10876 16980
rect 10827 16949 10839 16952
rect 10781 16943 10839 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12161 16983 12219 16989
rect 12161 16980 12173 16983
rect 12032 16952 12173 16980
rect 12032 16940 12038 16952
rect 12161 16949 12173 16952
rect 12207 16980 12219 16983
rect 12820 16980 12848 17011
rect 12207 16952 12848 16980
rect 12207 16949 12219 16952
rect 12161 16943 12219 16949
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 12952 16952 12997 16980
rect 12952 16940 12958 16952
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 14001 16983 14059 16989
rect 14001 16980 14013 16983
rect 13872 16952 14013 16980
rect 13872 16940 13878 16952
rect 14001 16949 14013 16952
rect 14047 16949 14059 16983
rect 14001 16943 14059 16949
rect 14369 16983 14427 16989
rect 14369 16949 14381 16983
rect 14415 16980 14427 16983
rect 14568 16980 14596 17088
rect 23382 17076 23388 17128
rect 23440 17116 23446 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 23440 17088 24593 17116
rect 23440 17076 23446 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24627 17088 25145 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 14826 17008 14832 17060
rect 14884 17048 14890 17060
rect 15565 17051 15623 17057
rect 15565 17048 15577 17051
rect 14884 17020 15577 17048
rect 14884 17008 14890 17020
rect 15565 17017 15577 17020
rect 15611 17017 15623 17051
rect 15565 17011 15623 17017
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 14415 16952 15117 16980
rect 14415 16949 14427 16952
rect 14369 16943 14427 16949
rect 15105 16949 15117 16952
rect 15151 16980 15163 16983
rect 15470 16980 15476 16992
rect 15151 16952 15476 16980
rect 15151 16949 15163 16952
rect 15105 16943 15163 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 24394 16980 24400 16992
rect 24355 16952 24400 16980
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 9306 16776 9312 16788
rect 9267 16748 9312 16776
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 11330 16776 11336 16788
rect 10459 16748 11336 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12526 16776 12532 16788
rect 12487 16748 12532 16776
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 13538 16776 13544 16788
rect 13499 16748 13544 16776
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 14148 16748 14193 16776
rect 14148 16736 14154 16748
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14700 16748 15025 16776
rect 14700 16736 14706 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15013 16739 15071 16745
rect 23753 16779 23811 16785
rect 23753 16745 23765 16779
rect 23799 16776 23811 16779
rect 24394 16776 24400 16788
rect 23799 16748 24400 16776
rect 23799 16745 23811 16748
rect 23753 16739 23811 16745
rect 10686 16668 10692 16720
rect 10744 16717 10750 16720
rect 10744 16711 10808 16717
rect 10744 16677 10762 16711
rect 10796 16677 10808 16711
rect 10744 16671 10808 16677
rect 10744 16668 10750 16671
rect 10870 16668 10876 16720
rect 10928 16708 10934 16720
rect 12894 16708 12900 16720
rect 10928 16680 12900 16708
rect 10928 16668 10934 16680
rect 12894 16668 12900 16680
rect 12952 16668 12958 16720
rect 13078 16668 13084 16720
rect 13136 16708 13142 16720
rect 13998 16708 14004 16720
rect 13136 16680 14004 16708
rect 13136 16668 13142 16680
rect 13998 16668 14004 16680
rect 14056 16668 14062 16720
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1486 16640 1492 16652
rect 1443 16612 1492 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1486 16600 1492 16612
rect 1544 16600 1550 16652
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 11330 16640 11336 16652
rect 10551 16612 11336 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 14108 16640 14136 16736
rect 15028 16708 15056 16739
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 24762 16776 24768 16788
rect 24723 16748 24768 16776
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 15534 16711 15592 16717
rect 15534 16708 15546 16711
rect 15028 16680 15546 16708
rect 15534 16677 15546 16680
rect 15580 16677 15592 16711
rect 15534 16671 15592 16677
rect 13832 16612 14136 16640
rect 23569 16643 23627 16649
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13832 16572 13860 16612
rect 23569 16609 23581 16643
rect 23615 16640 23627 16643
rect 23842 16640 23848 16652
rect 23615 16612 23848 16640
rect 23615 16609 23627 16612
rect 23569 16603 23627 16609
rect 23842 16600 23848 16612
rect 23900 16600 23906 16652
rect 24118 16600 24124 16652
rect 24176 16640 24182 16652
rect 24581 16643 24639 16649
rect 24581 16640 24593 16643
rect 24176 16612 24593 16640
rect 24176 16600 24182 16612
rect 24581 16609 24593 16612
rect 24627 16609 24639 16643
rect 24581 16603 24639 16609
rect 13412 16544 13860 16572
rect 14277 16575 14335 16581
rect 13412 16532 13418 16544
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 14642 16572 14648 16584
rect 14323 16544 14648 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 15286 16572 15292 16584
rect 15247 16544 15292 16572
rect 15286 16532 15292 16544
rect 15344 16532 15350 16584
rect 8849 16439 8907 16445
rect 8849 16405 8861 16439
rect 8895 16436 8907 16439
rect 9398 16436 9404 16448
rect 8895 16408 9404 16436
rect 8895 16405 8907 16408
rect 8849 16399 8907 16405
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 13630 16436 13636 16448
rect 13591 16408 13636 16436
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 16669 16439 16727 16445
rect 16669 16436 16681 16439
rect 15528 16408 16681 16436
rect 15528 16396 15534 16408
rect 16669 16405 16681 16408
rect 16715 16405 16727 16439
rect 16669 16399 16727 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2685 16235 2743 16241
rect 2685 16232 2697 16235
rect 2372 16204 2697 16232
rect 2372 16192 2378 16204
rect 2685 16201 2697 16204
rect 2731 16201 2743 16235
rect 2685 16195 2743 16201
rect 8757 16235 8815 16241
rect 8757 16201 8769 16235
rect 8803 16232 8815 16235
rect 9306 16232 9312 16244
rect 8803 16204 9312 16232
rect 8803 16201 8815 16204
rect 8757 16195 8815 16201
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 10134 16232 10140 16244
rect 10095 16204 10140 16232
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 11422 16232 11428 16244
rect 11383 16204 11428 16232
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 13265 16235 13323 16241
rect 13265 16201 13277 16235
rect 13311 16232 13323 16235
rect 13354 16232 13360 16244
rect 13311 16204 13360 16232
rect 13311 16201 13323 16204
rect 13265 16195 13323 16201
rect 13354 16192 13360 16204
rect 13412 16192 13418 16244
rect 13998 16192 14004 16244
rect 14056 16232 14062 16244
rect 14369 16235 14427 16241
rect 14369 16232 14381 16235
rect 14056 16204 14381 16232
rect 14056 16192 14062 16204
rect 14369 16201 14381 16204
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 24118 16192 24124 16244
rect 24176 16232 24182 16244
rect 24673 16235 24731 16241
rect 24673 16232 24685 16235
rect 24176 16204 24685 16232
rect 24176 16192 24182 16204
rect 24673 16201 24685 16204
rect 24719 16201 24731 16235
rect 24673 16195 24731 16201
rect 1581 16167 1639 16173
rect 1581 16133 1593 16167
rect 1627 16133 1639 16167
rect 1581 16127 1639 16133
rect 1596 16096 1624 16127
rect 2958 16096 2964 16108
rect 1596 16068 2964 16096
rect 2958 16056 2964 16068
rect 3016 16056 3022 16108
rect 8297 16099 8355 16105
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 9306 16096 9312 16108
rect 8343 16068 9312 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 10152 16096 10180 16192
rect 23842 16164 23848 16176
rect 23803 16136 23848 16164
rect 23842 16124 23848 16136
rect 23900 16124 23906 16176
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10152 16068 10885 16096
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 13688 16068 13829 16096
rect 13688 16056 13694 16068
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 14001 16099 14059 16105
rect 14001 16065 14013 16099
rect 14047 16096 14059 16099
rect 14047 16068 15056 16096
rect 14047 16065 14059 16068
rect 14001 16059 14059 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 2493 16031 2551 16037
rect 2493 16028 2505 16031
rect 1397 15991 1455 15997
rect 2424 16000 2505 16028
rect 1412 15892 1440 15991
rect 1486 15920 1492 15972
rect 1544 15960 1550 15972
rect 2317 15963 2375 15969
rect 2317 15960 2329 15963
rect 1544 15932 2329 15960
rect 1544 15920 1550 15932
rect 2317 15929 2329 15932
rect 2363 15929 2375 15963
rect 2424 15960 2452 16000
rect 2493 15997 2505 16000
rect 2539 15997 2551 16031
rect 2493 15991 2551 15997
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 16028 9275 16031
rect 9398 16028 9404 16040
rect 9263 16000 9404 16028
rect 9263 15997 9275 16000
rect 9217 15991 9275 15997
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 9861 16031 9919 16037
rect 9861 15997 9873 16031
rect 9907 16028 9919 16031
rect 10778 16028 10784 16040
rect 9907 16000 10784 16028
rect 9907 15997 9919 16000
rect 9861 15991 9919 15997
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 16028 12311 16031
rect 13722 16028 13728 16040
rect 12299 16000 13728 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 15028 16028 15056 16068
rect 15188 16031 15246 16037
rect 15188 16028 15200 16031
rect 15028 16000 15200 16028
rect 14921 15991 14979 15997
rect 15188 15997 15200 16000
rect 15234 16028 15246 16031
rect 15470 16028 15476 16040
rect 15234 16000 15476 16028
rect 15234 15997 15246 16000
rect 15188 15991 15246 15997
rect 2682 15960 2688 15972
rect 2424 15932 2688 15960
rect 2317 15923 2375 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 2774 15920 2780 15972
rect 2832 15960 2838 15972
rect 3053 15963 3111 15969
rect 3053 15960 3065 15963
rect 2832 15932 3065 15960
rect 2832 15920 2838 15932
rect 3053 15929 3065 15932
rect 3099 15960 3111 15963
rect 7558 15960 7564 15972
rect 3099 15932 7564 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 10689 15963 10747 15969
rect 10689 15929 10701 15963
rect 10735 15960 10747 15963
rect 10870 15960 10876 15972
rect 10735 15932 10876 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 10870 15920 10876 15932
rect 10928 15960 10934 15972
rect 11701 15963 11759 15969
rect 11701 15960 11713 15963
rect 10928 15932 11713 15960
rect 10928 15920 10934 15932
rect 11701 15929 11713 15932
rect 11747 15929 11759 15963
rect 11701 15923 11759 15929
rect 12897 15963 12955 15969
rect 12897 15929 12909 15963
rect 12943 15960 12955 15963
rect 14642 15960 14648 15972
rect 12943 15932 14648 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 14642 15920 14648 15932
rect 14700 15920 14706 15972
rect 14936 15960 14964 15991
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 18046 15988 18052 16000
rect 18104 16028 18110 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18104 16000 18521 16028
rect 18104 15988 18110 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 15286 15960 15292 15972
rect 14752 15932 15292 15960
rect 1854 15892 1860 15904
rect 1412 15864 1860 15892
rect 1854 15852 1860 15864
rect 1912 15892 1918 15904
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1912 15864 1961 15892
rect 1912 15852 1918 15864
rect 1949 15861 1961 15864
rect 1995 15861 2007 15895
rect 8570 15892 8576 15904
rect 8531 15864 8576 15892
rect 1949 15855 2007 15861
rect 8570 15852 8576 15864
rect 8628 15892 8634 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8628 15864 9137 15892
rect 8628 15852 8634 15864
rect 9125 15861 9137 15864
rect 9171 15861 9183 15895
rect 9125 15855 9183 15861
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 10321 15895 10379 15901
rect 10321 15892 10333 15895
rect 9732 15864 10333 15892
rect 9732 15852 9738 15864
rect 10321 15861 10333 15864
rect 10367 15861 10379 15895
rect 13354 15892 13360 15904
rect 13315 15864 13360 15892
rect 10321 15855 10379 15861
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 14752 15901 14780 15932
rect 15286 15920 15292 15932
rect 15344 15960 15350 15972
rect 16853 15963 16911 15969
rect 16853 15960 16865 15963
rect 15344 15932 16865 15960
rect 15344 15920 15350 15932
rect 16853 15929 16865 15932
rect 16899 15929 16911 15963
rect 16853 15923 16911 15929
rect 14737 15895 14795 15901
rect 14737 15892 14749 15895
rect 14608 15864 14749 15892
rect 14608 15852 14614 15864
rect 14737 15861 14749 15864
rect 14783 15861 14795 15895
rect 14737 15855 14795 15861
rect 15930 15852 15936 15904
rect 15988 15892 15994 15904
rect 16301 15895 16359 15901
rect 16301 15892 16313 15895
rect 15988 15864 16313 15892
rect 15988 15852 15994 15864
rect 16301 15861 16313 15864
rect 16347 15861 16359 15895
rect 16301 15855 16359 15861
rect 17770 15852 17776 15904
rect 17828 15892 17834 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 17828 15864 18245 15892
rect 17828 15852 17834 15864
rect 18233 15861 18245 15864
rect 18279 15861 18291 15895
rect 18233 15855 18291 15861
rect 22557 15895 22615 15901
rect 22557 15861 22569 15895
rect 22603 15892 22615 15895
rect 23014 15892 23020 15904
rect 22603 15864 23020 15892
rect 22603 15861 22615 15864
rect 22557 15855 22615 15861
rect 23014 15852 23020 15864
rect 23072 15852 23078 15904
rect 24213 15895 24271 15901
rect 24213 15861 24225 15895
rect 24259 15892 24271 15895
rect 24946 15892 24952 15904
rect 24259 15864 24952 15892
rect 24259 15861 24271 15864
rect 24213 15855 24271 15861
rect 24946 15852 24952 15864
rect 25004 15852 25010 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 8386 15648 8392 15700
rect 8444 15688 8450 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 8444 15660 8493 15688
rect 8444 15648 8450 15660
rect 8481 15657 8493 15660
rect 8527 15688 8539 15691
rect 9214 15688 9220 15700
rect 8527 15660 9220 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 10597 15691 10655 15697
rect 10597 15657 10609 15691
rect 10643 15688 10655 15691
rect 10686 15688 10692 15700
rect 10643 15660 10692 15688
rect 10643 15657 10655 15660
rect 10597 15651 10655 15657
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 11422 15648 11428 15700
rect 11480 15648 11486 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 13630 15688 13636 15700
rect 13127 15660 13636 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 13722 15648 13728 15700
rect 13780 15688 13786 15700
rect 14093 15691 14151 15697
rect 14093 15688 14105 15691
rect 13780 15660 14105 15688
rect 13780 15648 13786 15660
rect 14093 15657 14105 15660
rect 14139 15688 14151 15691
rect 15289 15691 15347 15697
rect 15289 15688 15301 15691
rect 14139 15660 15301 15688
rect 14139 15657 14151 15660
rect 14093 15651 14151 15657
rect 15289 15657 15301 15660
rect 15335 15657 15347 15691
rect 15654 15688 15660 15700
rect 15615 15660 15660 15688
rect 15289 15651 15347 15657
rect 15654 15648 15660 15660
rect 15712 15688 15718 15700
rect 16022 15688 16028 15700
rect 15712 15660 16028 15688
rect 15712 15648 15718 15660
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 24670 15648 24676 15700
rect 24728 15688 24734 15700
rect 24765 15691 24823 15697
rect 24765 15688 24777 15691
rect 24728 15660 24777 15688
rect 24728 15648 24734 15660
rect 24765 15657 24777 15660
rect 24811 15657 24823 15691
rect 24765 15651 24823 15657
rect 11440 15620 11468 15648
rect 10796 15592 11468 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1670 15552 1676 15564
rect 1443 15524 1676 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1670 15512 1676 15524
rect 1728 15512 1734 15564
rect 2593 15555 2651 15561
rect 2593 15521 2605 15555
rect 2639 15521 2651 15555
rect 6822 15552 6828 15564
rect 6783 15524 6828 15552
rect 2593 15515 2651 15521
rect 2608 15484 2636 15515
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 2682 15484 2688 15496
rect 2608 15456 2688 15484
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 6917 15487 6975 15493
rect 6917 15484 6929 15487
rect 6788 15456 6929 15484
rect 6788 15444 6794 15456
rect 6917 15453 6929 15456
rect 6963 15453 6975 15487
rect 7098 15484 7104 15496
rect 7059 15456 7104 15484
rect 6917 15447 6975 15453
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 6457 15419 6515 15425
rect 6457 15385 6469 15419
rect 6503 15416 6515 15419
rect 8404 15416 8432 15515
rect 10318 15512 10324 15564
rect 10376 15552 10382 15564
rect 10796 15561 10824 15592
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 14001 15623 14059 15629
rect 14001 15620 14013 15623
rect 13872 15592 14013 15620
rect 13872 15580 13878 15592
rect 14001 15589 14013 15592
rect 14047 15620 14059 15623
rect 14826 15620 14832 15632
rect 14047 15592 14832 15620
rect 14047 15589 14059 15592
rect 14001 15583 14059 15589
rect 14826 15580 14832 15592
rect 14884 15580 14890 15632
rect 15749 15623 15807 15629
rect 15749 15589 15761 15623
rect 15795 15620 15807 15623
rect 15838 15620 15844 15632
rect 15795 15592 15844 15620
rect 15795 15589 15807 15592
rect 15749 15583 15807 15589
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 10781 15555 10839 15561
rect 10781 15552 10793 15555
rect 10376 15524 10793 15552
rect 10376 15512 10382 15524
rect 10781 15521 10793 15524
rect 10827 15521 10839 15555
rect 10781 15515 10839 15521
rect 11048 15555 11106 15561
rect 11048 15521 11060 15555
rect 11094 15552 11106 15555
rect 11422 15552 11428 15564
rect 11094 15524 11428 15552
rect 11094 15521 11106 15524
rect 11048 15515 11106 15521
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 13044 15524 13461 15552
rect 13044 15512 13050 15524
rect 13449 15521 13461 15524
rect 13495 15552 13507 15555
rect 14737 15555 14795 15561
rect 14737 15552 14749 15555
rect 13495 15524 14749 15552
rect 13495 15521 13507 15524
rect 13449 15515 13507 15521
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 14292 15493 14320 15524
rect 14737 15521 14749 15524
rect 14783 15552 14795 15555
rect 15470 15552 15476 15564
rect 14783 15524 15476 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 17310 15552 17316 15564
rect 16899 15524 17316 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 18230 15512 18236 15564
rect 18288 15552 18294 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 18288 15524 18429 15552
rect 18288 15512 18294 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 19392 15524 19441 15552
rect 19392 15512 19398 15524
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 23566 15552 23572 15564
rect 23527 15524 23572 15552
rect 19429 15515 19487 15521
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 23992 15524 24593 15552
rect 23992 15512 23998 15524
rect 24581 15521 24593 15524
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 8536 15456 8585 15484
rect 8536 15444 8542 15456
rect 8573 15453 8585 15456
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14642 15444 14648 15496
rect 14700 15484 14706 15496
rect 15013 15487 15071 15493
rect 15013 15484 15025 15487
rect 14700 15456 15025 15484
rect 14700 15444 14706 15456
rect 15013 15453 15025 15456
rect 15059 15484 15071 15487
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15059 15456 15853 15484
rect 15059 15453 15071 15456
rect 15013 15447 15071 15453
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 15841 15447 15899 15453
rect 22278 15444 22284 15496
rect 22336 15484 22342 15496
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22336 15456 22569 15484
rect 22336 15444 22342 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 8662 15416 8668 15428
rect 6503 15388 8668 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 13630 15416 13636 15428
rect 13591 15388 13636 15416
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 2777 15351 2835 15357
rect 2777 15348 2789 15351
rect 2740 15320 2789 15348
rect 2740 15308 2746 15320
rect 2777 15317 2789 15320
rect 2823 15317 2835 15351
rect 4246 15348 4252 15360
rect 4207 15320 4252 15348
rect 2777 15311 2835 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15348 8079 15351
rect 9582 15348 9588 15360
rect 8067 15320 9588 15348
rect 8067 15317 8079 15320
rect 8021 15311 8079 15317
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 11756 15320 12173 15348
rect 11756 15308 11762 15320
rect 12161 15317 12173 15320
rect 12207 15317 12219 15351
rect 12161 15311 12219 15317
rect 16393 15351 16451 15357
rect 16393 15317 16405 15351
rect 16439 15348 16451 15351
rect 16482 15348 16488 15360
rect 16439 15320 16488 15348
rect 16439 15317 16451 15320
rect 16393 15311 16451 15317
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 16758 15348 16764 15360
rect 16719 15320 16764 15348
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 17034 15348 17040 15360
rect 16995 15320 17040 15348
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 18322 15308 18328 15360
rect 18380 15348 18386 15360
rect 18601 15351 18659 15357
rect 18601 15348 18613 15351
rect 18380 15320 18613 15348
rect 18380 15308 18386 15320
rect 18601 15317 18613 15320
rect 18647 15317 18659 15351
rect 18601 15311 18659 15317
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 19484 15320 19625 15348
rect 19484 15308 19490 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 23750 15348 23756 15360
rect 23711 15320 23756 15348
rect 19613 15311 19671 15317
rect 23750 15308 23756 15320
rect 23808 15308 23814 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2682 15144 2688 15156
rect 2547 15116 2688 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 2516 14940 2544 15107
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 2832 15116 3893 15144
rect 2832 15104 2838 15116
rect 3881 15113 3893 15116
rect 3927 15113 3939 15147
rect 7098 15144 7104 15156
rect 7011 15116 7104 15144
rect 3881 15107 3939 15113
rect 7098 15104 7104 15116
rect 7156 15144 7162 15156
rect 8202 15144 8208 15156
rect 7156 15116 8208 15144
rect 7156 15104 7162 15116
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 10318 15144 10324 15156
rect 9824 15116 10324 15144
rect 9824 15104 9830 15116
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 10870 15144 10876 15156
rect 10827 15116 10876 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 12986 15144 12992 15156
rect 12947 15116 12992 15144
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 13814 15144 13820 15156
rect 13403 15116 13820 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 15841 15147 15899 15153
rect 15841 15113 15853 15147
rect 15887 15144 15899 15147
rect 16022 15144 16028 15156
rect 15887 15116 16028 15144
rect 15887 15113 15899 15116
rect 15841 15107 15899 15113
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 24762 15144 24768 15156
rect 24723 15116 24768 15144
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 10686 15036 10692 15088
rect 10744 15076 10750 15088
rect 22281 15079 22339 15085
rect 10744 15048 11376 15076
rect 10744 15036 10750 15048
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 3835 14980 4445 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 4433 14977 4445 14980
rect 4479 15008 4491 15011
rect 5718 15008 5724 15020
rect 4479 14980 5724 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 5718 14968 5724 14980
rect 5776 14968 5782 15020
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 6822 15008 6828 15020
rect 6595 14980 6828 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 6822 14968 6828 14980
rect 6880 15008 6886 15020
rect 11348 15017 11376 15048
rect 22281 15045 22293 15079
rect 22327 15076 22339 15079
rect 22922 15076 22928 15088
rect 22327 15048 22928 15076
rect 22327 15045 22339 15048
rect 22281 15039 22339 15045
rect 22922 15036 22928 15048
rect 22980 15036 22986 15088
rect 11333 15011 11391 15017
rect 6880 14980 8064 15008
rect 6880 14968 6886 14980
rect 4246 14940 4252 14952
rect 1903 14912 2544 14940
rect 4207 14912 4252 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 8036 14940 8064 14980
rect 11333 14977 11345 15011
rect 11379 15008 11391 15011
rect 11606 15008 11612 15020
rect 11379 14980 11612 15008
rect 11379 14977 11391 14980
rect 11333 14971 11391 14977
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16724 14980 16865 15008
rect 16724 14968 16730 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 16853 14971 16911 14977
rect 19168 14980 19993 15008
rect 9490 14940 9496 14952
rect 8036 14912 9496 14940
rect 7929 14903 7987 14909
rect 4341 14875 4399 14881
rect 4341 14872 4353 14875
rect 3344 14844 4353 14872
rect 1670 14804 1676 14816
rect 1631 14776 1676 14804
rect 1670 14764 1676 14776
rect 1728 14764 1734 14816
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 3344 14813 3372 14844
rect 4341 14841 4353 14844
rect 4387 14841 4399 14875
rect 4341 14835 4399 14841
rect 6181 14875 6239 14881
rect 6181 14841 6193 14875
rect 6227 14872 6239 14875
rect 6730 14872 6736 14884
rect 6227 14844 6736 14872
rect 6227 14841 6239 14844
rect 6181 14835 6239 14841
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 7745 14875 7803 14881
rect 7745 14872 7757 14875
rect 7064 14844 7757 14872
rect 7064 14832 7070 14844
rect 7745 14841 7757 14844
rect 7791 14872 7803 14875
rect 7944 14872 7972 14903
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 12342 14900 12348 14952
rect 12400 14940 12406 14952
rect 12986 14940 12992 14952
rect 12400 14912 12992 14940
rect 12400 14900 12406 14912
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 13817 14943 13875 14949
rect 13817 14940 13829 14943
rect 13648 14912 13829 14940
rect 7791 14844 7972 14872
rect 7791 14841 7803 14844
rect 7745 14835 7803 14841
rect 8018 14832 8024 14884
rect 8076 14872 8082 14884
rect 8174 14875 8232 14881
rect 8174 14872 8186 14875
rect 8076 14844 8186 14872
rect 8076 14832 8082 14844
rect 8174 14841 8186 14844
rect 8220 14841 8232 14875
rect 8174 14835 8232 14841
rect 9953 14875 10011 14881
rect 9953 14841 9965 14875
rect 9999 14872 10011 14875
rect 11149 14875 11207 14881
rect 11149 14872 11161 14875
rect 9999 14844 11161 14872
rect 9999 14841 10011 14844
rect 9953 14835 10011 14841
rect 11149 14841 11161 14844
rect 11195 14872 11207 14875
rect 12437 14875 12495 14881
rect 12437 14872 12449 14875
rect 11195 14844 12449 14872
rect 11195 14841 11207 14844
rect 11149 14835 11207 14841
rect 12437 14841 12449 14844
rect 12483 14841 12495 14875
rect 12437 14835 12495 14841
rect 3329 14807 3387 14813
rect 3329 14804 3341 14807
rect 3200 14776 3341 14804
rect 3200 14764 3206 14776
rect 3329 14773 3341 14776
rect 3375 14773 3387 14807
rect 7374 14804 7380 14816
rect 7335 14776 7380 14804
rect 3329 14767 3387 14773
rect 7374 14764 7380 14776
rect 7432 14804 7438 14816
rect 8478 14804 8484 14816
rect 7432 14776 8484 14804
rect 7432 14764 7438 14776
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9309 14807 9367 14813
rect 9309 14773 9321 14807
rect 9355 14804 9367 14807
rect 9858 14804 9864 14816
rect 9355 14776 9864 14804
rect 9355 14773 9367 14776
rect 9309 14767 9367 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 10735 14776 11253 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 11241 14773 11253 14776
rect 11287 14804 11299 14807
rect 11330 14804 11336 14816
rect 11287 14776 11336 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11793 14807 11851 14813
rect 11793 14804 11805 14807
rect 11480 14776 11805 14804
rect 11480 14764 11486 14776
rect 11793 14773 11805 14776
rect 11839 14804 11851 14807
rect 12342 14804 12348 14816
rect 11839 14776 12348 14804
rect 11839 14773 11851 14776
rect 11793 14767 11851 14773
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 13446 14764 13452 14816
rect 13504 14804 13510 14816
rect 13648 14813 13676 14912
rect 13817 14909 13829 14912
rect 13863 14940 13875 14943
rect 14550 14940 14556 14952
rect 13863 14912 14556 14940
rect 13863 14909 13875 14912
rect 13817 14903 13875 14909
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16356 14912 16773 14940
rect 16356 14900 16362 14912
rect 16761 14909 16773 14912
rect 16807 14909 16819 14943
rect 16761 14903 16819 14909
rect 18506 14900 18512 14952
rect 18564 14940 18570 14952
rect 19168 14949 19196 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 19153 14943 19211 14949
rect 19153 14940 19165 14943
rect 18564 14912 19165 14940
rect 18564 14900 18570 14912
rect 19153 14909 19165 14912
rect 19199 14909 19211 14943
rect 19153 14903 19211 14909
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19392 14912 19625 14940
rect 19392 14900 19398 14912
rect 19613 14909 19625 14912
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 22097 14943 22155 14949
rect 22097 14909 22109 14943
rect 22143 14940 22155 14943
rect 24394 14940 24400 14952
rect 22143 14912 22692 14940
rect 24355 14912 24400 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 14084 14875 14142 14881
rect 14084 14872 14096 14875
rect 13964 14844 14096 14872
rect 13964 14832 13970 14844
rect 14084 14841 14096 14844
rect 14130 14872 14142 14875
rect 15930 14872 15936 14884
rect 14130 14844 15936 14872
rect 14130 14841 14142 14844
rect 14084 14835 14142 14841
rect 15930 14832 15936 14844
rect 15988 14832 15994 14884
rect 16209 14875 16267 14881
rect 16209 14841 16221 14875
rect 16255 14872 16267 14875
rect 16669 14875 16727 14881
rect 16669 14872 16681 14875
rect 16255 14844 16681 14872
rect 16255 14841 16267 14844
rect 16209 14835 16267 14841
rect 16669 14841 16681 14844
rect 16715 14872 16727 14875
rect 17218 14872 17224 14884
rect 16715 14844 17224 14872
rect 16715 14841 16727 14844
rect 16669 14835 16727 14841
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 18782 14832 18788 14884
rect 18840 14872 18846 14884
rect 20180 14872 20208 14903
rect 20625 14875 20683 14881
rect 20625 14872 20637 14875
rect 18840 14844 20637 14872
rect 18840 14832 18846 14844
rect 20625 14841 20637 14844
rect 20671 14841 20683 14875
rect 20625 14835 20683 14841
rect 13633 14807 13691 14813
rect 13633 14804 13645 14807
rect 13504 14776 13645 14804
rect 13504 14764 13510 14776
rect 13633 14773 13645 14776
rect 13679 14773 13691 14807
rect 13633 14767 13691 14773
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 15197 14807 15255 14813
rect 15197 14804 15209 14807
rect 13872 14776 15209 14804
rect 13872 14764 13878 14776
rect 15197 14773 15209 14776
rect 15243 14773 15255 14807
rect 15197 14767 15255 14773
rect 16301 14807 16359 14813
rect 16301 14773 16313 14807
rect 16347 14804 16359 14807
rect 16390 14804 16396 14816
rect 16347 14776 16396 14804
rect 16347 14773 16359 14776
rect 16301 14767 16359 14773
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 17310 14804 17316 14816
rect 17271 14776 17316 14804
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 17460 14776 18061 14804
rect 17460 14764 17466 14776
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 18049 14767 18107 14773
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 18509 14807 18567 14813
rect 18509 14804 18521 14807
rect 18288 14776 18521 14804
rect 18288 14764 18294 14776
rect 18509 14773 18521 14776
rect 18555 14773 18567 14807
rect 19334 14804 19340 14816
rect 19295 14776 19340 14804
rect 18509 14767 18567 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 20162 14764 20168 14816
rect 20220 14804 20226 14816
rect 22664 14813 22692 14912
rect 24394 14900 24400 14912
rect 24452 14900 24458 14952
rect 24578 14940 24584 14952
rect 24539 14912 24584 14940
rect 24578 14900 24584 14912
rect 24636 14940 24642 14952
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24636 14912 25145 14940
rect 24636 14900 24642 14912
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 20349 14807 20407 14813
rect 20349 14804 20361 14807
rect 20220 14776 20361 14804
rect 20220 14764 20226 14776
rect 20349 14773 20361 14776
rect 20395 14773 20407 14807
rect 20349 14767 20407 14773
rect 22649 14807 22707 14813
rect 22649 14773 22661 14807
rect 22695 14804 22707 14807
rect 23198 14804 23204 14816
rect 22695 14776 23204 14804
rect 22695 14773 22707 14776
rect 22649 14767 22707 14773
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 23566 14764 23572 14816
rect 23624 14804 23630 14816
rect 23845 14807 23903 14813
rect 23845 14804 23857 14807
rect 23624 14776 23857 14804
rect 23624 14764 23630 14776
rect 23845 14773 23857 14776
rect 23891 14773 23903 14807
rect 23845 14767 23903 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 2590 14560 2596 14612
rect 2648 14600 2654 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2648 14572 2697 14600
rect 2648 14560 2654 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 2685 14563 2743 14569
rect 4065 14603 4123 14609
rect 4065 14569 4077 14603
rect 4111 14600 4123 14603
rect 4246 14600 4252 14612
rect 4111 14572 4252 14600
rect 4111 14569 4123 14572
rect 4065 14563 4123 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 8018 14600 8024 14612
rect 7979 14572 8024 14600
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8386 14600 8392 14612
rect 8347 14572 8392 14600
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 8662 14600 8668 14612
rect 8623 14572 8668 14600
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 11606 14600 11612 14612
rect 11567 14572 11612 14600
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 13541 14603 13599 14609
rect 13541 14569 13553 14603
rect 13587 14600 13599 14603
rect 13722 14600 13728 14612
rect 13587 14572 13728 14600
rect 13587 14569 13599 14572
rect 13541 14563 13599 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 13906 14600 13912 14612
rect 13867 14572 13912 14600
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 17310 14600 17316 14612
rect 15335 14572 17316 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 18598 14600 18604 14612
rect 18559 14572 18604 14600
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 22738 14560 22744 14612
rect 22796 14600 22802 14612
rect 23753 14603 23811 14609
rect 23753 14600 23765 14603
rect 22796 14572 23765 14600
rect 22796 14560 22802 14572
rect 23753 14569 23765 14572
rect 23799 14569 23811 14603
rect 23753 14563 23811 14569
rect 24118 14560 24124 14612
rect 24176 14600 24182 14612
rect 24765 14603 24823 14609
rect 24765 14600 24777 14603
rect 24176 14572 24777 14600
rect 24176 14560 24182 14572
rect 24765 14569 24777 14572
rect 24811 14569 24823 14603
rect 24765 14563 24823 14569
rect 3881 14535 3939 14541
rect 3881 14501 3893 14535
rect 3927 14532 3939 14535
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 3927 14504 4537 14532
rect 3927 14501 3939 14504
rect 3881 14495 3939 14501
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2406 14464 2412 14476
rect 1443 14436 2412 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2406 14424 2412 14436
rect 2464 14424 2470 14476
rect 2501 14467 2559 14473
rect 2501 14433 2513 14467
rect 2547 14433 2559 14467
rect 2501 14427 2559 14433
rect 2314 14356 2320 14408
rect 2372 14396 2378 14408
rect 2516 14396 2544 14427
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 2372 14368 3065 14396
rect 2372 14356 2378 14368
rect 3053 14365 3065 14368
rect 3099 14365 3111 14399
rect 3053 14359 3111 14365
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 3896 14328 3924 14495
rect 5718 14492 5724 14544
rect 5776 14532 5782 14544
rect 5874 14535 5932 14541
rect 5874 14532 5886 14535
rect 5776 14504 5886 14532
rect 5776 14492 5782 14504
rect 5874 14501 5886 14504
rect 5920 14501 5932 14535
rect 15654 14532 15660 14544
rect 15615 14504 15660 14532
rect 5874 14495 5932 14501
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 15746 14492 15752 14544
rect 15804 14532 15810 14544
rect 16298 14532 16304 14544
rect 15804 14504 15849 14532
rect 16259 14504 16304 14532
rect 15804 14492 15810 14504
rect 16298 14492 16304 14504
rect 16356 14492 16362 14544
rect 4430 14464 4436 14476
rect 4391 14436 4436 14464
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 9766 14464 9772 14476
rect 9723 14436 9772 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 9950 14473 9956 14476
rect 9944 14464 9956 14473
rect 9911 14436 9956 14464
rect 9944 14427 9956 14436
rect 9950 14424 9956 14427
rect 10008 14424 10014 14476
rect 11974 14424 11980 14476
rect 12032 14464 12038 14476
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 12032 14436 12541 14464
rect 12032 14424 12038 14436
rect 12529 14433 12541 14436
rect 12575 14433 12587 14467
rect 12529 14427 12587 14433
rect 14185 14467 14243 14473
rect 14185 14433 14197 14467
rect 14231 14464 14243 14467
rect 14642 14464 14648 14476
rect 14231 14436 14648 14464
rect 14231 14433 14243 14436
rect 14185 14427 14243 14433
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 16114 14424 16120 14476
rect 16172 14464 16178 14476
rect 17221 14467 17279 14473
rect 17221 14464 17233 14467
rect 16172 14436 17233 14464
rect 16172 14424 16178 14436
rect 17221 14433 17233 14436
rect 17267 14433 17279 14467
rect 17221 14427 17279 14433
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14464 18475 14467
rect 19058 14464 19064 14476
rect 18463 14436 19064 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 19518 14464 19524 14476
rect 19479 14436 19524 14464
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21450 14464 21456 14476
rect 20947 14436 21456 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21450 14424 21456 14436
rect 21508 14424 21514 14476
rect 21542 14424 21548 14476
rect 21600 14464 21606 14476
rect 22554 14464 22560 14476
rect 21600 14436 22560 14464
rect 21600 14424 21606 14436
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 23569 14467 23627 14473
rect 23569 14433 23581 14467
rect 23615 14464 23627 14467
rect 24118 14464 24124 14476
rect 23615 14436 24124 14464
rect 23615 14433 23627 14436
rect 23569 14427 23627 14433
rect 24118 14424 24124 14436
rect 24176 14424 24182 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 4614 14396 4620 14408
rect 4575 14368 4620 14396
rect 4614 14356 4620 14368
rect 4672 14396 4678 14408
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4672 14368 5089 14396
rect 4672 14356 4678 14368
rect 5077 14365 5089 14368
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 2648 14300 3924 14328
rect 2648 14288 2654 14300
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 5644 14328 5672 14359
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 12492 14368 12633 14396
rect 12492 14356 12498 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14396 12863 14399
rect 12986 14396 12992 14408
rect 12851 14368 12992 14396
rect 12851 14365 12863 14368
rect 12805 14359 12863 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 17310 14396 17316 14408
rect 16684 14368 17316 14396
rect 4212 14300 5672 14328
rect 4212 14288 4218 14300
rect 3418 14260 3424 14272
rect 3379 14232 3424 14260
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 5644 14260 5672 14300
rect 15105 14331 15163 14337
rect 15105 14297 15117 14331
rect 15151 14328 15163 14331
rect 15838 14328 15844 14340
rect 15151 14300 15844 14328
rect 15151 14297 15163 14300
rect 15105 14291 15163 14297
rect 15838 14288 15844 14300
rect 15896 14328 15902 14340
rect 16684 14328 16712 14368
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 16850 14328 16856 14340
rect 15896 14300 16712 14328
rect 16811 14300 16856 14328
rect 15896 14288 15902 14300
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 5994 14260 6000 14272
rect 5644 14232 6000 14260
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 7009 14263 7067 14269
rect 7009 14229 7021 14263
rect 7055 14260 7067 14263
rect 7466 14260 7472 14272
rect 7055 14232 7472 14260
rect 7055 14229 7067 14232
rect 7009 14223 7067 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 11057 14263 11115 14269
rect 11057 14229 11069 14263
rect 11103 14260 11115 14263
rect 11422 14260 11428 14272
rect 11103 14232 11428 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 12161 14263 12219 14269
rect 12161 14260 12173 14263
rect 11756 14232 12173 14260
rect 11756 14220 11762 14232
rect 12161 14229 12173 14232
rect 12207 14229 12219 14263
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 12161 14223 12219 14229
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 14734 14260 14740 14272
rect 14695 14232 14740 14260
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 16666 14260 16672 14272
rect 16627 14232 16672 14260
rect 16666 14220 16672 14232
rect 16724 14260 16730 14272
rect 17420 14260 17448 14359
rect 17862 14260 17868 14272
rect 16724 14232 17868 14260
rect 16724 14220 16730 14232
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 18414 14260 18420 14272
rect 18187 14232 18420 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 19705 14263 19763 14269
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 20530 14260 20536 14272
rect 19751 14232 20536 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 21085 14263 21143 14269
rect 21085 14229 21097 14263
rect 21131 14260 21143 14263
rect 21726 14260 21732 14272
rect 21131 14232 21732 14260
rect 21131 14229 21143 14232
rect 21085 14223 21143 14229
rect 21726 14220 21732 14232
rect 21784 14220 21790 14272
rect 22370 14220 22376 14272
rect 22428 14260 22434 14272
rect 22741 14263 22799 14269
rect 22741 14260 22753 14263
rect 22428 14232 22753 14260
rect 22428 14220 22434 14232
rect 22741 14229 22753 14232
rect 22787 14229 22799 14263
rect 22741 14223 22799 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1946 14056 1952 14068
rect 1627 14028 1952 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 3789 14059 3847 14065
rect 3789 14025 3801 14059
rect 3835 14056 3847 14059
rect 4430 14056 4436 14068
rect 3835 14028 4436 14056
rect 3835 14025 3847 14028
rect 3789 14019 3847 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5592 14028 5641 14056
rect 5592 14016 5598 14028
rect 5629 14025 5641 14028
rect 5675 14056 5687 14059
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 5675 14028 6561 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8570 14056 8576 14068
rect 8076 14028 8576 14056
rect 8076 14016 8082 14028
rect 8570 14016 8576 14028
rect 8628 14056 8634 14068
rect 8665 14059 8723 14065
rect 8665 14056 8677 14059
rect 8628 14028 8677 14056
rect 8628 14016 8634 14028
rect 8665 14025 8677 14028
rect 8711 14025 8723 14059
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 8665 14019 8723 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 10778 14056 10784 14068
rect 10643 14028 10784 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11698 14056 11704 14068
rect 11659 14028 11704 14056
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 12986 14056 12992 14068
rect 12947 14028 12992 14056
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 15930 14056 15936 14068
rect 15611 14028 15936 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 17310 14056 17316 14068
rect 17271 14028 17316 14056
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 19058 14016 19064 14028
rect 19116 14056 19122 14068
rect 19797 14059 19855 14065
rect 19797 14056 19809 14059
rect 19116 14028 19809 14056
rect 19116 14016 19122 14028
rect 19797 14025 19809 14028
rect 19843 14025 19855 14059
rect 19797 14019 19855 14025
rect 22554 14016 22560 14068
rect 22612 14056 22618 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 22612 14028 23397 14056
rect 22612 14016 22618 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 2222 13948 2228 14000
rect 2280 13988 2286 14000
rect 2685 13991 2743 13997
rect 2685 13988 2697 13991
rect 2280 13960 2697 13988
rect 2280 13948 2286 13960
rect 2685 13957 2697 13960
rect 2731 13957 2743 13991
rect 4154 13988 4160 14000
rect 4115 13960 4160 13988
rect 2685 13951 2743 13957
rect 4154 13948 4160 13960
rect 4212 13988 4218 14000
rect 4212 13960 4292 13988
rect 4212 13948 4218 13960
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 2516 13892 3157 13920
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 2038 13852 2044 13864
rect 1443 13824 2044 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2516 13861 2544 13892
rect 3145 13889 3157 13892
rect 3191 13920 3203 13923
rect 3234 13920 3240 13932
rect 3191 13892 3240 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 4264 13929 4292 13960
rect 5994 13948 6000 14000
rect 6052 13988 6058 14000
rect 6181 13991 6239 13997
rect 6181 13988 6193 13991
rect 6052 13960 6193 13988
rect 6052 13948 6058 13960
rect 6181 13957 6193 13960
rect 6227 13988 6239 13991
rect 7006 13988 7012 14000
rect 6227 13960 7012 13988
rect 6227 13957 6239 13960
rect 6181 13951 6239 13957
rect 7006 13948 7012 13960
rect 7064 13988 7070 14000
rect 7101 13991 7159 13997
rect 7101 13988 7113 13991
rect 7064 13960 7113 13988
rect 7064 13948 7070 13960
rect 7101 13957 7113 13960
rect 7147 13957 7159 13991
rect 7101 13951 7159 13957
rect 10505 13991 10563 13997
rect 10505 13957 10517 13991
rect 10551 13988 10563 13991
rect 10686 13988 10692 14000
rect 10551 13960 10692 13988
rect 10551 13957 10563 13960
rect 10505 13951 10563 13957
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 7116 13920 7144 13951
rect 10686 13948 10692 13960
rect 10744 13988 10750 14000
rect 16114 13988 16120 14000
rect 10744 13960 11192 13988
rect 16075 13960 16120 13988
rect 10744 13948 10750 13960
rect 11164 13929 11192 13960
rect 16114 13948 16120 13960
rect 16172 13948 16178 14000
rect 16298 13988 16304 14000
rect 16259 13960 16304 13988
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 21085 13991 21143 13997
rect 17920 13960 18644 13988
rect 17920 13948 17926 13960
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7116 13892 7297 13920
rect 4249 13883 4307 13889
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15654 13920 15660 13932
rect 15160 13892 15660 13920
rect 15160 13880 15166 13892
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 16758 13920 16764 13932
rect 16719 13892 16764 13920
rect 16758 13880 16764 13892
rect 16816 13880 16822 13932
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13920 17003 13923
rect 17494 13920 17500 13932
rect 16991 13892 17500 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 18616 13929 18644 13960
rect 21085 13957 21097 13991
rect 21131 13988 21143 13991
rect 22094 13988 22100 14000
rect 21131 13960 22100 13988
rect 21131 13957 21143 13960
rect 21085 13951 21143 13957
rect 22094 13948 22100 13960
rect 22152 13948 22158 14000
rect 24762 13988 24768 14000
rect 24723 13960 24768 13988
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 17788 13892 18521 13920
rect 4522 13861 4528 13864
rect 2507 13855 2565 13861
rect 2507 13821 2519 13855
rect 2553 13821 2565 13855
rect 4505 13855 4528 13861
rect 4505 13852 4517 13855
rect 2507 13815 2565 13821
rect 4356 13824 4517 13852
rect 3786 13744 3792 13796
rect 3844 13784 3850 13796
rect 4356 13784 4384 13824
rect 4505 13821 4517 13824
rect 4580 13852 4586 13864
rect 9950 13852 9956 13864
rect 4580 13824 5488 13852
rect 4505 13815 4528 13821
rect 4522 13812 4528 13815
rect 4580 13812 4586 13824
rect 3844 13756 4384 13784
rect 5460 13784 5488 13824
rect 8220 13824 9956 13852
rect 5626 13784 5632 13796
rect 5460 13756 5632 13784
rect 3844 13744 3850 13756
rect 5626 13744 5632 13756
rect 5684 13744 5690 13796
rect 7466 13744 7472 13796
rect 7524 13793 7530 13796
rect 7524 13787 7588 13793
rect 7524 13753 7542 13787
rect 7576 13753 7588 13787
rect 7524 13747 7588 13753
rect 7524 13744 7530 13747
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 8220 13784 8248 13824
rect 9950 13812 9956 13824
rect 10008 13852 10014 13864
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 10008 13824 10057 13852
rect 10008 13812 10014 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 11698 13852 11704 13864
rect 11011 13824 11704 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 11974 13812 11980 13864
rect 12032 13852 12038 13864
rect 13814 13861 13820 13864
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 12032 13824 12173 13852
rect 12032 13812 12038 13824
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 12161 13815 12219 13821
rect 13464 13824 13553 13852
rect 8168 13756 8248 13784
rect 8168 13744 8174 13756
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 11057 13787 11115 13793
rect 11057 13784 11069 13787
rect 10836 13756 11069 13784
rect 10836 13744 10842 13756
rect 11057 13753 11069 13756
rect 11103 13753 11115 13787
rect 11057 13747 11115 13753
rect 13464 13728 13492 13824
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13808 13852 13820 13861
rect 13775 13824 13820 13852
rect 13541 13815 13599 13821
rect 13808 13815 13820 13824
rect 13814 13812 13820 13815
rect 13872 13812 13878 13864
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 14792 13824 15148 13852
rect 14792 13812 14798 13824
rect 15120 13784 15148 13824
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 17788 13861 17816 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19518 13920 19524 13932
rect 19300 13892 19524 13920
rect 19300 13880 19306 13892
rect 19518 13880 19524 13892
rect 19576 13920 19582 13932
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 19576 13892 20085 13920
rect 19576 13880 19582 13892
rect 20073 13889 20085 13892
rect 20119 13889 20131 13923
rect 20073 13883 20131 13889
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 23900 13892 24624 13920
rect 23900 13880 23906 13892
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17644 13824 17785 13852
rect 17644 13812 17650 13824
rect 17773 13821 17785 13824
rect 17819 13821 17831 13855
rect 19610 13852 19616 13864
rect 19571 13824 19616 13852
rect 17773 13815 17831 13821
rect 19610 13812 19616 13824
rect 19668 13852 19674 13864
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 19668 13824 20453 13852
rect 19668 13812 19674 13824
rect 20441 13821 20453 13824
rect 20487 13821 20499 13855
rect 20898 13852 20904 13864
rect 20859 13824 20904 13852
rect 20441 13815 20499 13821
rect 20898 13812 20904 13824
rect 20956 13852 20962 13864
rect 21729 13855 21787 13861
rect 21729 13852 21741 13855
rect 20956 13824 21741 13852
rect 20956 13812 20962 13824
rect 21729 13821 21741 13824
rect 21775 13821 21787 13855
rect 21729 13815 21787 13821
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13852 22615 13855
rect 23109 13855 23167 13861
rect 23109 13852 23121 13855
rect 22603 13824 23121 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 23109 13821 23121 13824
rect 23155 13852 23167 13855
rect 23290 13852 23296 13864
rect 23155 13824 23296 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 23937 13855 23995 13861
rect 23937 13821 23949 13855
rect 23983 13852 23995 13855
rect 24118 13852 24124 13864
rect 23983 13824 24124 13852
rect 23983 13821 23995 13824
rect 23937 13815 23995 13821
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 24596 13861 24624 13892
rect 24581 13855 24639 13861
rect 24581 13821 24593 13855
rect 24627 13852 24639 13855
rect 25133 13855 25191 13861
rect 25133 13852 25145 13855
rect 24627 13824 25145 13852
rect 24627 13821 24639 13824
rect 24581 13815 24639 13821
rect 25133 13821 25145 13824
rect 25179 13821 25191 13855
rect 25133 13815 25191 13821
rect 16298 13784 16304 13796
rect 15120 13756 16304 13784
rect 16298 13744 16304 13756
rect 16356 13784 16362 13796
rect 16669 13787 16727 13793
rect 16669 13784 16681 13787
rect 16356 13756 16681 13784
rect 16356 13744 16362 13756
rect 16669 13753 16681 13756
rect 16715 13753 16727 13787
rect 16669 13747 16727 13753
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12492 13688 12633 13716
rect 12492 13676 12498 13688
rect 12621 13685 12633 13688
rect 12667 13685 12679 13719
rect 13446 13716 13452 13728
rect 13407 13688 13452 13716
rect 12621 13679 12679 13685
rect 13446 13676 13452 13688
rect 13504 13676 13510 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 14921 13719 14979 13725
rect 14921 13716 14933 13719
rect 14884 13688 14933 13716
rect 14884 13676 14890 13688
rect 14921 13685 14933 13688
rect 14967 13685 14979 13719
rect 18046 13716 18052 13728
rect 18007 13688 18052 13716
rect 14921 13679 14979 13685
rect 18046 13676 18052 13688
rect 18104 13676 18110 13728
rect 18414 13716 18420 13728
rect 18375 13688 18420 13716
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 21450 13716 21456 13728
rect 21411 13688 21456 13716
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 22462 13676 22468 13728
rect 22520 13716 22526 13728
rect 22741 13719 22799 13725
rect 22741 13716 22753 13719
rect 22520 13688 22753 13716
rect 22520 13676 22526 13688
rect 22741 13685 22753 13688
rect 22787 13685 22799 13719
rect 24394 13716 24400 13728
rect 24355 13688 24400 13716
rect 22741 13679 22799 13685
rect 24394 13676 24400 13688
rect 24452 13716 24458 13728
rect 24670 13716 24676 13728
rect 24452 13688 24676 13716
rect 24452 13676 24458 13688
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1581 13515 1639 13521
rect 1581 13481 1593 13515
rect 1627 13512 1639 13515
rect 2498 13512 2504 13524
rect 1627 13484 2504 13512
rect 1627 13481 1639 13484
rect 1581 13475 1639 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 2682 13512 2688 13524
rect 2643 13484 2688 13512
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8570 13512 8576 13524
rect 8531 13484 8576 13512
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 10778 13512 10784 13524
rect 10735 13484 10784 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11514 13512 11520 13524
rect 11287 13484 11520 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 13630 13512 13636 13524
rect 13591 13484 13636 13512
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 15102 13512 15108 13524
rect 15063 13484 15108 13512
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 15746 13512 15752 13524
rect 15611 13484 15752 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17920 13484 18153 13512
rect 17920 13472 17926 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 18230 13472 18236 13524
rect 18288 13512 18294 13524
rect 18506 13512 18512 13524
rect 18288 13484 18512 13512
rect 18288 13472 18294 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 20070 13512 20076 13524
rect 18739 13484 20076 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 23753 13515 23811 13521
rect 23753 13481 23765 13515
rect 23799 13512 23811 13515
rect 24394 13512 24400 13524
rect 23799 13484 24400 13512
rect 23799 13481 23811 13484
rect 23753 13475 23811 13481
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 24762 13512 24768 13524
rect 24723 13484 24768 13512
rect 24762 13472 24768 13484
rect 24820 13472 24826 13524
rect 7377 13447 7435 13453
rect 7377 13413 7389 13447
rect 7423 13444 7435 13447
rect 7466 13444 7472 13456
rect 7423 13416 7472 13444
rect 7423 13413 7435 13416
rect 7377 13407 7435 13413
rect 7466 13404 7472 13416
rect 7524 13404 7530 13456
rect 8018 13444 8024 13456
rect 7979 13416 8024 13444
rect 8018 13404 8024 13416
rect 8076 13404 8082 13456
rect 13541 13447 13599 13453
rect 13541 13413 13553 13447
rect 13587 13444 13599 13447
rect 13814 13444 13820 13456
rect 13587 13416 13820 13444
rect 13587 13413 13599 13416
rect 13541 13407 13599 13413
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 14642 13444 14648 13456
rect 14603 13416 14648 13444
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1946 13376 1952 13388
rect 1443 13348 1952 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2280 13348 2513 13376
rect 2280 13336 2286 13348
rect 2501 13345 2513 13348
rect 2547 13376 2559 13379
rect 3053 13379 3111 13385
rect 3053 13376 3065 13379
rect 2547 13348 3065 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 3053 13345 3065 13348
rect 3099 13345 3111 13379
rect 3053 13339 3111 13345
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4522 13385 4528 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4212 13348 4261 13376
rect 4212 13336 4218 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 4516 13339 4528 13385
rect 4580 13376 4586 13388
rect 7009 13379 7067 13385
rect 4580 13348 4616 13376
rect 4522 13336 4528 13339
rect 4580 13336 4586 13348
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7929 13379 7987 13385
rect 7929 13376 7941 13379
rect 7055 13348 7941 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7929 13345 7941 13348
rect 7975 13376 7987 13379
rect 8202 13376 8208 13388
rect 7975 13348 8208 13376
rect 7975 13345 7987 13348
rect 7929 13339 7987 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 10778 13336 10784 13388
rect 10836 13376 10842 13388
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 10836 13348 11161 13376
rect 10836 13336 10842 13348
rect 11149 13345 11161 13348
rect 11195 13345 11207 13379
rect 12618 13376 12624 13388
rect 12579 13348 12624 13376
rect 11149 13339 11207 13345
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 13998 13376 14004 13388
rect 13959 13348 14004 13376
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 14093 13379 14151 13385
rect 14093 13345 14105 13379
rect 14139 13376 14151 13379
rect 14550 13376 14556 13388
rect 14139 13348 14556 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 14550 13336 14556 13348
rect 14608 13336 14614 13388
rect 16476 13379 16534 13385
rect 16476 13345 16488 13379
rect 16522 13376 16534 13379
rect 16942 13376 16948 13388
rect 16522 13348 16948 13376
rect 16522 13345 16534 13348
rect 16476 13339 16534 13345
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 18966 13336 18972 13388
rect 19024 13376 19030 13388
rect 19061 13379 19119 13385
rect 19061 13376 19073 13379
rect 19024 13348 19073 13376
rect 19024 13336 19030 13348
rect 19061 13345 19073 13348
rect 19107 13376 19119 13379
rect 19705 13379 19763 13385
rect 19705 13376 19717 13379
rect 19107 13348 19717 13376
rect 19107 13345 19119 13348
rect 19061 13339 19119 13345
rect 19705 13345 19717 13348
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 23569 13379 23627 13385
rect 23569 13376 23581 13379
rect 23532 13348 23581 13376
rect 23532 13336 23538 13348
rect 23569 13345 23581 13348
rect 23615 13345 23627 13379
rect 23569 13339 23627 13345
rect 24581 13379 24639 13385
rect 24581 13345 24593 13379
rect 24627 13376 24639 13379
rect 24670 13376 24676 13388
rect 24627 13348 24676 13376
rect 24627 13345 24639 13348
rect 24581 13339 24639 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2682 13308 2688 13320
rect 2455 13280 2688 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 8628 13280 9689 13308
rect 8628 13268 8634 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 11422 13308 11428 13320
rect 11335 13280 11428 13308
rect 9677 13271 9735 13277
rect 11422 13268 11428 13280
rect 11480 13308 11486 13320
rect 11790 13308 11796 13320
rect 11480 13280 11796 13308
rect 11480 13268 11486 13280
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14826 13308 14832 13320
rect 14323 13280 14832 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15896 13280 16221 13308
rect 15896 13268 15902 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 18598 13268 18604 13320
rect 18656 13308 18662 13320
rect 19153 13311 19211 13317
rect 19153 13308 19165 13311
rect 18656 13280 19165 13308
rect 18656 13268 18662 13280
rect 19153 13277 19165 13280
rect 19199 13277 19211 13311
rect 19153 13271 19211 13277
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13308 20959 13311
rect 21174 13308 21180 13320
rect 20947 13280 21180 13308
rect 20947 13277 20959 13280
rect 20901 13271 20959 13277
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 1949 13243 2007 13249
rect 1949 13240 1961 13243
rect 1452 13212 1961 13240
rect 1452 13200 1458 13212
rect 1949 13209 1961 13212
rect 1995 13209 2007 13243
rect 1949 13203 2007 13209
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 15746 13240 15752 13252
rect 10008 13212 15752 13240
rect 10008 13200 10014 13212
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 3510 13172 3516 13184
rect 3471 13144 3516 13172
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 3786 13172 3792 13184
rect 3747 13144 3792 13172
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 12802 13172 12808 13184
rect 12763 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13078 13172 13084 13184
rect 13039 13144 13084 13172
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 16117 13175 16175 13181
rect 16117 13141 16129 13175
rect 16163 13172 16175 13175
rect 17494 13172 17500 13184
rect 16163 13144 17500 13172
rect 16163 13141 16175 13144
rect 16117 13135 16175 13141
rect 17494 13132 17500 13144
rect 17552 13172 17558 13184
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 17552 13144 17601 13172
rect 17552 13132 17558 13144
rect 17589 13141 17601 13144
rect 17635 13141 17647 13175
rect 18506 13172 18512 13184
rect 18467 13144 18512 13172
rect 17589 13135 17647 13141
rect 18506 13132 18512 13144
rect 18564 13172 18570 13184
rect 19260 13172 19288 13271
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 22554 13308 22560 13320
rect 22515 13280 22560 13308
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 18564 13144 19288 13172
rect 18564 13132 18570 13144
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 3142 12968 3148 12980
rect 3103 12940 3148 12968
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 4246 12968 4252 12980
rect 4207 12940 4252 12968
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 7742 12968 7748 12980
rect 6687 12940 7748 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 7742 12928 7748 12940
rect 7800 12968 7806 12980
rect 8018 12968 8024 12980
rect 7800 12940 8024 12968
rect 7800 12928 7806 12940
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 8202 12968 8208 12980
rect 8163 12940 8208 12968
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 11241 12971 11299 12977
rect 11241 12937 11253 12971
rect 11287 12968 11299 12971
rect 11514 12968 11520 12980
rect 11287 12940 11520 12968
rect 11287 12937 11299 12940
rect 11241 12931 11299 12937
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13814 12968 13820 12980
rect 13727 12940 13820 12968
rect 13814 12928 13820 12940
rect 13872 12968 13878 12980
rect 13998 12968 14004 12980
rect 13872 12940 14004 12968
rect 13872 12928 13878 12940
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15804 12940 16037 12968
rect 15804 12928 15810 12940
rect 16025 12937 16037 12940
rect 16071 12968 16083 12971
rect 16117 12971 16175 12977
rect 16117 12968 16129 12971
rect 16071 12940 16129 12968
rect 16071 12937 16083 12940
rect 16025 12931 16083 12937
rect 16117 12937 16129 12940
rect 16163 12937 16175 12971
rect 16298 12968 16304 12980
rect 16259 12940 16304 12968
rect 16117 12931 16175 12937
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23532 12940 23857 12968
rect 23532 12928 23538 12940
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 23934 12928 23940 12980
rect 23992 12968 23998 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 23992 12940 24777 12968
rect 23992 12928 23998 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 4709 12903 4767 12909
rect 4709 12900 4721 12903
rect 3620 12872 4721 12900
rect 3510 12792 3516 12844
rect 3568 12832 3574 12844
rect 3620 12841 3648 12872
rect 4709 12869 4721 12872
rect 4755 12869 4767 12903
rect 4709 12863 4767 12869
rect 7377 12903 7435 12909
rect 7377 12869 7389 12903
rect 7423 12900 7435 12903
rect 8110 12900 8116 12912
rect 7423 12872 8116 12900
rect 7423 12869 7435 12872
rect 7377 12863 7435 12869
rect 8110 12860 8116 12872
rect 8168 12860 8174 12912
rect 10778 12900 10784 12912
rect 10739 12872 10784 12900
rect 10778 12860 10784 12872
rect 10836 12860 10842 12912
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 11388 12872 13093 12900
rect 11388 12860 11394 12872
rect 13081 12869 13093 12872
rect 13127 12869 13139 12903
rect 13081 12863 13139 12869
rect 18049 12903 18107 12909
rect 18049 12869 18061 12903
rect 18095 12869 18107 12903
rect 18049 12863 18107 12869
rect 19613 12903 19671 12909
rect 19613 12869 19625 12903
rect 19659 12900 19671 12903
rect 22741 12903 22799 12909
rect 19659 12872 22600 12900
rect 19659 12869 19671 12872
rect 19613 12863 19671 12869
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3568 12804 3617 12832
rect 3568 12792 3574 12804
rect 3605 12801 3617 12804
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3786 12832 3792 12844
rect 3743 12804 3792 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1854 12764 1860 12776
rect 1443 12736 1860 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3712 12764 3740 12795
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4522 12792 4528 12844
rect 4580 12832 4586 12844
rect 5166 12832 5172 12844
rect 4580 12804 5172 12832
rect 4580 12792 4586 12804
rect 5166 12792 5172 12804
rect 5224 12832 5230 12844
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 5224 12804 5273 12832
rect 5224 12792 5230 12804
rect 5261 12801 5273 12804
rect 5307 12832 5319 12835
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5307 12804 5733 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8662 12832 8668 12844
rect 8444 12804 8668 12832
rect 8444 12792 8450 12804
rect 8662 12792 8668 12804
rect 8720 12832 8726 12844
rect 8757 12835 8815 12841
rect 8757 12832 8769 12835
rect 8720 12804 8769 12832
rect 8720 12792 8726 12804
rect 8757 12801 8769 12804
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 9916 12804 10333 12832
rect 9916 12792 9922 12804
rect 10321 12801 10333 12804
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 13906 12832 13912 12844
rect 12400 12804 13912 12832
rect 12400 12792 12406 12804
rect 13906 12792 13912 12804
rect 13964 12832 13970 12844
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 13964 12804 14381 12832
rect 13964 12792 13970 12804
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14884 12804 14933 12832
rect 14884 12792 14890 12804
rect 14921 12801 14933 12804
rect 14967 12832 14979 12835
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 14967 12804 15485 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 15473 12801 15485 12804
rect 15519 12832 15531 12835
rect 16942 12832 16948 12844
rect 15519 12804 16948 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 16942 12792 16948 12804
rect 17000 12832 17006 12844
rect 17313 12835 17371 12841
rect 17313 12832 17325 12835
rect 17000 12804 17325 12832
rect 17000 12792 17006 12804
rect 17313 12801 17325 12804
rect 17359 12801 17371 12835
rect 17313 12795 17371 12801
rect 4614 12764 4620 12776
rect 3099 12736 3740 12764
rect 4527 12736 4620 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 4614 12724 4620 12736
rect 4672 12764 4678 12776
rect 5074 12764 5080 12776
rect 4672 12736 5080 12764
rect 4672 12724 4678 12736
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 8570 12764 8576 12776
rect 7791 12736 8576 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 9306 12764 9312 12776
rect 9219 12736 9312 12764
rect 9306 12724 9312 12736
rect 9364 12764 9370 12776
rect 10686 12764 10692 12776
rect 9364 12736 10692 12764
rect 9364 12724 9370 12736
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 11333 12767 11391 12773
rect 11333 12733 11345 12767
rect 11379 12764 11391 12767
rect 12805 12767 12863 12773
rect 11379 12736 12296 12764
rect 11379 12733 11391 12736
rect 11333 12727 11391 12733
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 3513 12699 3571 12705
rect 3513 12696 3525 12699
rect 3476 12668 3525 12696
rect 3476 12656 3482 12668
rect 3513 12665 3525 12668
rect 3559 12696 3571 12699
rect 4246 12696 4252 12708
rect 3559 12668 4252 12696
rect 3559 12665 3571 12668
rect 3513 12659 3571 12665
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 4798 12656 4804 12708
rect 4856 12696 4862 12708
rect 5169 12699 5227 12705
rect 5169 12696 5181 12699
rect 4856 12668 5181 12696
rect 4856 12656 4862 12668
rect 5169 12665 5181 12668
rect 5215 12665 5227 12699
rect 5169 12659 5227 12665
rect 8113 12699 8171 12705
rect 8113 12665 8125 12699
rect 8159 12696 8171 12699
rect 8665 12699 8723 12705
rect 8665 12696 8677 12699
rect 8159 12668 8677 12696
rect 8159 12665 8171 12668
rect 8113 12659 8171 12665
rect 8665 12665 8677 12668
rect 8711 12696 8723 12699
rect 8754 12696 8760 12708
rect 8711 12668 8760 12696
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 8754 12656 8760 12668
rect 8812 12656 8818 12708
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 10137 12699 10195 12705
rect 10137 12696 10149 12699
rect 9723 12668 10149 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 10137 12665 10149 12668
rect 10183 12696 10195 12699
rect 11606 12696 11612 12708
rect 10183 12668 11612 12696
rect 10183 12665 10195 12668
rect 10137 12659 10195 12665
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 12268 12640 12296 12736
rect 12805 12733 12817 12767
rect 12851 12764 12863 12767
rect 13078 12764 13084 12776
rect 12851 12736 13084 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 13078 12724 13084 12736
rect 13136 12764 13142 12776
rect 13630 12764 13636 12776
rect 13136 12736 13636 12764
rect 13136 12724 13142 12736
rect 13630 12724 13636 12736
rect 13688 12724 13694 12776
rect 13725 12767 13783 12773
rect 13725 12733 13737 12767
rect 13771 12764 13783 12767
rect 14090 12764 14096 12776
rect 13771 12736 14096 12764
rect 13771 12733 13783 12736
rect 13725 12727 13783 12733
rect 14090 12724 14096 12736
rect 14148 12764 14154 12776
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 14148 12736 14197 12764
rect 14148 12724 14154 12736
rect 14185 12733 14197 12736
rect 14231 12764 14243 12767
rect 16482 12764 16488 12776
rect 14231 12736 16488 12764
rect 14231 12733 14243 12736
rect 14185 12727 14243 12733
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 16669 12767 16727 12773
rect 16669 12764 16681 12767
rect 16632 12736 16681 12764
rect 16632 12724 16638 12736
rect 16669 12733 16681 12736
rect 16715 12764 16727 12767
rect 17402 12764 17408 12776
rect 16715 12736 17408 12764
rect 16715 12733 16727 12736
rect 16669 12727 16727 12733
rect 17402 12724 17408 12736
rect 17460 12724 17466 12776
rect 18064 12764 18092 12863
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18564 12804 18613 12832
rect 18564 12792 18570 12804
rect 18601 12801 18613 12804
rect 18647 12832 18659 12835
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18647 12804 19073 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 20070 12832 20076 12844
rect 20031 12804 20076 12832
rect 19061 12795 19119 12801
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12832 20223 12835
rect 20211 12804 20392 12832
rect 20211 12801 20223 12804
rect 20165 12795 20223 12801
rect 19981 12767 20039 12773
rect 19981 12764 19993 12767
rect 18064 12736 19993 12764
rect 19981 12733 19993 12736
rect 20027 12764 20039 12767
rect 20254 12764 20260 12776
rect 20027 12736 20260 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 12713 12699 12771 12705
rect 12713 12696 12725 12699
rect 12676 12668 12725 12696
rect 12676 12656 12682 12668
rect 12713 12665 12725 12668
rect 12759 12696 12771 12699
rect 13354 12696 13360 12708
rect 12759 12668 13360 12696
rect 12759 12665 12771 12668
rect 12713 12659 12771 12665
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 15286 12656 15292 12708
rect 15344 12696 15350 12708
rect 17773 12699 17831 12705
rect 17773 12696 17785 12699
rect 15344 12668 17785 12696
rect 15344 12656 15350 12668
rect 17773 12665 17785 12668
rect 17819 12696 17831 12699
rect 18417 12699 18475 12705
rect 18417 12696 18429 12699
rect 17819 12668 18429 12696
rect 17819 12665 17831 12668
rect 17773 12659 17831 12665
rect 18417 12665 18429 12668
rect 18463 12665 18475 12699
rect 18417 12659 18475 12665
rect 18506 12656 18512 12708
rect 18564 12696 18570 12708
rect 19518 12696 19524 12708
rect 18564 12668 19196 12696
rect 19479 12668 19524 12696
rect 18564 12656 18570 12668
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2958 12628 2964 12640
rect 2547 12600 2964 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12628 9827 12631
rect 9950 12628 9956 12640
rect 9815 12600 9956 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10686 12628 10692 12640
rect 10275 12600 10692 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11296 12600 11529 12628
rect 11296 12588 11302 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 12250 12628 12256 12640
rect 12211 12600 12256 12628
rect 11517 12591 11575 12597
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12986 12628 12992 12640
rect 12947 12600 12992 12628
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13081 12631 13139 12637
rect 13081 12597 13093 12631
rect 13127 12628 13139 12631
rect 13265 12631 13323 12637
rect 13265 12628 13277 12631
rect 13127 12600 13277 12628
rect 13127 12597 13139 12600
rect 13081 12591 13139 12597
rect 13265 12597 13277 12600
rect 13311 12628 13323 12631
rect 14277 12631 14335 12637
rect 14277 12628 14289 12631
rect 13311 12600 14289 12628
rect 13311 12597 13323 12600
rect 13265 12591 13323 12597
rect 14277 12597 14289 12600
rect 14323 12628 14335 12631
rect 15378 12628 15384 12640
rect 14323 12600 15384 12628
rect 14323 12597 14335 12600
rect 14277 12591 14335 12597
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 15838 12628 15844 12640
rect 15799 12600 15844 12628
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 16025 12631 16083 12637
rect 16025 12597 16037 12631
rect 16071 12628 16083 12631
rect 16758 12628 16764 12640
rect 16071 12600 16764 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 19168 12628 19196 12668
rect 19518 12656 19524 12668
rect 19576 12696 19582 12708
rect 20364 12696 20392 12804
rect 22572 12773 22600 12872
rect 22741 12869 22753 12903
rect 22787 12900 22799 12903
rect 24397 12903 24455 12909
rect 24397 12900 24409 12903
rect 22787 12872 24409 12900
rect 22787 12869 22799 12872
rect 22741 12863 22799 12869
rect 24397 12869 24409 12872
rect 24443 12900 24455 12903
rect 24670 12900 24676 12912
rect 24443 12872 24676 12900
rect 24443 12869 24455 12872
rect 24397 12863 24455 12869
rect 24670 12860 24676 12872
rect 24728 12860 24734 12912
rect 22549 12767 22607 12773
rect 22549 12733 22561 12767
rect 22595 12733 22607 12767
rect 22549 12727 22607 12733
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 24670 12764 24676 12776
rect 24627 12736 24676 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 19576 12668 20392 12696
rect 22572 12696 22600 12727
rect 24670 12724 24676 12736
rect 24728 12764 24734 12776
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24728 12736 25145 12764
rect 24728 12724 24734 12736
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 23017 12699 23075 12705
rect 23017 12696 23029 12699
rect 22572 12668 23029 12696
rect 19576 12656 19582 12668
rect 23017 12665 23029 12668
rect 23063 12665 23075 12699
rect 23017 12659 23075 12665
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 19168 12600 20729 12628
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 20717 12591 20775 12597
rect 21177 12631 21235 12637
rect 21177 12597 21189 12631
rect 21223 12628 21235 12631
rect 21358 12628 21364 12640
rect 21223 12600 21364 12628
rect 21223 12597 21235 12600
rect 21177 12591 21235 12597
rect 21358 12588 21364 12600
rect 21416 12588 21422 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 2314 12424 2320 12436
rect 1627 12396 2320 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 2590 12424 2596 12436
rect 2455 12396 2596 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4430 12424 4436 12436
rect 4295 12396 4436 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 7742 12424 7748 12436
rect 7703 12396 7748 12424
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 14185 12427 14243 12433
rect 14185 12424 14197 12427
rect 13964 12396 14197 12424
rect 13964 12384 13970 12396
rect 14185 12393 14197 12396
rect 14231 12393 14243 12427
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 14185 12387 14243 12393
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 16022 12384 16028 12436
rect 16080 12424 16086 12436
rect 16117 12427 16175 12433
rect 16117 12424 16129 12427
rect 16080 12396 16129 12424
rect 16080 12384 16086 12396
rect 16117 12393 16129 12396
rect 16163 12393 16175 12427
rect 16574 12424 16580 12436
rect 16535 12396 16580 12424
rect 16117 12387 16175 12393
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18690 12424 18696 12436
rect 18104 12396 18696 12424
rect 18104 12384 18110 12396
rect 18690 12384 18696 12396
rect 18748 12424 18754 12436
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 18748 12396 19625 12424
rect 18748 12384 18754 12396
rect 19613 12393 19625 12396
rect 19659 12393 19671 12427
rect 20254 12424 20260 12436
rect 20215 12396 20260 12424
rect 19613 12387 19671 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 24026 12384 24032 12436
rect 24084 12424 24090 12436
rect 24765 12427 24823 12433
rect 24765 12424 24777 12427
rect 24084 12396 24777 12424
rect 24084 12384 24090 12396
rect 24765 12393 24777 12396
rect 24811 12393 24823 12427
rect 24765 12387 24823 12393
rect 2777 12359 2835 12365
rect 2777 12325 2789 12359
rect 2823 12356 2835 12359
rect 2866 12356 2872 12368
rect 2823 12328 2872 12356
rect 2823 12325 2835 12328
rect 2777 12319 2835 12325
rect 2866 12316 2872 12328
rect 2924 12356 2930 12368
rect 3326 12356 3332 12368
rect 2924 12328 3332 12356
rect 2924 12316 2930 12328
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 5629 12359 5687 12365
rect 5629 12325 5641 12359
rect 5675 12356 5687 12359
rect 6178 12356 6184 12368
rect 5675 12328 6184 12356
rect 5675 12325 5687 12328
rect 5629 12319 5687 12325
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 11572 12328 13768 12356
rect 11572 12316 11578 12328
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 2682 12288 2688 12300
rect 1443 12260 2688 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 3418 12288 3424 12300
rect 2884 12260 3424 12288
rect 2884 12229 2912 12260
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 6086 12288 6092 12300
rect 5767 12260 6092 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 6086 12248 6092 12260
rect 6144 12288 6150 12300
rect 6362 12288 6368 12300
rect 6144 12260 6368 12288
rect 6144 12248 6150 12260
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12288 7343 12291
rect 8110 12288 8116 12300
rect 7331 12260 8116 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 10502 12288 10508 12300
rect 10463 12260 10508 12288
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 10761 12291 10819 12297
rect 10761 12288 10773 12291
rect 10612 12260 10773 12288
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 5074 12220 5080 12232
rect 3016 12192 5080 12220
rect 3016 12180 3022 12192
rect 5074 12180 5080 12192
rect 5132 12220 5138 12232
rect 5813 12223 5871 12229
rect 5132 12192 5672 12220
rect 5132 12180 5138 12192
rect 3326 12112 3332 12164
rect 3384 12152 3390 12164
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 3384 12124 3801 12152
rect 3384 12112 3390 12124
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 5261 12155 5319 12161
rect 5261 12152 5273 12155
rect 4304 12124 5273 12152
rect 4304 12112 4310 12124
rect 5261 12121 5273 12124
rect 5307 12121 5319 12155
rect 5644 12152 5672 12192
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 7653 12223 7711 12229
rect 7653 12189 7665 12223
rect 7699 12220 7711 12223
rect 7926 12220 7932 12232
rect 7699 12192 7932 12220
rect 7699 12189 7711 12192
rect 7653 12183 7711 12189
rect 5828 12152 5856 12183
rect 7926 12180 7932 12192
rect 7984 12220 7990 12232
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 7984 12192 8217 12220
rect 7984 12180 7990 12192
rect 8205 12189 8217 12192
rect 8251 12189 8263 12223
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 8205 12183 8263 12189
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10612 12220 10640 12260
rect 10761 12257 10773 12260
rect 10807 12288 10819 12291
rect 12066 12288 12072 12300
rect 10807 12260 12072 12288
rect 10807 12257 10819 12260
rect 10761 12251 10819 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 13538 12288 13544 12300
rect 13499 12260 13544 12288
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 13740 12288 13768 12328
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 14921 12359 14979 12365
rect 14921 12356 14933 12359
rect 13872 12328 14933 12356
rect 13872 12316 13878 12328
rect 14921 12325 14933 12328
rect 14967 12325 14979 12359
rect 14921 12319 14979 12325
rect 18874 12316 18880 12368
rect 18932 12356 18938 12368
rect 19242 12356 19248 12368
rect 18932 12328 19248 12356
rect 18932 12316 18938 12328
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 22278 12356 22284 12368
rect 21928 12328 22284 12356
rect 14182 12288 14188 12300
rect 13740 12260 14188 12288
rect 14182 12248 14188 12260
rect 14240 12248 14246 12300
rect 17028 12291 17086 12297
rect 17028 12257 17040 12291
rect 17074 12288 17086 12291
rect 17494 12288 17500 12300
rect 17074 12260 17500 12288
rect 17074 12257 17086 12260
rect 17028 12251 17086 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 19058 12288 19064 12300
rect 19019 12260 19064 12288
rect 19058 12248 19064 12260
rect 19116 12288 19122 12300
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19116 12260 19717 12288
rect 19116 12248 19122 12260
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 21928 12297 21956 12328
rect 22278 12316 22284 12328
rect 22336 12316 22342 12368
rect 21913 12291 21971 12297
rect 21913 12288 21925 12291
rect 20772 12260 21925 12288
rect 20772 12248 20778 12260
rect 21913 12257 21925 12260
rect 21959 12257 21971 12291
rect 21913 12251 21971 12257
rect 22002 12248 22008 12300
rect 22060 12288 22066 12300
rect 22169 12291 22227 12297
rect 22169 12288 22181 12291
rect 22060 12260 22181 12288
rect 22060 12248 22066 12260
rect 22169 12257 22181 12260
rect 22215 12257 22227 12291
rect 22169 12251 22227 12257
rect 24210 12248 24216 12300
rect 24268 12288 24274 12300
rect 24581 12291 24639 12297
rect 24581 12288 24593 12291
rect 24268 12260 24593 12288
rect 24268 12248 24274 12260
rect 24581 12257 24593 12260
rect 24627 12257 24639 12291
rect 24581 12251 24639 12257
rect 9732 12192 10640 12220
rect 9732 12180 9738 12192
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 13633 12223 13691 12229
rect 13633 12220 13645 12223
rect 13136 12192 13645 12220
rect 13136 12180 13142 12192
rect 13633 12189 13645 12192
rect 13679 12189 13691 12223
rect 13633 12183 13691 12189
rect 13817 12223 13875 12229
rect 13817 12189 13829 12223
rect 13863 12220 13875 12223
rect 13906 12220 13912 12232
rect 13863 12192 13912 12220
rect 13863 12189 13875 12192
rect 13817 12183 13875 12189
rect 5644 12124 5856 12152
rect 5261 12115 5319 12121
rect 7466 12112 7472 12164
rect 7524 12152 7530 12164
rect 9858 12152 9864 12164
rect 7524 12124 9864 12152
rect 7524 12112 7530 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 11514 12112 11520 12164
rect 11572 12152 11578 12164
rect 11885 12155 11943 12161
rect 11885 12152 11897 12155
rect 11572 12124 11897 12152
rect 11572 12112 11578 12124
rect 11885 12121 11897 12124
rect 11931 12121 11943 12155
rect 11885 12115 11943 12121
rect 12989 12155 13047 12161
rect 12989 12121 13001 12155
rect 13035 12152 13047 12155
rect 13832 12152 13860 12183
rect 13906 12180 13912 12192
rect 13964 12180 13970 12232
rect 14550 12220 14556 12232
rect 14511 12192 14556 12220
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16758 12220 16764 12232
rect 15896 12192 16764 12220
rect 15896 12180 15902 12192
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 18984 12192 19809 12220
rect 13035 12124 13860 12152
rect 13035 12121 13047 12124
rect 12989 12115 13047 12121
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 2314 12084 2320 12096
rect 2275 12056 2320 12084
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 3421 12087 3479 12093
rect 3421 12084 3433 12087
rect 3292 12056 3433 12084
rect 3292 12044 3298 12056
rect 3421 12053 3433 12056
rect 3467 12053 3479 12087
rect 4798 12084 4804 12096
rect 4759 12056 4804 12084
rect 3421 12047 3479 12053
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 6270 12084 6276 12096
rect 6231 12056 6276 12084
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 6638 12084 6644 12096
rect 6599 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 13170 12084 13176 12096
rect 13131 12056 13176 12084
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 18141 12087 18199 12093
rect 18141 12084 18153 12087
rect 18012 12056 18153 12084
rect 18012 12044 18018 12056
rect 18141 12053 18153 12056
rect 18187 12053 18199 12087
rect 18141 12047 18199 12053
rect 18598 12044 18604 12096
rect 18656 12084 18662 12096
rect 18693 12087 18751 12093
rect 18693 12084 18705 12087
rect 18656 12056 18705 12084
rect 18656 12044 18662 12056
rect 18693 12053 18705 12056
rect 18739 12053 18751 12087
rect 18984 12084 19012 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 20901 12223 20959 12229
rect 20901 12189 20913 12223
rect 20947 12220 20959 12223
rect 21266 12220 21272 12232
rect 20947 12192 21272 12220
rect 20947 12189 20959 12192
rect 20901 12183 20959 12189
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 19058 12084 19064 12096
rect 18984 12056 19064 12084
rect 18693 12047 18751 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19242 12084 19248 12096
rect 19203 12056 19248 12084
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 21361 12087 21419 12093
rect 21361 12084 21373 12087
rect 21048 12056 21373 12084
rect 21048 12044 21054 12056
rect 21361 12053 21373 12056
rect 21407 12053 21419 12087
rect 21361 12047 21419 12053
rect 21821 12087 21879 12093
rect 21821 12053 21833 12087
rect 21867 12084 21879 12087
rect 21910 12084 21916 12096
rect 21867 12056 21916 12084
rect 21867 12053 21879 12056
rect 21821 12047 21879 12053
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 23293 12087 23351 12093
rect 23293 12053 23305 12087
rect 23339 12084 23351 12087
rect 23934 12084 23940 12096
rect 23339 12056 23940 12084
rect 23339 12053 23351 12056
rect 23293 12047 23351 12053
rect 23934 12044 23940 12056
rect 23992 12044 23998 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11880 1823 11883
rect 2866 11880 2872 11892
rect 1811 11852 2872 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11880 3387 11883
rect 3418 11880 3424 11892
rect 3375 11852 3424 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 5132 11852 5181 11880
rect 5132 11840 5138 11852
rect 5169 11849 5181 11852
rect 5215 11880 5227 11883
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5215 11852 6469 11880
rect 5215 11849 5227 11852
rect 5169 11843 5227 11849
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7101 11883 7159 11889
rect 7101 11880 7113 11883
rect 7064 11852 7113 11880
rect 7064 11840 7070 11852
rect 7101 11849 7113 11852
rect 7147 11849 7159 11883
rect 7101 11843 7159 11849
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2777 11747 2835 11753
rect 2777 11744 2789 11747
rect 2372 11716 2789 11744
rect 2372 11704 2378 11716
rect 2777 11713 2789 11716
rect 2823 11713 2835 11747
rect 7116 11744 7144 11843
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 8444 11852 9229 11880
rect 8444 11840 8450 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9674 11880 9680 11892
rect 9635 11852 9680 11880
rect 9217 11843 9275 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 10778 11880 10784 11892
rect 10739 11852 10784 11880
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 12342 11880 12348 11892
rect 11931 11852 12348 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7116 11716 7297 11744
rect 2777 11707 2835 11713
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 11425 11747 11483 11753
rect 9732 11716 10272 11744
rect 9732 11704 9738 11716
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3743 11648 3801 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 3789 11645 3801 11648
rect 3835 11676 3847 11679
rect 4338 11676 4344 11688
rect 3835 11648 4344 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 7374 11636 7380 11688
rect 7432 11676 7438 11688
rect 7552 11679 7610 11685
rect 7552 11676 7564 11679
rect 7432 11648 7564 11676
rect 7432 11636 7438 11648
rect 7552 11645 7564 11648
rect 7598 11676 7610 11679
rect 7834 11676 7840 11688
rect 7598 11648 7840 11676
rect 7598 11645 7610 11648
rect 7552 11639 7610 11645
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 9769 11679 9827 11685
rect 9769 11645 9781 11679
rect 9815 11676 9827 11679
rect 10134 11676 10140 11688
rect 9815 11648 10140 11676
rect 9815 11645 9827 11648
rect 9769 11639 9827 11645
rect 10134 11636 10140 11648
rect 10192 11636 10198 11688
rect 10244 11676 10272 11716
rect 11425 11713 11437 11747
rect 11471 11744 11483 11747
rect 11900 11744 11928 11843
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11880 13323 11883
rect 13538 11880 13544 11892
rect 13311 11852 13544 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 16114 11880 16120 11892
rect 16075 11852 16120 11880
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 21726 11840 21732 11892
rect 21784 11880 21790 11892
rect 22002 11880 22008 11892
rect 21784 11852 22008 11880
rect 21784 11840 21790 11852
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 22278 11840 22284 11892
rect 22336 11880 22342 11892
rect 22833 11883 22891 11889
rect 22833 11880 22845 11883
rect 22336 11852 22845 11880
rect 22336 11840 22342 11852
rect 22833 11849 22845 11852
rect 22879 11880 22891 11883
rect 23385 11883 23443 11889
rect 23385 11880 23397 11883
rect 22879 11852 23397 11880
rect 22879 11849 22891 11852
rect 22833 11843 22891 11849
rect 23385 11849 23397 11852
rect 23431 11880 23443 11883
rect 24026 11880 24032 11892
rect 23431 11852 24032 11880
rect 23431 11849 23443 11852
rect 23385 11843 23443 11849
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 14734 11772 14740 11824
rect 14792 11812 14798 11824
rect 18785 11815 18843 11821
rect 18785 11812 18797 11815
rect 14792 11784 18797 11812
rect 14792 11772 14798 11784
rect 18785 11781 18797 11784
rect 18831 11812 18843 11815
rect 19058 11812 19064 11824
rect 18831 11784 19064 11812
rect 18831 11781 18843 11784
rect 18785 11775 18843 11781
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 20990 11772 20996 11824
rect 21048 11812 21054 11824
rect 21048 11784 22212 11812
rect 21048 11772 21054 11784
rect 11471 11716 11928 11744
rect 11471 11713 11483 11716
rect 11425 11707 11483 11713
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16577 11747 16635 11753
rect 16577 11744 16589 11747
rect 16080 11716 16589 11744
rect 16080 11704 16086 11716
rect 16577 11713 16589 11716
rect 16623 11713 16635 11747
rect 16577 11707 16635 11713
rect 16761 11747 16819 11753
rect 16761 11713 16773 11747
rect 16807 11744 16819 11747
rect 17954 11744 17960 11756
rect 16807 11716 17960 11744
rect 16807 11713 16819 11716
rect 16761 11707 16819 11713
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 10244 11648 12449 11676
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 13446 11676 13452 11688
rect 12584 11648 13452 11676
rect 12584 11636 12590 11648
rect 13446 11636 13452 11648
rect 13504 11676 13510 11688
rect 13906 11685 13912 11688
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13504 11648 13645 11676
rect 13504 11636 13510 11648
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13900 11676 13912 11685
rect 13819 11648 13912 11676
rect 13633 11639 13691 11645
rect 13900 11639 13912 11648
rect 13964 11676 13970 11688
rect 14642 11676 14648 11688
rect 13964 11648 14648 11676
rect 2685 11611 2743 11617
rect 2685 11608 2697 11611
rect 2056 11580 2697 11608
rect 2056 11552 2084 11580
rect 2685 11577 2697 11580
rect 2731 11577 2743 11611
rect 2685 11571 2743 11577
rect 3970 11568 3976 11620
rect 4028 11617 4034 11620
rect 4028 11611 4092 11617
rect 4028 11577 4046 11611
rect 4080 11577 4092 11611
rect 4028 11571 4092 11577
rect 5813 11611 5871 11617
rect 5813 11577 5825 11611
rect 5859 11608 5871 11611
rect 6086 11608 6092 11620
rect 5859 11580 6092 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 4028 11568 4034 11571
rect 6086 11568 6092 11580
rect 6144 11568 6150 11620
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 10735 11580 11161 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 11149 11577 11161 11580
rect 11195 11608 11207 11611
rect 11514 11608 11520 11620
rect 11195 11580 11520 11608
rect 11195 11577 11207 11580
rect 11149 11571 11207 11577
rect 11514 11568 11520 11580
rect 11572 11608 11578 11620
rect 11974 11608 11980 11620
rect 11572 11580 11980 11608
rect 11572 11568 11578 11580
rect 11974 11568 11980 11580
rect 12032 11568 12038 11620
rect 13648 11608 13676 11639
rect 13906 11636 13912 11639
rect 13964 11636 13970 11648
rect 14642 11636 14648 11648
rect 14700 11676 14706 11688
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 14700 11648 15669 11676
rect 14700 11636 14706 11648
rect 15657 11645 15669 11648
rect 15703 11676 15715 11679
rect 16776 11676 16804 11707
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 22184 11744 22212 11784
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 22184 11716 22385 11744
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 15703 11648 16804 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 17920 11648 19165 11676
rect 17920 11636 17926 11648
rect 19153 11645 19165 11648
rect 19199 11676 19211 11679
rect 19337 11679 19395 11685
rect 19337 11676 19349 11679
rect 19199 11648 19349 11676
rect 19199 11645 19211 11648
rect 19153 11639 19211 11645
rect 19337 11645 19349 11648
rect 19383 11676 19395 11679
rect 20714 11676 20720 11688
rect 19383 11648 20720 11676
rect 19383 11645 19395 11648
rect 19337 11639 19395 11645
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 22189 11679 22247 11685
rect 22189 11676 22201 11679
rect 21652 11648 22201 11676
rect 14274 11608 14280 11620
rect 13648 11580 14280 11608
rect 14274 11568 14280 11580
rect 14332 11568 14338 11620
rect 19518 11568 19524 11620
rect 19576 11617 19582 11620
rect 19576 11611 19640 11617
rect 19576 11577 19594 11611
rect 19628 11577 19640 11611
rect 19576 11571 19640 11577
rect 19576 11568 19582 11571
rect 20346 11568 20352 11620
rect 20404 11608 20410 11620
rect 21652 11617 21680 11648
rect 22189 11645 22201 11648
rect 22235 11676 22247 11679
rect 23661 11679 23719 11685
rect 22235 11648 23520 11676
rect 22235 11645 22247 11648
rect 22189 11639 22247 11645
rect 21637 11611 21695 11617
rect 21637 11608 21649 11611
rect 20404 11580 21649 11608
rect 20404 11568 20410 11580
rect 21637 11577 21649 11580
rect 21683 11577 21695 11611
rect 23492 11608 23520 11648
rect 23661 11645 23673 11679
rect 23707 11676 23719 11679
rect 23707 11648 24072 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 24044 11620 24072 11648
rect 23934 11617 23940 11620
rect 23928 11608 23940 11617
rect 23492 11580 23796 11608
rect 23895 11580 23940 11608
rect 21637 11571 21695 11577
rect 2038 11540 2044 11552
rect 1999 11512 2044 11540
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 2314 11540 2320 11552
rect 2271 11512 2320 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2590 11540 2596 11552
rect 2551 11512 2596 11540
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 6178 11540 6184 11552
rect 6139 11512 6184 11540
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 8352 11512 8677 11540
rect 8352 11500 8358 11512
rect 8665 11509 8677 11512
rect 8711 11509 8723 11543
rect 9950 11540 9956 11552
rect 9911 11512 9956 11540
rect 8665 11503 8723 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 10100 11512 10241 11540
rect 10100 11500 10106 11512
rect 10229 11509 10241 11512
rect 10275 11540 10287 11543
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 10275 11512 11253 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 11241 11509 11253 11512
rect 11287 11540 11299 11543
rect 12434 11540 12440 11552
rect 11287 11512 12440 11540
rect 11287 11509 11299 11512
rect 11241 11503 11299 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 14090 11540 14096 11552
rect 12676 11512 14096 11540
rect 12676 11500 12682 11512
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 15010 11540 15016 11552
rect 14971 11512 15016 11540
rect 15010 11500 15016 11512
rect 15068 11540 15074 11552
rect 15470 11540 15476 11552
rect 15068 11512 15476 11540
rect 15068 11500 15074 11512
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16390 11540 16396 11552
rect 16071 11512 16396 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16390 11500 16396 11512
rect 16448 11540 16454 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 16448 11512 16497 11540
rect 16448 11500 16454 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16485 11503 16543 11509
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 16816 11512 17233 11540
rect 16816 11500 16822 11512
rect 17221 11509 17233 11512
rect 17267 11540 17279 11543
rect 17862 11540 17868 11552
rect 17267 11512 17868 11540
rect 17267 11509 17279 11512
rect 17221 11503 17279 11509
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 20128 11512 20729 11540
rect 20128 11500 20134 11512
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 20717 11503 20775 11509
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21082 11540 21088 11552
rect 20864 11512 21088 11540
rect 20864 11500 20870 11512
rect 21082 11500 21088 11512
rect 21140 11540 21146 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 21140 11512 21281 11540
rect 21140 11500 21146 11512
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21818 11540 21824 11552
rect 21779 11512 21824 11540
rect 21269 11503 21327 11509
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 23474 11540 23480 11552
rect 22336 11512 23480 11540
rect 22336 11500 22342 11512
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 23768 11540 23796 11580
rect 23928 11571 23940 11580
rect 23934 11568 23940 11571
rect 23992 11568 23998 11620
rect 24026 11568 24032 11620
rect 24084 11568 24090 11620
rect 24578 11540 24584 11552
rect 23768 11512 24584 11540
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 25038 11540 25044 11552
rect 24999 11512 25044 11540
rect 25038 11500 25044 11512
rect 25096 11500 25102 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 2222 11336 2228 11348
rect 1627 11308 2228 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2682 11336 2688 11348
rect 2455 11308 2688 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 2832 11308 4077 11336
rect 2832 11296 2838 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 4433 11339 4491 11345
rect 4433 11336 4445 11339
rect 4396 11308 4445 11336
rect 4396 11296 4402 11308
rect 4433 11305 4445 11308
rect 4479 11336 4491 11339
rect 6638 11336 6644 11348
rect 4479 11308 6644 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 7374 11336 7380 11348
rect 7335 11308 7380 11336
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7926 11336 7932 11348
rect 7887 11308 7932 11336
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 12066 11336 12072 11348
rect 12027 11308 12072 11336
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 13078 11336 13084 11348
rect 13039 11308 13084 11336
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 14642 11336 14648 11348
rect 13228 11308 13273 11336
rect 14603 11308 14648 11336
rect 13228 11296 13234 11308
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16540 11308 16681 11336
rect 16540 11296 16546 11308
rect 16669 11305 16681 11308
rect 16715 11336 16727 11339
rect 16850 11336 16856 11348
rect 16715 11308 16856 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19245 11339 19303 11345
rect 19245 11305 19257 11339
rect 19291 11336 19303 11339
rect 20717 11339 20775 11345
rect 20717 11336 20729 11339
rect 19291 11308 20729 11336
rect 19291 11305 19303 11308
rect 19245 11299 19303 11305
rect 20717 11305 20729 11308
rect 20763 11336 20775 11339
rect 21082 11336 21088 11348
rect 20763 11308 21088 11336
rect 20763 11305 20775 11308
rect 20717 11299 20775 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 22554 11296 22560 11348
rect 22612 11336 22618 11348
rect 22833 11339 22891 11345
rect 22833 11336 22845 11339
rect 22612 11308 22845 11336
rect 22612 11296 22618 11308
rect 22833 11305 22845 11308
rect 22879 11305 22891 11339
rect 22833 11299 22891 11305
rect 23109 11339 23167 11345
rect 23109 11305 23121 11339
rect 23155 11336 23167 11339
rect 23845 11339 23903 11345
rect 23845 11336 23857 11339
rect 23155 11308 23857 11336
rect 23155 11305 23167 11308
rect 23109 11299 23167 11305
rect 23845 11305 23857 11308
rect 23891 11336 23903 11339
rect 24854 11336 24860 11348
rect 23891 11308 24860 11336
rect 23891 11305 23903 11308
rect 23845 11299 23903 11305
rect 2866 11228 2872 11280
rect 2924 11268 2930 11280
rect 4525 11271 4583 11277
rect 4525 11268 4537 11271
rect 2924 11240 4537 11268
rect 2924 11228 2930 11240
rect 4525 11237 4537 11240
rect 4571 11268 4583 11271
rect 6270 11268 6276 11280
rect 4571 11240 6276 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 7650 11268 7656 11280
rect 7064 11240 7656 11268
rect 7064 11228 7070 11240
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 8018 11228 8024 11280
rect 8076 11268 8082 11280
rect 8297 11271 8355 11277
rect 8297 11268 8309 11271
rect 8076 11240 8309 11268
rect 8076 11228 8082 11240
rect 8297 11237 8309 11240
rect 8343 11268 8355 11271
rect 8386 11268 8392 11280
rect 8343 11240 8392 11268
rect 8343 11237 8355 11240
rect 8297 11231 8355 11237
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 12434 11268 12440 11280
rect 11664 11240 12440 11268
rect 11664 11228 11670 11240
rect 12434 11228 12440 11240
rect 12492 11268 12498 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 12492 11240 13645 11268
rect 12492 11228 12498 11240
rect 13188 11212 13216 11240
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 18506 11228 18512 11280
rect 18564 11268 18570 11280
rect 18966 11268 18972 11280
rect 18564 11240 18972 11268
rect 18564 11228 18570 11240
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 20438 11228 20444 11280
rect 20496 11268 20502 11280
rect 20496 11240 22508 11268
rect 20496 11228 20502 11240
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 2777 11203 2835 11209
rect 2777 11200 2789 11203
rect 1995 11172 2789 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 2777 11169 2789 11172
rect 2823 11200 2835 11203
rect 3602 11200 3608 11212
rect 2823 11172 3608 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3602 11160 3608 11172
rect 3660 11160 3666 11212
rect 5994 11200 6000 11212
rect 5907 11172 6000 11200
rect 5994 11160 6000 11172
rect 6052 11200 6058 11212
rect 6546 11200 6552 11212
rect 6052 11172 6552 11200
rect 6052 11160 6058 11172
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 10597 11203 10655 11209
rect 7616 11172 8524 11200
rect 7616 11160 7622 11172
rect 8496 11144 8524 11172
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 10686 11200 10692 11212
rect 10643 11172 10692 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 10962 11209 10968 11212
rect 10956 11200 10968 11209
rect 10875 11172 10968 11200
rect 10956 11163 10968 11172
rect 11020 11200 11026 11212
rect 11020 11172 12848 11200
rect 10962 11160 10968 11163
rect 11020 11160 11026 11172
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 2372 11104 2881 11132
rect 2372 11092 2378 11104
rect 2869 11101 2881 11104
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 2961 11095 3019 11101
rect 2222 11064 2228 11076
rect 2183 11036 2228 11064
rect 2222 11024 2228 11036
rect 2280 11064 2286 11076
rect 2590 11064 2596 11076
rect 2280 11036 2596 11064
rect 2280 11024 2286 11036
rect 2590 11024 2596 11036
rect 2648 11024 2654 11076
rect 2976 11064 3004 11095
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6178 11132 6184 11144
rect 6135 11104 6184 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11132 6331 11135
rect 6454 11132 6460 11144
rect 6319 11104 6460 11132
rect 6319 11101 6331 11104
rect 6273 11095 6331 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 8386 11132 8392 11144
rect 8347 11104 8392 11132
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 9677 11135 9735 11141
rect 8536 11104 8629 11132
rect 8536 11092 8542 11104
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 9723 11104 10732 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 2884 11036 3004 11064
rect 2406 10956 2412 11008
rect 2464 10996 2470 11008
rect 2884 10996 2912 11036
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 3421 11067 3479 11073
rect 3421 11064 3433 11067
rect 3200 11036 3433 11064
rect 3200 11024 3206 11036
rect 3421 11033 3433 11036
rect 3467 11033 3479 11067
rect 3421 11027 3479 11033
rect 3881 11067 3939 11073
rect 3881 11033 3893 11067
rect 3927 11064 3939 11067
rect 3970 11064 3976 11076
rect 3927 11036 3976 11064
rect 3927 11033 3939 11036
rect 3881 11027 3939 11033
rect 3970 11024 3976 11036
rect 4028 11064 4034 11076
rect 4632 11064 4660 11092
rect 4028 11036 4660 11064
rect 4028 11024 4034 11036
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5629 11067 5687 11073
rect 5629 11064 5641 11067
rect 5592 11036 5641 11064
rect 5592 11024 5598 11036
rect 5629 11033 5641 11036
rect 5675 11064 5687 11067
rect 6641 11067 6699 11073
rect 6641 11064 6653 11067
rect 5675 11036 6653 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 6641 11033 6653 11036
rect 6687 11033 6699 11067
rect 10134 11064 10140 11076
rect 10095 11036 10140 11064
rect 6641 11027 6699 11033
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 5074 10996 5080 11008
rect 2464 10968 2912 10996
rect 5035 10968 5080 10996
rect 2464 10956 2470 10968
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5445 10999 5503 11005
rect 5445 10965 5457 10999
rect 5491 10996 5503 10999
rect 5994 10996 6000 11008
rect 5491 10968 6000 10996
rect 5491 10965 5503 10968
rect 5445 10959 5503 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 10704 10996 10732 11104
rect 11330 10996 11336 11008
rect 10704 10968 11336 10996
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 12710 10996 12716 11008
rect 12671 10968 12716 10996
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 12820 10996 12848 11172
rect 13170 11160 13176 11212
rect 13228 11160 13234 11212
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 13722 11200 13728 11212
rect 13587 11172 13728 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 15556 11203 15614 11209
rect 15556 11200 15568 11203
rect 15068 11172 15568 11200
rect 15068 11160 15074 11172
rect 15556 11169 15568 11172
rect 15602 11200 15614 11203
rect 16114 11200 16120 11212
rect 15602 11172 16120 11200
rect 15602 11169 15614 11172
rect 15556 11163 15614 11169
rect 16114 11160 16120 11172
rect 16172 11160 16178 11212
rect 19610 11200 19616 11212
rect 19571 11172 19616 11200
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 19702 11160 19708 11212
rect 19760 11200 19766 11212
rect 19978 11200 19984 11212
rect 19760 11172 19984 11200
rect 19760 11160 19766 11172
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 21157 11203 21215 11209
rect 21157 11200 21169 11203
rect 20088 11172 21169 11200
rect 20088 11144 20116 11172
rect 21157 11169 21169 11172
rect 21203 11169 21215 11203
rect 21157 11163 21215 11169
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11132 13875 11135
rect 13906 11132 13912 11144
rect 13863 11104 13912 11132
rect 13863 11101 13875 11104
rect 13817 11095 13875 11101
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 14274 11132 14280 11144
rect 14187 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11132 14338 11144
rect 15286 11132 15292 11144
rect 14332 11104 15292 11132
rect 14332 11092 14338 11104
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11132 18199 11135
rect 18506 11132 18512 11144
rect 18187 11104 18512 11132
rect 18187 11101 18199 11104
rect 18141 11095 18199 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11132 19947 11135
rect 20070 11132 20076 11144
rect 19935 11104 20076 11132
rect 19935 11101 19947 11104
rect 19889 11095 19947 11101
rect 20070 11092 20076 11104
rect 20128 11092 20134 11144
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 20901 11135 20959 11141
rect 20901 11132 20913 11135
rect 20772 11104 20913 11132
rect 20772 11092 20778 11104
rect 20901 11101 20913 11104
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 20349 11067 20407 11073
rect 20349 11033 20361 11067
rect 20395 11064 20407 11067
rect 20395 11036 20760 11064
rect 20395 11033 20407 11036
rect 20349 11027 20407 11033
rect 20732 11008 20760 11036
rect 21910 11024 21916 11076
rect 21968 11064 21974 11076
rect 22281 11067 22339 11073
rect 22281 11064 22293 11067
rect 21968 11036 22293 11064
rect 21968 11024 21974 11036
rect 22281 11033 22293 11036
rect 22327 11033 22339 11067
rect 22480 11064 22508 11240
rect 22738 11228 22744 11280
rect 22796 11228 22802 11280
rect 22848 11268 22876 11299
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25130 11336 25136 11348
rect 25091 11308 25136 11336
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 23474 11268 23480 11280
rect 22848 11240 23480 11268
rect 23474 11228 23480 11240
rect 23532 11228 23538 11280
rect 22554 11160 22560 11212
rect 22612 11200 22618 11212
rect 22756 11200 22784 11228
rect 22612 11172 22784 11200
rect 22612 11160 22618 11172
rect 23566 11160 23572 11212
rect 23624 11200 23630 11212
rect 23753 11203 23811 11209
rect 23753 11200 23765 11203
rect 23624 11172 23765 11200
rect 23624 11160 23630 11172
rect 23753 11169 23765 11172
rect 23799 11200 23811 11203
rect 23842 11200 23848 11212
rect 23799 11172 23848 11200
rect 23799 11169 23811 11172
rect 23753 11163 23811 11169
rect 23842 11160 23848 11172
rect 23900 11160 23906 11212
rect 24578 11160 24584 11212
rect 24636 11200 24642 11212
rect 24946 11200 24952 11212
rect 24636 11172 24952 11200
rect 24636 11160 24642 11172
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 22738 11092 22744 11144
rect 22796 11132 22802 11144
rect 23934 11132 23940 11144
rect 22796 11104 23940 11132
rect 22796 11092 22802 11104
rect 23934 11092 23940 11104
rect 23992 11092 23998 11144
rect 23109 11067 23167 11073
rect 23109 11064 23121 11067
rect 22480 11036 23121 11064
rect 22281 11027 22339 11033
rect 23109 11033 23121 11036
rect 23155 11064 23167 11067
rect 23201 11067 23259 11073
rect 23201 11064 23213 11067
rect 23155 11036 23213 11064
rect 23155 11033 23167 11036
rect 23109 11027 23167 11033
rect 23201 11033 23213 11036
rect 23247 11033 23259 11067
rect 23201 11027 23259 11033
rect 24210 11024 24216 11076
rect 24268 11064 24274 11076
rect 24581 11067 24639 11073
rect 24581 11064 24593 11067
rect 24268 11036 24593 11064
rect 24268 11024 24274 11036
rect 24581 11033 24593 11036
rect 24627 11033 24639 11067
rect 24581 11027 24639 11033
rect 16850 10996 16856 11008
rect 12820 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 18049 10999 18107 11005
rect 18049 10965 18061 10999
rect 18095 10996 18107 10999
rect 18598 10996 18604 11008
rect 18095 10968 18604 10996
rect 18095 10965 18107 10968
rect 18049 10959 18107 10965
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 19153 10999 19211 11005
rect 19153 10965 19165 10999
rect 19199 10996 19211 10999
rect 19518 10996 19524 11008
rect 19199 10968 19524 10996
rect 19199 10965 19211 10968
rect 19153 10959 19211 10965
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 20714 10956 20720 11008
rect 20772 10956 20778 11008
rect 23382 10996 23388 11008
rect 23343 10968 23388 10996
rect 23382 10956 23388 10968
rect 23440 10956 23446 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 2130 10792 2136 10804
rect 1627 10764 2136 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4614 10792 4620 10804
rect 4019 10764 4620 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4890 10752 4896 10804
rect 4948 10792 4954 10804
rect 5077 10795 5135 10801
rect 5077 10792 5089 10795
rect 4948 10764 5089 10792
rect 4948 10752 4954 10764
rect 5077 10761 5089 10764
rect 5123 10761 5135 10795
rect 5077 10755 5135 10761
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 7156 10764 7573 10792
rect 7156 10752 7162 10764
rect 7561 10761 7573 10764
rect 7607 10792 7619 10795
rect 8018 10792 8024 10804
rect 7607 10764 8024 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 11425 10795 11483 10801
rect 11425 10792 11437 10795
rect 10744 10764 11437 10792
rect 10744 10752 10750 10764
rect 11425 10761 11437 10764
rect 11471 10792 11483 10795
rect 12526 10792 12532 10804
rect 11471 10764 12532 10792
rect 11471 10761 11483 10764
rect 11425 10755 11483 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 13228 10764 13461 10792
rect 13228 10752 13234 10764
rect 13449 10761 13461 10764
rect 13495 10761 13507 10795
rect 13449 10755 13507 10761
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 13964 10764 14197 10792
rect 13964 10752 13970 10764
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 14185 10755 14243 10761
rect 15013 10795 15071 10801
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15286 10792 15292 10804
rect 15059 10764 15292 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15286 10752 15292 10764
rect 15344 10792 15350 10804
rect 15381 10795 15439 10801
rect 15381 10792 15393 10795
rect 15344 10764 15393 10792
rect 15344 10752 15350 10764
rect 15381 10761 15393 10764
rect 15427 10792 15439 10795
rect 16758 10792 16764 10804
rect 15427 10764 16764 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 7190 10724 7196 10736
rect 7151 10696 7196 10724
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 10321 10727 10379 10733
rect 10321 10724 10333 10727
rect 9548 10696 10333 10724
rect 9548 10684 9554 10696
rect 10321 10693 10333 10696
rect 10367 10724 10379 10727
rect 11606 10724 11612 10736
rect 10367 10696 11612 10724
rect 10367 10693 10379 10696
rect 10321 10687 10379 10693
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 12437 10727 12495 10733
rect 12437 10693 12449 10727
rect 12483 10724 12495 10727
rect 12894 10724 12900 10736
rect 12483 10696 12900 10724
rect 12483 10693 12495 10696
rect 12437 10687 12495 10693
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 5074 10616 5080 10668
rect 5132 10656 5138 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5132 10628 5549 10656
rect 5132 10616 5138 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 5994 10656 6000 10668
rect 5767 10628 6000 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 5994 10616 6000 10628
rect 6052 10656 6058 10668
rect 6454 10656 6460 10668
rect 6052 10628 6460 10656
rect 6052 10616 6058 10628
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 7650 10656 7656 10668
rect 7611 10628 7656 10656
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10275 10628 10885 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10873 10625 10885 10628
rect 10919 10656 10931 10659
rect 11422 10656 11428 10668
rect 10919 10628 11428 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 12250 10656 12256 10668
rect 12163 10628 12256 10656
rect 12250 10616 12256 10628
rect 12308 10656 12314 10668
rect 15488 10665 15516 10764
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 16850 10752 16856 10804
rect 16908 10792 16914 10804
rect 16908 10764 16953 10792
rect 16908 10752 16914 10764
rect 19242 10752 19248 10804
rect 19300 10792 19306 10804
rect 19610 10792 19616 10804
rect 19300 10764 19616 10792
rect 19300 10752 19306 10764
rect 19610 10752 19616 10764
rect 19668 10792 19674 10804
rect 20073 10795 20131 10801
rect 20073 10792 20085 10795
rect 19668 10764 20085 10792
rect 19668 10752 19674 10764
rect 20073 10761 20085 10764
rect 20119 10761 20131 10795
rect 20073 10755 20131 10761
rect 20625 10795 20683 10801
rect 20625 10761 20637 10795
rect 20671 10792 20683 10795
rect 21450 10792 21456 10804
rect 20671 10764 21456 10792
rect 20671 10761 20683 10764
rect 20625 10755 20683 10761
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 22646 10792 22652 10804
rect 22607 10764 22652 10792
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 24946 10792 24952 10804
rect 24907 10764 24952 10792
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 25409 10795 25467 10801
rect 25409 10761 25421 10795
rect 25455 10792 25467 10795
rect 25498 10792 25504 10804
rect 25455 10764 25504 10792
rect 25455 10761 25467 10764
rect 25409 10755 25467 10761
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 20533 10727 20591 10733
rect 20533 10693 20545 10727
rect 20579 10724 20591 10727
rect 21910 10724 21916 10736
rect 20579 10696 21916 10724
rect 20579 10693 20591 10696
rect 20533 10687 20591 10693
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12308 10628 13001 10656
rect 12308 10616 12314 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 21082 10656 21088 10668
rect 21043 10628 21088 10656
rect 15473 10619 15531 10625
rect 21082 10616 21088 10628
rect 21140 10616 21146 10668
rect 21192 10665 21220 10696
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 23477 10727 23535 10733
rect 23477 10693 23489 10727
rect 23523 10724 23535 10727
rect 23658 10724 23664 10736
rect 23523 10696 23664 10724
rect 23523 10693 23535 10696
rect 23477 10687 23535 10693
rect 23658 10684 23664 10696
rect 23716 10724 23722 10736
rect 23716 10696 24164 10724
rect 23716 10684 23722 10696
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10625 21235 10659
rect 21177 10619 21235 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 2501 10591 2559 10597
rect 1443 10560 1716 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1688 10464 1716 10560
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2593 10591 2651 10597
rect 2593 10588 2605 10591
rect 2547 10560 2605 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2593 10557 2605 10560
rect 2639 10588 2651 10591
rect 4430 10588 4436 10600
rect 2639 10560 4436 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 7920 10591 7978 10597
rect 7920 10557 7932 10591
rect 7966 10588 7978 10591
rect 8202 10588 8208 10600
rect 7966 10560 8208 10588
rect 7966 10557 7978 10560
rect 7920 10551 7978 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 12526 10588 12532 10600
rect 11808 10560 12532 10588
rect 2860 10523 2918 10529
rect 2860 10489 2872 10523
rect 2906 10520 2918 10523
rect 3418 10520 3424 10532
rect 2906 10492 3424 10520
rect 2906 10489 2918 10492
rect 2860 10483 2918 10489
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 4985 10523 5043 10529
rect 4985 10489 4997 10523
rect 5031 10520 5043 10523
rect 5350 10520 5356 10532
rect 5031 10492 5356 10520
rect 5031 10489 5043 10492
rect 4985 10483 5043 10489
rect 5350 10480 5356 10492
rect 5408 10520 5414 10532
rect 5445 10523 5503 10529
rect 5445 10520 5457 10523
rect 5408 10492 5457 10520
rect 5408 10480 5414 10492
rect 5445 10489 5457 10492
rect 5491 10489 5503 10523
rect 6178 10520 6184 10532
rect 6091 10492 6184 10520
rect 5445 10483 5503 10489
rect 6178 10480 6184 10492
rect 6236 10520 6242 10532
rect 8110 10520 8116 10532
rect 6236 10492 8116 10520
rect 6236 10480 6242 10492
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 9784 10492 10793 10520
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 1949 10455 2007 10461
rect 1949 10452 1961 10455
rect 1728 10424 1961 10452
rect 1728 10412 1734 10424
rect 1949 10421 1961 10424
rect 1995 10421 2007 10455
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 1949 10415 2007 10421
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 9030 10452 9036 10464
rect 8991 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9784 10461 9812 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 10781 10483 10839 10489
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 11808 10529 11836 10560
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 15746 10597 15752 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12768 10560 12817 10588
rect 12768 10548 12774 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 15740 10588 15752 10597
rect 15659 10560 15752 10588
rect 12805 10551 12863 10557
rect 15740 10551 15752 10560
rect 15804 10588 15810 10600
rect 16482 10588 16488 10600
rect 15804 10560 16488 10588
rect 15746 10548 15752 10551
rect 15804 10548 15810 10560
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 18138 10588 18144 10600
rect 18099 10560 18144 10588
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 20993 10591 21051 10597
rect 20993 10588 21005 10591
rect 20772 10560 21005 10588
rect 20772 10548 20778 10560
rect 20993 10557 21005 10560
rect 21039 10557 21051 10591
rect 20993 10551 21051 10557
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22465 10591 22523 10597
rect 22465 10588 22477 10591
rect 22244 10560 22477 10588
rect 22244 10548 22250 10560
rect 22465 10557 22477 10560
rect 22511 10588 22523 10591
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22511 10560 23029 10588
rect 22511 10557 22523 10560
rect 22465 10551 22523 10557
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 23017 10551 23075 10557
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 24136 10597 24164 10696
rect 24305 10659 24363 10665
rect 24305 10625 24317 10659
rect 24351 10656 24363 10659
rect 25038 10656 25044 10668
rect 24351 10628 25044 10656
rect 24351 10625 24363 10628
rect 24305 10619 24363 10625
rect 25038 10616 25044 10628
rect 25096 10616 25102 10668
rect 24029 10591 24087 10597
rect 24029 10588 24041 10591
rect 23532 10560 24041 10588
rect 23532 10548 23538 10560
rect 24029 10557 24041 10560
rect 24075 10557 24087 10591
rect 24029 10551 24087 10557
rect 24121 10591 24179 10597
rect 24121 10557 24133 10591
rect 24167 10588 24179 10591
rect 24670 10588 24676 10600
rect 24167 10560 24676 10588
rect 24167 10557 24179 10560
rect 24121 10551 24179 10557
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 25222 10588 25228 10600
rect 25183 10560 25228 10588
rect 25222 10548 25228 10560
rect 25280 10588 25286 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25280 10560 25789 10588
rect 25280 10548 25286 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 11793 10523 11851 10529
rect 11793 10520 11805 10523
rect 11204 10492 11805 10520
rect 11204 10480 11210 10492
rect 11793 10489 11805 10492
rect 11839 10489 11851 10523
rect 18386 10523 18444 10529
rect 18386 10520 18398 10523
rect 11793 10483 11851 10489
rect 17420 10492 18398 10520
rect 17420 10464 17448 10492
rect 18386 10489 18398 10492
rect 18432 10489 18444 10523
rect 18386 10483 18444 10489
rect 20622 10480 20628 10532
rect 20680 10520 20686 10532
rect 21637 10523 21695 10529
rect 21637 10520 21649 10523
rect 20680 10492 21649 10520
rect 20680 10480 20686 10492
rect 21637 10489 21649 10492
rect 21683 10520 21695 10523
rect 21818 10520 21824 10532
rect 21683 10492 21824 10520
rect 21683 10489 21695 10492
rect 21637 10483 21695 10489
rect 21818 10480 21824 10492
rect 21876 10480 21882 10532
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 9732 10424 9781 10452
rect 9732 10412 9738 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 10686 10452 10692 10464
rect 10647 10424 10692 10452
rect 9769 10415 9827 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12584 10424 12909 10452
rect 12584 10412 12590 10424
rect 12897 10421 12909 10424
rect 12943 10421 12955 10455
rect 12897 10415 12955 10421
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 13780 10424 13921 10452
rect 13780 10412 13786 10424
rect 13909 10421 13921 10424
rect 13955 10452 13967 10455
rect 14366 10452 14372 10464
rect 13955 10424 14372 10452
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 17402 10452 17408 10464
rect 14516 10424 14561 10452
rect 17363 10424 17408 10452
rect 14516 10412 14522 10424
rect 17402 10412 17408 10424
rect 17460 10412 17466 10464
rect 17862 10452 17868 10464
rect 17775 10424 17868 10452
rect 17862 10412 17868 10424
rect 17920 10452 17926 10464
rect 18138 10452 18144 10464
rect 17920 10424 18144 10452
rect 17920 10412 17926 10424
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 19518 10452 19524 10464
rect 19479 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 22002 10452 22008 10464
rect 21963 10424 22008 10452
rect 22002 10412 22008 10424
rect 22060 10412 22066 10464
rect 22462 10412 22468 10464
rect 22520 10452 22526 10464
rect 22646 10452 22652 10464
rect 22520 10424 22652 10452
rect 22520 10412 22526 10424
rect 22646 10412 22652 10424
rect 22704 10412 22710 10464
rect 23658 10452 23664 10464
rect 23619 10424 23664 10452
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 1854 10248 1860 10260
rect 1627 10220 1860 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2314 10248 2320 10260
rect 1995 10220 2320 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 2590 10248 2596 10260
rect 2455 10220 2596 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2832 10220 2877 10248
rect 2832 10208 2838 10220
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7432 10220 7573 10248
rect 7432 10208 7438 10220
rect 7561 10217 7573 10220
rect 7607 10248 7619 10251
rect 8294 10248 8300 10260
rect 7607 10220 8300 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8536 10220 8585 10248
rect 8536 10208 8542 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 9490 10248 9496 10260
rect 9451 10220 9496 10248
rect 8573 10211 8631 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10686 10248 10692 10260
rect 10091 10220 10692 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 10962 10248 10968 10260
rect 10923 10220 10968 10248
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11606 10248 11612 10260
rect 11567 10220 11612 10248
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 12710 10248 12716 10260
rect 12671 10220 12716 10248
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13170 10248 13176 10260
rect 13131 10220 13176 10248
rect 13170 10208 13176 10220
rect 13228 10208 13234 10260
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16114 10248 16120 10260
rect 16075 10220 16120 10248
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 17310 10248 17316 10260
rect 17175 10220 17316 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18230 10248 18236 10260
rect 18191 10220 18236 10248
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 19334 10208 19340 10260
rect 19392 10248 19398 10260
rect 20530 10248 20536 10260
rect 19392 10220 20536 10248
rect 19392 10208 19398 10220
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20772 10220 20913 10248
rect 20772 10208 20778 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 21266 10248 21272 10260
rect 21227 10220 21272 10248
rect 20901 10211 20959 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 22097 10251 22155 10257
rect 22097 10217 22109 10251
rect 22143 10248 22155 10251
rect 22278 10248 22284 10260
rect 22143 10220 22284 10248
rect 22143 10217 22155 10220
rect 22097 10211 22155 10217
rect 22278 10208 22284 10220
rect 22336 10248 22342 10260
rect 23382 10248 23388 10260
rect 22336 10220 23388 10248
rect 22336 10208 22342 10220
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 25038 10208 25044 10260
rect 25096 10248 25102 10260
rect 25133 10251 25191 10257
rect 25133 10248 25145 10251
rect 25096 10220 25145 10248
rect 25096 10208 25102 10220
rect 25133 10217 25145 10220
rect 25179 10217 25191 10251
rect 25133 10211 25191 10217
rect 2498 10140 2504 10192
rect 2556 10180 2562 10192
rect 6270 10180 6276 10192
rect 2556 10152 6276 10180
rect 2556 10140 2562 10152
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 12250 10140 12256 10192
rect 12308 10180 12314 10192
rect 13081 10183 13139 10189
rect 13081 10180 13093 10183
rect 12308 10152 13093 10180
rect 12308 10140 12314 10152
rect 13081 10149 13093 10152
rect 13127 10149 13139 10183
rect 13081 10143 13139 10149
rect 13538 10140 13544 10192
rect 13596 10180 13602 10192
rect 17770 10180 17776 10192
rect 13596 10152 17776 10180
rect 13596 10140 13602 10152
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 19978 10180 19984 10192
rect 19352 10152 19984 10180
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10081 1455 10115
rect 1397 10075 1455 10081
rect 1412 10044 1440 10075
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 3878 10112 3884 10124
rect 1636 10084 3884 10112
rect 1636 10072 1642 10084
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4792 10115 4850 10121
rect 4792 10112 4804 10115
rect 4212 10084 4804 10112
rect 4212 10072 4218 10084
rect 4792 10081 4804 10084
rect 4838 10112 4850 10115
rect 6454 10112 6460 10124
rect 4838 10084 6460 10112
rect 4838 10081 4850 10084
rect 4792 10075 4850 10081
rect 6454 10072 6460 10084
rect 6512 10072 6518 10124
rect 7926 10112 7932 10124
rect 7887 10084 7932 10112
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8110 10112 8116 10124
rect 8067 10084 8116 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 11112 10084 11529 10112
rect 11112 10072 11118 10084
rect 11517 10081 11529 10084
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 19352 10121 19380 10152
rect 19978 10140 19984 10152
rect 20036 10140 20042 10192
rect 22738 10180 22744 10192
rect 22699 10152 22744 10180
rect 22738 10140 22744 10152
rect 22796 10140 22802 10192
rect 23109 10183 23167 10189
rect 23109 10149 23121 10183
rect 23155 10180 23167 10183
rect 23566 10180 23572 10192
rect 23155 10152 23572 10180
rect 23155 10149 23167 10152
rect 23109 10143 23167 10149
rect 23566 10140 23572 10152
rect 23624 10140 23630 10192
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 17000 10084 17049 10112
rect 17000 10072 17006 10084
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 19337 10115 19395 10121
rect 19337 10081 19349 10115
rect 19383 10081 19395 10115
rect 19794 10112 19800 10124
rect 19755 10084 19800 10112
rect 19337 10075 19395 10081
rect 19794 10072 19800 10084
rect 19852 10072 19858 10124
rect 21818 10072 21824 10124
rect 21876 10112 21882 10124
rect 23014 10112 23020 10124
rect 21876 10084 23020 10112
rect 21876 10072 21882 10084
rect 23014 10072 23020 10084
rect 23072 10112 23078 10124
rect 23201 10115 23259 10121
rect 23201 10112 23213 10115
rect 23072 10084 23213 10112
rect 23072 10072 23078 10084
rect 23201 10081 23213 10084
rect 23247 10081 23259 10115
rect 23468 10115 23526 10121
rect 23468 10112 23480 10115
rect 23201 10075 23259 10081
rect 23308 10084 23480 10112
rect 2590 10044 2596 10056
rect 1412 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 3016 10016 3065 10044
rect 3016 10004 3022 10016
rect 3053 10013 3065 10016
rect 3099 10044 3111 10047
rect 3602 10044 3608 10056
rect 3099 10016 3608 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 4430 10004 4436 10056
rect 4488 10044 4494 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4488 10016 4537 10044
rect 4488 10004 4494 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 8202 10044 8208 10056
rect 8163 10016 8208 10044
rect 4525 10007 4583 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10013 11759 10047
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 11701 10007 11759 10013
rect 3418 9936 3424 9988
rect 3476 9976 3482 9988
rect 3513 9979 3571 9985
rect 3513 9976 3525 9979
rect 3476 9948 3525 9976
rect 3476 9936 3482 9948
rect 3513 9945 3525 9948
rect 3559 9976 3571 9979
rect 7098 9976 7104 9988
rect 3559 9948 4476 9976
rect 7011 9948 7104 9976
rect 3559 9945 3571 9948
rect 3513 9939 3571 9945
rect 2314 9908 2320 9920
rect 2275 9880 2320 9908
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4448 9917 4476 9948
rect 7098 9936 7104 9948
rect 7156 9976 7162 9988
rect 7469 9979 7527 9985
rect 7469 9976 7481 9979
rect 7156 9948 7481 9976
rect 7156 9936 7162 9948
rect 7469 9945 7481 9948
rect 7515 9976 7527 9979
rect 8220 9976 8248 10004
rect 8938 9976 8944 9988
rect 7515 9948 8248 9976
rect 8899 9948 8944 9976
rect 7515 9945 7527 9948
rect 7469 9939 7527 9945
rect 8938 9936 8944 9948
rect 8996 9936 9002 9988
rect 10321 9979 10379 9985
rect 10321 9945 10333 9979
rect 10367 9976 10379 9979
rect 10962 9976 10968 9988
rect 10367 9948 10968 9976
rect 10367 9945 10379 9948
rect 10321 9939 10379 9945
rect 10962 9936 10968 9948
rect 11020 9936 11026 9988
rect 11146 9976 11152 9988
rect 11107 9948 11152 9976
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11514 9936 11520 9988
rect 11572 9976 11578 9988
rect 11716 9976 11744 10007
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 14884 10016 15301 10044
rect 14884 10004 14890 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 17402 10044 17408 10056
rect 17359 10016 17408 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10044 17831 10047
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 17819 10016 18705 10044
rect 17819 10013 17831 10016
rect 17773 10007 17831 10013
rect 18693 10013 18705 10016
rect 18739 10013 18751 10047
rect 18693 10007 18751 10013
rect 18877 10047 18935 10053
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 19518 10044 19524 10056
rect 18923 10016 19524 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 11572 9948 11744 9976
rect 16669 9979 16727 9985
rect 11572 9936 11578 9948
rect 16669 9945 16681 9979
rect 16715 9976 16727 9979
rect 17788 9976 17816 10007
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 21082 10004 21088 10056
rect 21140 10044 21146 10056
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 21140 10016 21373 10044
rect 21140 10004 21146 10016
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 21361 10007 21419 10013
rect 21453 10047 21511 10053
rect 21453 10013 21465 10047
rect 21499 10044 21511 10047
rect 22002 10044 22008 10056
rect 21499 10016 22008 10044
rect 21499 10013 21511 10016
rect 21453 10007 21511 10013
rect 19978 9976 19984 9988
rect 16715 9948 17816 9976
rect 19939 9948 19984 9976
rect 16715 9945 16727 9948
rect 16669 9939 16727 9945
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 21468 9976 21496 10007
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 23308 10044 23336 10084
rect 23468 10081 23480 10084
rect 23514 10112 23526 10115
rect 25056 10112 25084 10208
rect 23514 10084 25084 10112
rect 23514 10081 23526 10084
rect 23468 10075 23526 10081
rect 23164 10016 23336 10044
rect 23164 10004 23170 10016
rect 20364 9948 21496 9976
rect 20364 9920 20392 9948
rect 4433 9911 4491 9917
rect 4433 9877 4445 9911
rect 4479 9908 4491 9911
rect 5166 9908 5172 9920
rect 4479 9880 5172 9908
rect 4479 9877 4491 9880
rect 4433 9871 4491 9877
rect 5166 9868 5172 9880
rect 5224 9908 5230 9920
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 5224 9880 5917 9908
rect 5224 9868 5230 9880
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 6454 9908 6460 9920
rect 6415 9880 6460 9908
rect 5905 9871 5963 9877
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 10594 9908 10600 9920
rect 10555 9880 10600 9908
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12802 9908 12808 9920
rect 12575 9880 12808 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 13817 9911 13875 9917
rect 13817 9908 13829 9911
rect 13780 9880 13829 9908
rect 13780 9868 13786 9880
rect 13817 9877 13829 9880
rect 13863 9877 13875 9911
rect 14090 9908 14096 9920
rect 14051 9880 14096 9908
rect 13817 9871 13875 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14550 9908 14556 9920
rect 14511 9880 14556 9908
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 16574 9908 16580 9920
rect 16535 9880 16580 9908
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 20070 9908 20076 9920
rect 19751 9880 20076 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 20070 9868 20076 9880
rect 20128 9908 20134 9920
rect 20346 9908 20352 9920
rect 20128 9880 20352 9908
rect 20128 9868 20134 9880
rect 20346 9868 20352 9880
rect 20404 9868 20410 9920
rect 24581 9911 24639 9917
rect 24581 9877 24593 9911
rect 24627 9908 24639 9911
rect 24670 9908 24676 9920
rect 24627 9880 24676 9908
rect 24627 9877 24639 9880
rect 24581 9871 24639 9877
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1578 9704 1584 9716
rect 1539 9676 1584 9704
rect 1578 9664 1584 9676
rect 1636 9664 1642 9716
rect 2314 9664 2320 9716
rect 2372 9704 2378 9716
rect 5994 9704 6000 9716
rect 2372 9676 6000 9704
rect 2372 9664 2378 9676
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 9858 9704 9864 9716
rect 9732 9676 9864 9704
rect 9732 9664 9738 9676
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 10413 9707 10471 9713
rect 10413 9673 10425 9707
rect 10459 9704 10471 9707
rect 10686 9704 10692 9716
rect 10459 9676 10692 9704
rect 10459 9673 10471 9676
rect 10413 9667 10471 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 11112 9676 12388 9704
rect 11112 9664 11118 9676
rect 2774 9636 2780 9648
rect 2735 9608 2780 9636
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 3881 9639 3939 9645
rect 3881 9605 3893 9639
rect 3927 9636 3939 9639
rect 4154 9636 4160 9648
rect 3927 9608 4160 9636
rect 3927 9605 3939 9608
rect 3881 9599 3939 9605
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 4338 9636 4344 9648
rect 4299 9608 4344 9636
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 4908 9608 6561 9636
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 3418 9568 3424 9580
rect 2731 9540 3424 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 4908 9568 4936 9608
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 9306 9636 9312 9648
rect 9267 9608 9312 9636
rect 6549 9599 6607 9605
rect 4080 9540 4936 9568
rect 4985 9571 5043 9577
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 3234 9500 3240 9512
rect 1443 9472 2084 9500
rect 3195 9472 3240 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 2056 9376 2084 9472
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 2038 9364 2044 9376
rect 1999 9336 2044 9364
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3234 9364 3240 9376
rect 3191 9336 3240 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 4080 9364 4108 9540
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5166 9568 5172 9580
rect 5031 9540 5172 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 6564 9568 6592 9599
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 11330 9596 11336 9648
rect 11388 9636 11394 9648
rect 11793 9639 11851 9645
rect 11793 9636 11805 9639
rect 11388 9608 11805 9636
rect 11388 9596 11394 9608
rect 11793 9605 11805 9608
rect 11839 9636 11851 9639
rect 12250 9636 12256 9648
rect 11839 9608 12256 9636
rect 11839 9605 11851 9608
rect 11793 9599 11851 9605
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 6564 9540 8064 9568
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9500 4859 9503
rect 5442 9500 5448 9512
rect 4847 9472 5448 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7929 9503 7987 9509
rect 7929 9500 7941 9503
rect 7708 9472 7941 9500
rect 7708 9460 7714 9472
rect 7929 9469 7941 9472
rect 7975 9469 7987 9503
rect 8036 9500 8064 9540
rect 10686 9528 10692 9580
rect 10744 9568 10750 9580
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10744 9540 10977 9568
rect 10744 9528 10750 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11480 9540 11621 9568
rect 11480 9528 11486 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 12360 9568 12388 9676
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 13412 9676 13768 9704
rect 13412 9664 13418 9676
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9605 12495 9639
rect 12437 9599 12495 9605
rect 12452 9568 12480 9599
rect 13170 9596 13176 9648
rect 13228 9636 13234 9648
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 13228 9608 13461 9636
rect 13228 9596 13234 9608
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 13740 9636 13768 9676
rect 17310 9664 17316 9716
rect 17368 9704 17374 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 17368 9676 17417 9704
rect 17368 9664 17374 9676
rect 17405 9673 17417 9676
rect 17451 9673 17463 9707
rect 17405 9667 17463 9673
rect 17865 9707 17923 9713
rect 17865 9673 17877 9707
rect 17911 9704 17923 9707
rect 18230 9704 18236 9716
rect 17911 9676 18236 9704
rect 17911 9673 17923 9676
rect 17865 9667 17923 9673
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13740 9608 13829 9636
rect 13449 9599 13507 9605
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 13817 9599 13875 9605
rect 14461 9639 14519 9645
rect 14461 9605 14473 9639
rect 14507 9636 14519 9639
rect 14507 9608 15148 9636
rect 14507 9605 14519 9608
rect 14461 9599 14519 9605
rect 12360 9540 12480 9568
rect 13081 9571 13139 9577
rect 11609 9531 11667 9537
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13722 9568 13728 9580
rect 13127 9540 13728 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 8185 9503 8243 9509
rect 8185 9500 8197 9503
rect 8036 9472 8197 9500
rect 7929 9463 7987 9469
rect 8185 9469 8197 9472
rect 8231 9500 8243 9503
rect 9030 9500 9036 9512
rect 8231 9472 9036 9500
rect 8231 9469 8243 9472
rect 8185 9463 8243 9469
rect 4249 9435 4307 9441
rect 4249 9401 4261 9435
rect 4295 9432 4307 9435
rect 4709 9435 4767 9441
rect 4709 9432 4721 9435
rect 4295 9404 4721 9432
rect 4295 9401 4307 9404
rect 4249 9395 4307 9401
rect 4709 9401 4721 9404
rect 4755 9432 4767 9435
rect 6825 9435 6883 9441
rect 6825 9432 6837 9435
rect 4755 9404 6837 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 6825 9401 6837 9404
rect 6871 9401 6883 9435
rect 7944 9432 7972 9463
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 9916 9472 10333 9500
rect 9916 9460 9922 9472
rect 10321 9469 10333 9472
rect 10367 9500 10379 9503
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 10367 9472 10793 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 10781 9469 10793 9472
rect 10827 9500 10839 9503
rect 10870 9500 10876 9512
rect 10827 9472 10876 9500
rect 10827 9469 10839 9472
rect 10781 9463 10839 9469
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 12158 9500 12164 9512
rect 12119 9472 12164 9500
rect 12158 9460 12164 9472
rect 12216 9500 12222 9512
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12216 9472 12909 9500
rect 12216 9460 12222 9472
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 8570 9432 8576 9444
rect 7944 9404 8576 9432
rect 6825 9395 6883 9401
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 11330 9392 11336 9444
rect 11388 9432 11394 9444
rect 12802 9432 12808 9444
rect 11388 9404 12808 9432
rect 11388 9392 11394 9404
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 3568 9336 4108 9364
rect 3568 9324 3574 9336
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 4212 9336 5365 9364
rect 4212 9324 4218 9336
rect 5353 9333 5365 9336
rect 5399 9333 5411 9367
rect 5353 9327 5411 9333
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 5994 9364 6000 9376
rect 5859 9336 6000 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6362 9364 6368 9376
rect 6227 9336 6368 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 7064 9336 7573 9364
rect 7064 9324 7070 9336
rect 7561 9333 7573 9336
rect 7607 9364 7619 9367
rect 7926 9364 7932 9376
rect 7607 9336 7932 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10778 9364 10784 9376
rect 9999 9336 10784 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10778 9324 10784 9336
rect 10836 9364 10842 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10836 9336 10885 9364
rect 10836 9324 10842 9336
rect 10873 9333 10885 9336
rect 10919 9333 10931 9367
rect 11514 9364 11520 9376
rect 11475 9336 11520 9364
rect 10873 9327 10931 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11609 9367 11667 9373
rect 11609 9333 11621 9367
rect 11655 9364 11667 9367
rect 13096 9364 13124 9531
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 15010 9568 15016 9580
rect 14608 9540 15016 9568
rect 14608 9528 14614 9540
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 14826 9500 14832 9512
rect 14787 9472 14832 9500
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 15120 9500 15148 9608
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 16025 9639 16083 9645
rect 16025 9636 16037 9639
rect 15712 9608 16037 9636
rect 15712 9596 15718 9608
rect 16025 9605 16037 9608
rect 16071 9605 16083 9639
rect 16025 9599 16083 9605
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16577 9571 16635 9577
rect 16577 9568 16589 9571
rect 16172 9540 16589 9568
rect 16172 9528 16178 9540
rect 16577 9537 16589 9540
rect 16623 9537 16635 9571
rect 16577 9531 16635 9537
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 15120 9472 16405 9500
rect 16393 9469 16405 9472
rect 16439 9500 16451 9503
rect 16482 9500 16488 9512
rect 16439 9472 16488 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18064 9509 18092 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 19981 9707 20039 9713
rect 19981 9704 19993 9707
rect 19576 9676 19993 9704
rect 19576 9664 19582 9676
rect 19981 9673 19993 9676
rect 20027 9673 20039 9707
rect 20346 9704 20352 9716
rect 20307 9676 20352 9704
rect 19981 9667 20039 9673
rect 20346 9664 20352 9676
rect 20404 9664 20410 9716
rect 21082 9704 21088 9716
rect 21043 9676 21088 9704
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 21266 9664 21272 9716
rect 21324 9704 21330 9716
rect 21453 9707 21511 9713
rect 21453 9704 21465 9707
rect 21324 9676 21465 9704
rect 21324 9664 21330 9676
rect 21453 9673 21465 9676
rect 21499 9673 21511 9707
rect 21453 9667 21511 9673
rect 23014 9664 23020 9716
rect 23072 9704 23078 9716
rect 23293 9707 23351 9713
rect 23293 9704 23305 9707
rect 23072 9676 23305 9704
rect 23072 9664 23078 9676
rect 23293 9673 23305 9676
rect 23339 9673 23351 9707
rect 23293 9667 23351 9673
rect 23198 9596 23204 9648
rect 23256 9636 23262 9648
rect 23661 9639 23719 9645
rect 23661 9636 23673 9639
rect 23256 9608 23673 9636
rect 23256 9596 23262 9608
rect 23661 9605 23673 9608
rect 23707 9605 23719 9639
rect 25406 9636 25412 9648
rect 25367 9608 25412 9636
rect 23661 9599 23719 9605
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 22278 9528 22284 9580
rect 22336 9568 22342 9580
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 22336 9540 22477 9568
rect 22336 9528 22342 9540
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9568 22707 9571
rect 23106 9568 23112 9580
rect 22695 9540 23112 9568
rect 22695 9537 22707 9540
rect 22649 9531 22707 9537
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9568 24363 9571
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 24351 9540 24501 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 24489 9537 24501 9540
rect 24535 9568 24547 9571
rect 24670 9568 24676 9580
rect 24535 9540 24676 9568
rect 24535 9537 24547 9540
rect 24489 9531 24547 9537
rect 24670 9528 24676 9540
rect 24728 9528 24734 9580
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 18012 9472 18061 9500
rect 18012 9460 18018 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 18305 9503 18363 9509
rect 18305 9500 18317 9503
rect 18196 9472 18317 9500
rect 18196 9460 18202 9472
rect 18305 9469 18317 9472
rect 18351 9469 18363 9503
rect 20530 9500 20536 9512
rect 20491 9472 20536 9500
rect 18305 9463 18363 9469
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 21913 9503 21971 9509
rect 21913 9500 21925 9503
rect 20772 9472 21925 9500
rect 20772 9460 20778 9472
rect 21913 9469 21925 9472
rect 21959 9500 21971 9503
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 21959 9472 22385 9500
rect 21959 9469 21971 9472
rect 21913 9463 21971 9469
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 23658 9460 23664 9512
rect 23716 9500 23722 9512
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 23716 9472 24041 9500
rect 23716 9460 23722 9472
rect 24029 9469 24041 9472
rect 24075 9469 24087 9503
rect 25222 9500 25228 9512
rect 25183 9472 25228 9500
rect 24029 9463 24087 9469
rect 25222 9460 25228 9472
rect 25280 9500 25286 9512
rect 25777 9503 25835 9509
rect 25777 9500 25789 9503
rect 25280 9472 25789 9500
rect 25280 9460 25286 9472
rect 25777 9469 25789 9472
rect 25823 9469 25835 9503
rect 25777 9463 25835 9469
rect 14921 9435 14979 9441
rect 14921 9432 14933 9435
rect 14292 9404 14933 9432
rect 14292 9376 14320 9404
rect 14921 9401 14933 9404
rect 14967 9401 14979 9435
rect 14921 9395 14979 9401
rect 15565 9435 15623 9441
rect 15565 9401 15577 9435
rect 15611 9432 15623 9435
rect 16298 9432 16304 9444
rect 15611 9404 16304 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 16298 9392 16304 9404
rect 16356 9432 16362 9444
rect 24121 9435 24179 9441
rect 24121 9432 24133 9435
rect 16356 9404 16528 9432
rect 16356 9392 16362 9404
rect 14274 9364 14280 9376
rect 11655 9336 13124 9364
rect 14235 9336 14280 9364
rect 11655 9333 11667 9336
rect 11609 9327 11667 9333
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 15933 9367 15991 9373
rect 15933 9333 15945 9367
rect 15979 9364 15991 9367
rect 16114 9364 16120 9376
rect 15979 9336 16120 9364
rect 15979 9333 15991 9336
rect 15933 9327 15991 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16500 9373 16528 9404
rect 22020 9404 24133 9432
rect 16485 9367 16543 9373
rect 16485 9333 16497 9367
rect 16531 9333 16543 9367
rect 16485 9327 16543 9333
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17037 9367 17095 9373
rect 17037 9364 17049 9367
rect 17000 9336 17049 9364
rect 17000 9324 17006 9336
rect 17037 9333 17049 9336
rect 17083 9333 17095 9367
rect 17037 9327 17095 9333
rect 19242 9324 19248 9376
rect 19300 9364 19306 9376
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 19300 9336 19441 9364
rect 19300 9324 19306 9336
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19429 9327 19487 9333
rect 20717 9367 20775 9373
rect 20717 9333 20729 9367
rect 20763 9364 20775 9367
rect 20990 9364 20996 9376
rect 20763 9336 20996 9364
rect 20763 9333 20775 9336
rect 20717 9327 20775 9333
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 22020 9373 22048 9404
rect 24121 9401 24133 9404
rect 24167 9432 24179 9435
rect 25041 9435 25099 9441
rect 25041 9432 25053 9435
rect 24167 9404 25053 9432
rect 24167 9401 24179 9404
rect 24121 9395 24179 9401
rect 25041 9401 25053 9404
rect 25087 9401 25099 9435
rect 25041 9395 25099 9401
rect 22005 9367 22063 9373
rect 22005 9333 22017 9367
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 24489 9367 24547 9373
rect 24489 9333 24501 9367
rect 24535 9364 24547 9367
rect 24765 9367 24823 9373
rect 24765 9364 24777 9367
rect 24535 9336 24777 9364
rect 24535 9333 24547 9336
rect 24489 9327 24547 9333
rect 24765 9333 24777 9336
rect 24811 9364 24823 9367
rect 24946 9364 24952 9376
rect 24811 9336 24952 9364
rect 24811 9333 24823 9336
rect 24765 9327 24823 9333
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2498 9160 2504 9172
rect 2455 9132 2504 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 2774 9120 2780 9172
rect 2832 9160 2838 9172
rect 7098 9160 7104 9172
rect 2832 9132 2877 9160
rect 7059 9132 7104 9160
rect 2832 9120 2838 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 7190 9120 7196 9172
rect 7248 9160 7254 9172
rect 7561 9163 7619 9169
rect 7248 9132 7293 9160
rect 7248 9120 7254 9132
rect 7561 9129 7573 9163
rect 7607 9160 7619 9163
rect 8018 9160 8024 9172
rect 7607 9132 8024 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 8352 9132 9321 9160
rect 8352 9120 8358 9132
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 9309 9123 9367 9129
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11701 9163 11759 9169
rect 11701 9160 11713 9163
rect 11480 9132 11713 9160
rect 11480 9120 11486 9132
rect 11701 9129 11713 9132
rect 11747 9129 11759 9163
rect 11701 9123 11759 9129
rect 14553 9163 14611 9169
rect 14553 9129 14565 9163
rect 14599 9160 14611 9163
rect 14826 9160 14832 9172
rect 14599 9132 14832 9160
rect 14599 9129 14611 9132
rect 14553 9123 14611 9129
rect 14826 9120 14832 9132
rect 14884 9120 14890 9172
rect 15010 9160 15016 9172
rect 14971 9132 15016 9160
rect 15010 9120 15016 9132
rect 15068 9160 15074 9172
rect 15286 9160 15292 9172
rect 15068 9132 15292 9160
rect 15068 9120 15074 9132
rect 15286 9120 15292 9132
rect 15344 9160 15350 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 15344 9132 16681 9160
rect 15344 9120 15350 9132
rect 16669 9129 16681 9132
rect 16715 9160 16727 9163
rect 17034 9160 17040 9172
rect 16715 9132 17040 9160
rect 16715 9129 16727 9132
rect 16669 9123 16727 9129
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 17313 9163 17371 9169
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17402 9160 17408 9172
rect 17359 9132 17408 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17402 9120 17408 9132
rect 17460 9160 17466 9172
rect 17589 9163 17647 9169
rect 17589 9160 17601 9163
rect 17460 9132 17601 9160
rect 17460 9120 17466 9132
rect 17589 9129 17601 9132
rect 17635 9129 17647 9163
rect 17589 9123 17647 9129
rect 18141 9163 18199 9169
rect 18141 9129 18153 9163
rect 18187 9160 18199 9163
rect 18598 9160 18604 9172
rect 18187 9132 18604 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 2958 9092 2964 9104
rect 1995 9064 2964 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 7116 9092 7144 9120
rect 7116 9064 7696 9092
rect 2866 9024 2872 9036
rect 2827 8996 2872 9024
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4154 9024 4160 9036
rect 4111 8996 4160 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4338 9033 4344 9036
rect 4332 9024 4344 9033
rect 4299 8996 4344 9024
rect 4332 8987 4344 8996
rect 4338 8984 4344 8987
rect 4396 8984 4402 9036
rect 7668 9024 7696 9064
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 10100 9064 10824 9092
rect 10100 9052 10106 9064
rect 9033 9027 9091 9033
rect 7668 8996 7788 9024
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 1946 8956 1952 8968
rect 1443 8928 1952 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 7760 8965 7788 8996
rect 9033 8993 9045 9027
rect 9079 9024 9091 9027
rect 9306 9024 9312 9036
rect 9079 8996 9312 9024
rect 9079 8993 9091 8996
rect 9033 8987 9091 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 10594 9033 10600 9036
rect 10588 9024 10600 9033
rect 10555 8996 10600 9024
rect 10588 8987 10600 8996
rect 10594 8984 10600 8987
rect 10652 8984 10658 9036
rect 10796 9024 10824 9064
rect 10870 9052 10876 9104
rect 10928 9092 10934 9104
rect 10928 9064 13860 9092
rect 10928 9052 10934 9064
rect 12250 9024 12256 9036
rect 10796 8996 12256 9024
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 13170 9024 13176 9036
rect 13131 8996 13176 9024
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13722 9024 13728 9036
rect 13311 8996 13728 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 6604 8928 7665 8956
rect 6604 8916 6610 8928
rect 7653 8925 7665 8928
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 10318 8956 10324 8968
rect 8628 8928 10324 8956
rect 8628 8916 8634 8928
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 13280 8956 13308 8987
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13832 9024 13860 9064
rect 15470 9052 15476 9104
rect 15528 9101 15534 9104
rect 15528 9095 15592 9101
rect 15528 9061 15546 9095
rect 15580 9061 15592 9095
rect 15528 9055 15592 9061
rect 15528 9052 15534 9055
rect 15838 9024 15844 9036
rect 13832 8996 15844 9024
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 17604 9024 17632 9123
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 21358 9160 21364 9172
rect 21319 9132 21364 9160
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 22370 9160 22376 9172
rect 22331 9132 22376 9160
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 22830 9160 22836 9172
rect 22791 9132 22836 9160
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 23106 9120 23112 9172
rect 23164 9160 23170 9172
rect 23201 9163 23259 9169
rect 23201 9160 23213 9163
rect 23164 9132 23213 9160
rect 23164 9120 23170 9132
rect 23201 9129 23213 9132
rect 23247 9129 23259 9163
rect 23658 9160 23664 9172
rect 23619 9132 23664 9160
rect 23201 9123 23259 9129
rect 23658 9120 23664 9132
rect 23716 9120 23722 9172
rect 18506 9092 18512 9104
rect 18467 9064 18512 9092
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 18616 9064 18828 9092
rect 18616 9024 18644 9064
rect 17604 8996 18644 9024
rect 12216 8928 13308 8956
rect 13357 8959 13415 8965
rect 12216 8916 12222 8928
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 3513 8891 3571 8897
rect 3513 8857 3525 8891
rect 3559 8888 3571 8891
rect 3970 8888 3976 8900
rect 3559 8860 3976 8888
rect 3559 8857 3571 8860
rect 3513 8851 3571 8857
rect 2314 8820 2320 8832
rect 2275 8792 2320 8820
rect 2314 8780 2320 8792
rect 2372 8780 2378 8832
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 3528 8820 3556 8851
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 13078 8848 13084 8900
rect 13136 8888 13142 8900
rect 13372 8888 13400 8919
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14792 8928 15301 8956
rect 14792 8916 14798 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 18322 8956 18328 8968
rect 17920 8928 18328 8956
rect 17920 8916 17926 8928
rect 18322 8916 18328 8928
rect 18380 8956 18386 8968
rect 18800 8965 18828 9064
rect 20162 9052 20168 9104
rect 20220 9092 20226 9104
rect 21266 9092 21272 9104
rect 20220 9064 21272 9092
rect 20220 9052 20226 9064
rect 21266 9052 21272 9064
rect 21324 9052 21330 9104
rect 22097 9095 22155 9101
rect 22097 9061 22109 9095
rect 22143 9092 22155 9095
rect 23124 9092 23152 9120
rect 22143 9064 23152 9092
rect 24020 9095 24078 9101
rect 22143 9061 22155 9064
rect 22097 9055 22155 9061
rect 24020 9061 24032 9095
rect 24066 9092 24078 9095
rect 24946 9092 24952 9104
rect 24066 9064 24952 9092
rect 24066 9061 24078 9064
rect 24020 9055 24078 9061
rect 24946 9052 24952 9064
rect 25004 9052 25010 9104
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 19484 8996 19717 9024
rect 19484 8984 19490 8996
rect 19705 8993 19717 8996
rect 19751 9024 19763 9027
rect 20257 9027 20315 9033
rect 20257 9024 20269 9027
rect 19751 8996 20269 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20257 8993 20269 8996
rect 20303 8993 20315 9027
rect 22646 9024 22652 9036
rect 22607 8996 22652 9024
rect 20257 8987 20315 8993
rect 22646 8984 22652 8996
rect 22704 8984 22710 9036
rect 23014 8984 23020 9036
rect 23072 9024 23078 9036
rect 23753 9027 23811 9033
rect 23753 9024 23765 9027
rect 23072 8996 23765 9024
rect 23072 8984 23078 8996
rect 23753 8993 23765 8996
rect 23799 8993 23811 9027
rect 23753 8987 23811 8993
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 18380 8928 18613 8956
rect 18380 8916 18386 8928
rect 18601 8925 18613 8928
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8956 18843 8959
rect 19242 8956 19248 8968
rect 18831 8928 19248 8956
rect 18831 8925 18843 8928
rect 18785 8919 18843 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21453 8959 21511 8965
rect 21453 8956 21465 8959
rect 21232 8928 21465 8956
rect 21232 8916 21238 8928
rect 21453 8925 21465 8928
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 13136 8860 13400 8888
rect 19337 8891 19395 8897
rect 13136 8848 13142 8860
rect 19337 8857 19349 8891
rect 19383 8888 19395 8891
rect 19518 8888 19524 8900
rect 19383 8860 19524 8888
rect 19383 8857 19395 8860
rect 19337 8851 19395 8857
rect 19518 8848 19524 8860
rect 19576 8888 19582 8900
rect 20901 8891 20959 8897
rect 20901 8888 20913 8891
rect 19576 8860 20913 8888
rect 19576 8848 19582 8860
rect 20901 8857 20913 8860
rect 20947 8857 20959 8891
rect 20901 8851 20959 8857
rect 2648 8792 3556 8820
rect 3881 8823 3939 8829
rect 2648 8780 2654 8792
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 4062 8820 4068 8832
rect 3927 8792 4068 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 5442 8820 5448 8832
rect 5403 8792 5448 8820
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8820 6147 8823
rect 6270 8820 6276 8832
rect 6135 8792 6276 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 6730 8820 6736 8832
rect 6691 8792 6736 8820
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 8294 8820 8300 8832
rect 8255 8792 8300 8820
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 10229 8823 10287 8829
rect 10229 8820 10241 8823
rect 10192 8792 10241 8820
rect 10192 8780 10198 8792
rect 10229 8789 10241 8792
rect 10275 8820 10287 8823
rect 10686 8820 10692 8832
rect 10275 8792 10692 8820
rect 10275 8789 10287 8792
rect 10229 8783 10287 8789
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 12437 8823 12495 8829
rect 12437 8820 12449 8823
rect 12400 8792 12449 8820
rect 12400 8780 12406 8792
rect 12437 8789 12449 8792
rect 12483 8789 12495 8823
rect 12437 8783 12495 8789
rect 12805 8823 12863 8829
rect 12805 8789 12817 8823
rect 12851 8820 12863 8823
rect 13722 8820 13728 8832
rect 12851 8792 13728 8820
rect 12851 8789 12863 8792
rect 12805 8783 12863 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 18049 8823 18107 8829
rect 13872 8792 13917 8820
rect 13872 8780 13878 8792
rect 18049 8789 18061 8823
rect 18095 8820 18107 8823
rect 18322 8820 18328 8832
rect 18095 8792 18328 8820
rect 18095 8789 18107 8792
rect 18049 8783 18107 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 19889 8823 19947 8829
rect 19889 8789 19901 8823
rect 19935 8820 19947 8823
rect 19978 8820 19984 8832
rect 19935 8792 19984 8820
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20714 8820 20720 8832
rect 20675 8792 20720 8820
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 25130 8820 25136 8832
rect 25091 8792 25136 8820
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 3605 8619 3663 8625
rect 3605 8616 3617 8619
rect 2556 8588 3617 8616
rect 2556 8576 2562 8588
rect 3605 8585 3617 8588
rect 3651 8616 3663 8619
rect 4338 8616 4344 8628
rect 3651 8588 4344 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 4338 8576 4344 8588
rect 4396 8616 4402 8628
rect 4525 8619 4583 8625
rect 4525 8616 4537 8619
rect 4396 8588 4537 8616
rect 4396 8576 4402 8588
rect 4525 8585 4537 8588
rect 4571 8585 4583 8619
rect 4525 8579 4583 8585
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7558 8616 7564 8628
rect 7147 8588 7564 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 7668 8588 10057 8616
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 3292 8520 5181 8548
rect 3292 8508 3298 8520
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5500 8452 5825 8480
rect 5500 8440 5506 8452
rect 5813 8449 5825 8452
rect 5859 8480 5871 8483
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5859 8452 6193 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6181 8449 6193 8452
rect 6227 8480 6239 8483
rect 6454 8480 6460 8492
rect 6227 8452 6460 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7668 8489 7696 8588
rect 10045 8585 10057 8588
rect 10091 8616 10103 8619
rect 10594 8616 10600 8628
rect 10091 8588 10600 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10594 8576 10600 8588
rect 10652 8616 10658 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10652 8588 10977 8616
rect 10652 8576 10658 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 13078 8576 13084 8628
rect 13136 8616 13142 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13136 8588 13829 8616
rect 13136 8576 13142 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 13817 8579 13875 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 18288 8588 19441 8616
rect 18288 8576 18294 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 20162 8616 20168 8628
rect 20123 8588 20168 8616
rect 19429 8579 19487 8585
rect 20162 8576 20168 8588
rect 20220 8576 20226 8628
rect 20533 8619 20591 8625
rect 20533 8585 20545 8619
rect 20579 8616 20591 8619
rect 21358 8616 21364 8628
rect 20579 8588 21364 8616
rect 20579 8585 20591 8588
rect 20533 8579 20591 8585
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 24946 8616 24952 8628
rect 24907 8588 24952 8616
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 25130 8576 25136 8628
rect 25188 8616 25194 8628
rect 25317 8619 25375 8625
rect 25317 8616 25329 8619
rect 25188 8588 25329 8616
rect 25188 8576 25194 8588
rect 25317 8585 25329 8588
rect 25363 8585 25375 8619
rect 25682 8616 25688 8628
rect 25643 8588 25688 8616
rect 25317 8579 25375 8585
rect 25682 8576 25688 8588
rect 25740 8576 25746 8628
rect 16114 8508 16120 8560
rect 16172 8548 16178 8560
rect 16301 8551 16359 8557
rect 16301 8548 16313 8551
rect 16172 8520 16313 8548
rect 16172 8508 16178 8520
rect 16301 8517 16313 8520
rect 16347 8517 16359 8551
rect 22002 8548 22008 8560
rect 21963 8520 22008 8548
rect 16301 8511 16359 8517
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 6788 8452 7665 8480
rect 6788 8440 6794 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 10318 8440 10324 8492
rect 10376 8480 10382 8492
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 10376 8452 10609 8480
rect 10376 8440 10382 8452
rect 10597 8449 10609 8452
rect 10643 8480 10655 8483
rect 11146 8480 11152 8492
rect 10643 8452 11152 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11330 8480 11336 8492
rect 11291 8452 11336 8480
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11572 8452 11897 8480
rect 11572 8440 11578 8452
rect 11885 8449 11897 8452
rect 11931 8480 11943 8483
rect 23109 8483 23167 8489
rect 11931 8452 12572 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 2130 8412 2136 8424
rect 2043 8384 2136 8412
rect 2130 8372 2136 8384
rect 2188 8412 2194 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 2188 8384 2237 8412
rect 2188 8372 2194 8384
rect 2225 8381 2237 8384
rect 2271 8412 2283 8415
rect 2271 8384 4292 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 4264 8356 4292 8384
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5316 8384 5549 8412
rect 5316 8372 5322 8384
rect 5537 8381 5549 8384
rect 5583 8412 5595 8415
rect 8018 8412 8024 8424
rect 5583 8384 8024 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8381 8723 8415
rect 8665 8375 8723 8381
rect 8932 8415 8990 8421
rect 8932 8381 8944 8415
rect 8978 8412 8990 8415
rect 9306 8412 9312 8424
rect 8978 8384 9312 8412
rect 8978 8381 8990 8384
rect 8932 8375 8990 8381
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 2470 8347 2528 8353
rect 2470 8344 2482 8347
rect 2372 8316 2482 8344
rect 2372 8304 2378 8316
rect 2470 8313 2482 8316
rect 2516 8313 2528 8347
rect 4246 8344 4252 8356
rect 4207 8316 4252 8344
rect 2470 8307 2528 8313
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 5077 8347 5135 8353
rect 5077 8313 5089 8347
rect 5123 8344 5135 8347
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5123 8316 5641 8344
rect 5123 8313 5135 8316
rect 5077 8307 5135 8313
rect 5629 8313 5641 8316
rect 5675 8344 5687 8347
rect 6546 8344 6552 8356
rect 5675 8316 6552 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7098 8304 7104 8356
rect 7156 8344 7162 8356
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 7156 8316 7573 8344
rect 7156 8304 7162 8316
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 7561 8307 7619 8313
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8481 8347 8539 8353
rect 8481 8344 8493 8347
rect 8352 8316 8493 8344
rect 8352 8304 8358 8316
rect 8481 8313 8493 8316
rect 8527 8344 8539 8347
rect 8570 8344 8576 8356
rect 8527 8316 8576 8344
rect 8527 8313 8539 8316
rect 8481 8307 8539 8313
rect 8570 8304 8576 8316
rect 8628 8344 8634 8356
rect 8680 8344 8708 8375
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 11164 8412 11192 8440
rect 12544 8424 12572 8452
rect 23109 8449 23121 8483
rect 23155 8480 23167 8483
rect 24210 8480 24216 8492
rect 23155 8452 24216 8480
rect 23155 8449 23167 8452
rect 23109 8443 23167 8449
rect 24210 8440 24216 8452
rect 24268 8480 24274 8492
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 24268 8452 24409 8480
rect 24268 8440 24274 8452
rect 24397 8449 24409 8452
rect 24443 8449 24455 8483
rect 24578 8480 24584 8492
rect 24491 8452 24584 8480
rect 24397 8443 24455 8449
rect 24578 8440 24584 8452
rect 24636 8480 24642 8492
rect 25148 8480 25176 8576
rect 24636 8452 25176 8480
rect 24636 8440 24642 8452
rect 12342 8412 12348 8424
rect 11164 8384 12348 8412
rect 12342 8372 12348 8384
rect 12400 8412 12406 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12400 8384 12449 8412
rect 12400 8372 12406 8384
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 12158 8344 12164 8356
rect 8628 8316 8708 8344
rect 12119 8316 12164 8344
rect 8628 8304 8634 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 1765 8279 1823 8285
rect 1765 8245 1777 8279
rect 1811 8276 1823 8279
rect 3050 8276 3056 8288
rect 1811 8248 3056 8276
rect 1811 8245 1823 8248
rect 1765 8239 1823 8245
rect 3050 8236 3056 8248
rect 3108 8236 3114 8288
rect 7466 8276 7472 8288
rect 7427 8248 7472 8276
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 8110 8276 8116 8288
rect 8071 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 12452 8276 12480 8375
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 12693 8415 12751 8421
rect 12693 8412 12705 8415
rect 12584 8384 12705 8412
rect 12584 8372 12590 8384
rect 12693 8381 12705 8384
rect 12739 8381 12751 8415
rect 12693 8375 12751 8381
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8412 14703 8415
rect 14734 8412 14740 8424
rect 14691 8384 14740 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 14734 8372 14740 8384
rect 14792 8412 14798 8424
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14792 8384 14933 8412
rect 14792 8372 14798 8384
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 17954 8412 17960 8424
rect 17543 8384 17960 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 17954 8372 17960 8384
rect 18012 8412 18018 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 18012 8384 18061 8412
rect 18012 8372 18018 8384
rect 18049 8381 18061 8384
rect 18095 8412 18107 8415
rect 20622 8412 20628 8424
rect 18095 8384 20628 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 25498 8412 25504 8424
rect 25459 8384 25504 8412
rect 25498 8372 25504 8384
rect 25556 8412 25562 8424
rect 26053 8415 26111 8421
rect 26053 8412 26065 8415
rect 25556 8384 26065 8412
rect 25556 8372 25562 8384
rect 26053 8381 26065 8384
rect 26099 8381 26111 8415
rect 26053 8375 26111 8381
rect 14461 8347 14519 8353
rect 14461 8313 14473 8347
rect 14507 8344 14519 8347
rect 15188 8347 15246 8353
rect 14507 8316 15148 8344
rect 14507 8313 14519 8316
rect 14461 8307 14519 8313
rect 14645 8279 14703 8285
rect 14645 8276 14657 8279
rect 12452 8248 14657 8276
rect 14645 8245 14657 8248
rect 14691 8276 14703 8279
rect 14737 8279 14795 8285
rect 14737 8276 14749 8279
rect 14691 8248 14749 8276
rect 14691 8245 14703 8248
rect 14645 8239 14703 8245
rect 14737 8245 14749 8248
rect 14783 8245 14795 8279
rect 15120 8276 15148 8316
rect 15188 8313 15200 8347
rect 15234 8344 15246 8347
rect 15286 8344 15292 8356
rect 15234 8316 15292 8344
rect 15234 8313 15246 8316
rect 15188 8307 15246 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17037 8347 17095 8353
rect 17037 8344 17049 8347
rect 16632 8316 17049 8344
rect 16632 8304 16638 8316
rect 17037 8313 17049 8316
rect 17083 8344 17095 8347
rect 17862 8344 17868 8356
rect 17083 8316 17868 8344
rect 17083 8313 17095 8316
rect 17037 8307 17095 8313
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 18322 8353 18328 8356
rect 18316 8344 18328 8353
rect 18235 8316 18328 8344
rect 18316 8307 18328 8316
rect 18380 8344 18386 8356
rect 19242 8344 19248 8356
rect 18380 8316 19248 8344
rect 18322 8304 18328 8307
rect 18380 8304 18386 8316
rect 19242 8304 19248 8316
rect 19300 8304 19306 8356
rect 20714 8304 20720 8356
rect 20772 8344 20778 8356
rect 20870 8347 20928 8353
rect 20870 8344 20882 8347
rect 20772 8316 20882 8344
rect 20772 8304 20778 8316
rect 20870 8313 20882 8316
rect 20916 8344 20928 8347
rect 22646 8344 22652 8356
rect 20916 8316 22140 8344
rect 22607 8316 22652 8344
rect 20916 8313 20928 8316
rect 20870 8307 20928 8313
rect 15470 8276 15476 8288
rect 15120 8248 15476 8276
rect 14737 8239 14795 8245
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 22112 8276 22140 8316
rect 22646 8304 22652 8316
rect 22704 8304 22710 8356
rect 23474 8344 23480 8356
rect 23435 8316 23480 8344
rect 23474 8304 23480 8316
rect 23532 8344 23538 8356
rect 24305 8347 24363 8353
rect 24305 8344 24317 8347
rect 23532 8316 24317 8344
rect 23532 8304 23538 8316
rect 24305 8313 24317 8316
rect 24351 8313 24363 8347
rect 24305 8307 24363 8313
rect 22278 8276 22284 8288
rect 22112 8248 22284 8276
rect 22278 8236 22284 8248
rect 22336 8236 22342 8288
rect 23934 8276 23940 8288
rect 23895 8248 23940 8276
rect 23934 8236 23940 8248
rect 23992 8236 23998 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 1452 8044 2237 8072
rect 1452 8032 1458 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3237 8075 3295 8081
rect 3237 8072 3249 8075
rect 2924 8044 3249 8072
rect 2924 8032 2930 8044
rect 3237 8041 3249 8044
rect 3283 8041 3295 8075
rect 3237 8035 3295 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4706 8072 4712 8084
rect 4571 8044 4712 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5810 8072 5816 8084
rect 5771 8044 5816 8072
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 7524 8044 7573 8072
rect 7524 8032 7530 8044
rect 7561 8041 7573 8044
rect 7607 8072 7619 8075
rect 8754 8072 8760 8084
rect 7607 8044 8760 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 10686 8072 10692 8084
rect 10647 8044 10692 8072
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13170 8072 13176 8084
rect 13131 8044 13176 8072
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13320 8044 13645 8072
rect 13320 8032 13326 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14001 8075 14059 8081
rect 14001 8072 14013 8075
rect 13780 8044 14013 8072
rect 13780 8032 13786 8044
rect 14001 8041 14013 8044
rect 14047 8041 14059 8075
rect 14001 8035 14059 8041
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 14792 8044 15485 8072
rect 14792 8032 14798 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 15473 8035 15531 8041
rect 16117 8075 16175 8081
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16574 8072 16580 8084
rect 16163 8044 16580 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 17092 8044 17141 8072
rect 17092 8032 17098 8044
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 17129 8035 17187 8041
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 17770 8072 17776 8084
rect 17727 8044 17776 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18141 8075 18199 8081
rect 18141 8072 18153 8075
rect 18012 8044 18153 8072
rect 18012 8032 18018 8044
rect 18141 8041 18153 8044
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 18564 8044 18705 8072
rect 18564 8032 18570 8044
rect 18693 8041 18705 8044
rect 18739 8041 18751 8075
rect 18693 8035 18751 8041
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 18840 8044 19257 8072
rect 18840 8032 18846 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 19245 8035 19303 8041
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 19576 8044 19625 8072
rect 19576 8032 19582 8044
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 20622 8032 20628 8084
rect 20680 8072 20686 8084
rect 20717 8075 20775 8081
rect 20717 8072 20729 8075
rect 20680 8044 20729 8072
rect 20680 8032 20686 8044
rect 20717 8041 20729 8044
rect 20763 8072 20775 8075
rect 20806 8072 20812 8084
rect 20763 8044 20812 8072
rect 20763 8041 20775 8044
rect 20717 8035 20775 8041
rect 20806 8032 20812 8044
rect 20864 8032 20870 8084
rect 22278 8072 22284 8084
rect 22239 8044 22284 8072
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 23477 8075 23535 8081
rect 23477 8041 23489 8075
rect 23523 8072 23535 8075
rect 23934 8072 23940 8084
rect 23523 8044 23940 8072
rect 23523 8041 23535 8044
rect 23477 8035 23535 8041
rect 23934 8032 23940 8044
rect 23992 8032 23998 8084
rect 2133 8007 2191 8013
rect 2133 7973 2145 8007
rect 2179 8004 2191 8007
rect 2682 8004 2688 8016
rect 2179 7976 2688 8004
rect 2179 7973 2191 7976
rect 2133 7967 2191 7973
rect 2682 7964 2688 7976
rect 2740 7964 2746 8016
rect 3050 7964 3056 8016
rect 3108 8004 3114 8016
rect 8662 8004 8668 8016
rect 3108 7976 8668 8004
rect 3108 7964 3114 7976
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 10134 8004 10140 8016
rect 10095 7976 10140 8004
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 11422 8013 11428 8016
rect 11416 8004 11428 8013
rect 11383 7976 11428 8004
rect 11416 7967 11428 7976
rect 11422 7964 11428 7967
rect 11480 7964 11486 8016
rect 24204 8007 24262 8013
rect 24204 7973 24216 8007
rect 24250 8004 24262 8007
rect 24578 8004 24584 8016
rect 24250 7976 24584 8004
rect 24250 7973 24262 7976
rect 24204 7967 24262 7973
rect 24578 7964 24584 7976
rect 24636 7964 24642 8016
rect 2590 7936 2596 7948
rect 2551 7908 2596 7936
rect 2590 7896 2596 7908
rect 2648 7896 2654 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4212 7908 4445 7936
rect 4212 7896 4218 7908
rect 4433 7905 4445 7908
rect 4479 7905 4491 7939
rect 6178 7936 6184 7948
rect 6139 7908 6184 7936
rect 4433 7899 4491 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 6454 7936 6460 7948
rect 6319 7908 6460 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 6454 7896 6460 7908
rect 6512 7936 6518 7948
rect 6638 7936 6644 7948
rect 6512 7908 6644 7936
rect 6512 7896 6518 7908
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 8018 7936 8024 7948
rect 7979 7908 8024 7936
rect 8018 7896 8024 7908
rect 8076 7896 8082 7948
rect 12618 7936 12624 7948
rect 8128 7908 12624 7936
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 4614 7868 4620 7880
rect 4575 7840 4620 7868
rect 2777 7831 2835 7837
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2498 7800 2504 7812
rect 2372 7772 2504 7800
rect 2372 7760 2378 7772
rect 2498 7760 2504 7772
rect 2556 7800 2562 7812
rect 2792 7800 2820 7831
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 2556 7772 2820 7800
rect 2556 7760 2562 7772
rect 3326 7760 3332 7812
rect 3384 7800 3390 7812
rect 3878 7800 3884 7812
rect 3384 7772 3884 7800
rect 3384 7760 3390 7772
rect 3878 7760 3884 7772
rect 3936 7800 3942 7812
rect 4065 7803 4123 7809
rect 4065 7800 4077 7803
rect 3936 7772 4077 7800
rect 3936 7760 3942 7772
rect 4065 7769 4077 7772
rect 4111 7769 4123 7803
rect 4065 7763 4123 7769
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7800 5779 7803
rect 6380 7800 6408 7831
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 8128 7877 8156 7908
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 14090 7936 14096 7948
rect 14003 7908 14096 7936
rect 14090 7896 14096 7908
rect 14148 7936 14154 7948
rect 14550 7936 14556 7948
rect 14148 7908 14556 7936
rect 14148 7896 14154 7908
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 16022 7896 16028 7948
rect 16080 7936 16086 7948
rect 16485 7939 16543 7945
rect 16485 7936 16497 7939
rect 16080 7908 16497 7936
rect 16080 7896 16086 7908
rect 16485 7905 16497 7908
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 16666 7936 16672 7948
rect 16623 7908 16672 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 18012 7908 18061 7936
rect 18012 7896 18018 7908
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7936 19211 7939
rect 19242 7936 19248 7948
rect 19199 7908 19248 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 21174 7945 21180 7948
rect 20349 7939 20407 7945
rect 20349 7905 20361 7939
rect 20395 7936 20407 7939
rect 21168 7936 21180 7945
rect 20395 7908 21180 7936
rect 20395 7905 20407 7908
rect 20349 7899 20407 7905
rect 21168 7899 21180 7908
rect 21174 7896 21180 7899
rect 21232 7896 21238 7948
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7800 7840 8125 7868
rect 7800 7828 7806 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7868 8355 7871
rect 11146 7868 11152 7880
rect 8343 7840 8800 7868
rect 11107 7840 11152 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 6914 7800 6920 7812
rect 5767 7772 6920 7800
rect 5767 7769 5779 7772
rect 5721 7763 5779 7769
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 8772 7809 8800 7840
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 16761 7871 16819 7877
rect 14240 7840 14285 7868
rect 14240 7828 14246 7840
rect 16761 7837 16773 7871
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 18138 7868 18144 7880
rect 17635 7840 18144 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 8757 7803 8815 7809
rect 8757 7769 8769 7803
rect 8803 7800 8815 7803
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8803 7772 9321 7800
rect 8803 7769 8815 7772
rect 8757 7763 8815 7769
rect 9309 7769 9321 7772
rect 9355 7800 9367 7803
rect 10134 7800 10140 7812
rect 9355 7772 10140 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 16025 7803 16083 7809
rect 16025 7769 16037 7803
rect 16071 7800 16083 7803
rect 16776 7800 16804 7831
rect 18138 7828 18144 7840
rect 18196 7868 18202 7880
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 18196 7840 18245 7868
rect 18196 7828 18202 7840
rect 18233 7837 18245 7840
rect 18279 7837 18291 7871
rect 19702 7868 19708 7880
rect 19663 7840 19708 7868
rect 18233 7831 18291 7837
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 19794 7828 19800 7880
rect 19852 7868 19858 7880
rect 20714 7868 20720 7880
rect 19852 7840 20720 7868
rect 19852 7828 19858 7840
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20864 7840 20913 7868
rect 20864 7828 20870 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 23937 7871 23995 7877
rect 23937 7868 23949 7871
rect 20901 7831 20959 7837
rect 23768 7840 23949 7868
rect 18322 7800 18328 7812
rect 16071 7772 18328 7800
rect 16071 7769 16083 7772
rect 16025 7763 16083 7769
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 1394 7692 1400 7744
rect 1452 7732 1458 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1452 7704 1593 7732
rect 1452 7692 1458 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 3786 7732 3792 7744
rect 3747 7704 3792 7732
rect 1581 7695 1639 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 7098 7732 7104 7744
rect 7059 7704 7104 7732
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7650 7732 7656 7744
rect 7611 7704 7656 7732
rect 7650 7692 7656 7704
rect 7708 7692 7714 7744
rect 9858 7732 9864 7744
rect 9819 7704 9864 7732
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13449 7735 13507 7741
rect 13449 7732 13461 7735
rect 13044 7704 13461 7732
rect 13044 7692 13050 7704
rect 13449 7701 13461 7704
rect 13495 7701 13507 7735
rect 14642 7732 14648 7744
rect 14603 7704 14648 7732
rect 13449 7695 13507 7701
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14792 7704 15025 7732
rect 14792 7692 14798 7704
rect 15013 7701 15025 7704
rect 15059 7701 15071 7735
rect 22830 7732 22836 7744
rect 22791 7704 22836 7732
rect 15013 7695 15071 7701
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 23474 7692 23480 7744
rect 23532 7732 23538 7744
rect 23768 7741 23796 7840
rect 23937 7837 23949 7840
rect 23983 7837 23995 7871
rect 23937 7831 23995 7837
rect 23753 7735 23811 7741
rect 23753 7732 23765 7735
rect 23532 7704 23765 7732
rect 23532 7692 23538 7704
rect 23753 7701 23765 7704
rect 23799 7701 23811 7735
rect 25314 7732 25320 7744
rect 25275 7704 25320 7732
rect 23753 7695 23811 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 2130 7528 2136 7540
rect 2087 7500 2136 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 4522 7528 4528 7540
rect 4435 7500 4528 7528
rect 4522 7488 4528 7500
rect 4580 7528 4586 7540
rect 4706 7528 4712 7540
rect 4580 7500 4712 7528
rect 4580 7488 4586 7500
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 6196 7500 8217 7528
rect 2148 7401 2176 7488
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 5169 7463 5227 7469
rect 5169 7460 5181 7463
rect 4028 7432 5181 7460
rect 4028 7420 4034 7432
rect 5169 7429 5181 7432
rect 5215 7429 5227 7463
rect 5169 7423 5227 7429
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7361 2191 7395
rect 4154 7392 4160 7404
rect 4115 7364 4160 7392
rect 2133 7355 2191 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 5810 7392 5816 7404
rect 5723 7364 5816 7392
rect 5810 7352 5816 7364
rect 5868 7392 5874 7404
rect 6196 7392 6224 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 10689 7531 10747 7537
rect 10689 7528 10701 7531
rect 9732 7500 10701 7528
rect 9732 7488 9738 7500
rect 10689 7497 10701 7500
rect 10735 7497 10747 7531
rect 10689 7491 10747 7497
rect 11146 7488 11152 7540
rect 11204 7488 11210 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11977 7531 12035 7537
rect 11977 7528 11989 7531
rect 11480 7500 11989 7528
rect 11480 7488 11486 7500
rect 11977 7497 11989 7500
rect 12023 7497 12035 7531
rect 13354 7528 13360 7540
rect 13267 7500 13360 7528
rect 11977 7491 12035 7497
rect 13354 7488 13360 7500
rect 13412 7528 13418 7540
rect 14182 7528 14188 7540
rect 13412 7500 14188 7528
rect 13412 7488 13418 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 16298 7528 16304 7540
rect 16259 7500 16304 7528
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 17313 7531 17371 7537
rect 17313 7528 17325 7531
rect 16724 7500 17325 7528
rect 16724 7488 16730 7500
rect 17313 7497 17325 7500
rect 17359 7497 17371 7531
rect 17313 7491 17371 7497
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 17773 7531 17831 7537
rect 17773 7528 17785 7531
rect 17644 7500 17785 7528
rect 17644 7488 17650 7500
rect 17773 7497 17785 7500
rect 17819 7528 17831 7531
rect 17819 7500 18552 7528
rect 17819 7497 17831 7500
rect 17773 7491 17831 7497
rect 6273 7463 6331 7469
rect 6273 7429 6285 7463
rect 6319 7460 6331 7463
rect 6454 7460 6460 7472
rect 6319 7432 6460 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 6454 7420 6460 7432
rect 6512 7420 6518 7472
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 8757 7463 8815 7469
rect 8757 7460 8769 7463
rect 8076 7432 8769 7460
rect 8076 7420 8082 7432
rect 8757 7429 8769 7432
rect 8803 7429 8815 7463
rect 9306 7460 9312 7472
rect 9267 7432 9312 7460
rect 8757 7423 8815 7429
rect 9306 7420 9312 7432
rect 9364 7420 9370 7472
rect 11164 7460 11192 7488
rect 11609 7463 11667 7469
rect 11609 7460 11621 7463
rect 11164 7432 11621 7460
rect 11609 7429 11621 7432
rect 11655 7460 11667 7463
rect 13633 7463 13691 7469
rect 13633 7460 13645 7463
rect 11655 7432 13645 7460
rect 11655 7429 11667 7432
rect 11609 7423 11667 7429
rect 13633 7429 13645 7432
rect 13679 7460 13691 7463
rect 15197 7463 15255 7469
rect 13679 7432 13860 7460
rect 13679 7429 13691 7432
rect 13633 7423 13691 7429
rect 5868 7364 6224 7392
rect 9953 7395 10011 7401
rect 5868 7352 5874 7364
rect 9953 7361 9965 7395
rect 9999 7392 10011 7395
rect 10134 7392 10140 7404
rect 9999 7364 10140 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 13170 7392 13176 7404
rect 11195 7364 13176 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13832 7401 13860 7432
rect 15197 7429 15209 7463
rect 15243 7460 15255 7463
rect 15470 7460 15476 7472
rect 15243 7432 15476 7460
rect 15243 7429 15255 7432
rect 15197 7423 15255 7429
rect 15470 7420 15476 7432
rect 15528 7460 15534 7472
rect 16390 7460 16396 7472
rect 15528 7432 16396 7460
rect 15528 7420 15534 7432
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17034 7392 17040 7404
rect 16991 7364 17040 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 18524 7401 18552 7500
rect 19702 7488 19708 7540
rect 19760 7528 19766 7540
rect 20254 7528 20260 7540
rect 19760 7500 20260 7528
rect 19760 7488 19766 7500
rect 20254 7488 20260 7500
rect 20312 7528 20318 7540
rect 20717 7531 20775 7537
rect 20717 7528 20729 7531
rect 20312 7500 20729 7528
rect 20312 7488 20318 7500
rect 20717 7497 20729 7500
rect 20763 7497 20775 7531
rect 20717 7491 20775 7497
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 21729 7531 21787 7537
rect 21729 7528 21741 7531
rect 20864 7500 21741 7528
rect 20864 7488 20870 7500
rect 21729 7497 21741 7500
rect 21775 7497 21787 7531
rect 21729 7491 21787 7497
rect 23566 7488 23572 7540
rect 23624 7528 23630 7540
rect 23661 7531 23719 7537
rect 23661 7528 23673 7531
rect 23624 7500 23673 7528
rect 23624 7488 23630 7500
rect 23661 7497 23673 7500
rect 23707 7497 23719 7531
rect 25130 7528 25136 7540
rect 25091 7500 25136 7528
rect 23661 7491 23719 7497
rect 25130 7488 25136 7500
rect 25188 7488 25194 7540
rect 19337 7463 19395 7469
rect 19337 7429 19349 7463
rect 19383 7460 19395 7463
rect 19794 7460 19800 7472
rect 19383 7432 19800 7460
rect 19383 7429 19395 7432
rect 19337 7423 19395 7429
rect 19794 7420 19800 7432
rect 19852 7420 19858 7472
rect 23477 7463 23535 7469
rect 23477 7429 23489 7463
rect 23523 7460 23535 7463
rect 23750 7460 23756 7472
rect 23523 7432 23756 7460
rect 23523 7429 23535 7432
rect 23477 7423 23535 7429
rect 23750 7420 23756 7432
rect 23808 7420 23814 7472
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 19242 7392 19248 7404
rect 18739 7364 19248 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 21174 7352 21180 7404
rect 21232 7392 21238 7404
rect 21361 7395 21419 7401
rect 21361 7392 21373 7395
rect 21232 7364 21373 7392
rect 21232 7352 21238 7364
rect 21361 7361 21373 7364
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 5534 7324 5540 7336
rect 5495 7296 5540 7324
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 5994 7324 6000 7336
rect 5675 7296 6000 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6178 7284 6184 7336
rect 6236 7284 6242 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6564 7296 6837 7324
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 2378 7259 2436 7265
rect 2378 7256 2390 7259
rect 1719 7228 2390 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 2378 7225 2390 7228
rect 2424 7256 2436 7259
rect 3234 7256 3240 7268
rect 2424 7228 3240 7256
rect 2424 7225 2436 7228
rect 2378 7219 2436 7225
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 6196 7256 6224 7284
rect 5123 7228 6224 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 3510 7188 3516 7200
rect 3471 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 6564 7197 6592 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7081 7327 7139 7333
rect 7081 7324 7093 7327
rect 6972 7296 7093 7324
rect 6972 7284 6978 7296
rect 7081 7293 7093 7296
rect 7127 7293 7139 7327
rect 7081 7287 7139 7293
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10321 7327 10379 7333
rect 10321 7324 10333 7327
rect 9732 7296 10333 7324
rect 9732 7284 9738 7296
rect 10321 7293 10333 7296
rect 10367 7293 10379 7327
rect 14084 7327 14142 7333
rect 10321 7287 10379 7293
rect 10428 7296 13584 7324
rect 9769 7259 9827 7265
rect 9769 7256 9781 7259
rect 9140 7228 9781 7256
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 5592 7160 6561 7188
rect 5592 7148 5598 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 6549 7151 6607 7157
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 9140 7197 9168 7228
rect 9769 7225 9781 7228
rect 9815 7225 9827 7259
rect 9769 7219 9827 7225
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 8352 7160 9137 7188
rect 8352 7148 8358 7160
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 9125 7151 9183 7157
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 9677 7191 9735 7197
rect 9677 7188 9689 7191
rect 9364 7160 9689 7188
rect 9364 7148 9370 7160
rect 9677 7157 9689 7160
rect 9723 7188 9735 7191
rect 10428 7188 10456 7296
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 13078 7256 13084 7268
rect 12759 7228 13084 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 13078 7216 13084 7228
rect 13136 7216 13142 7268
rect 13556 7256 13584 7296
rect 14084 7293 14096 7327
rect 14130 7324 14142 7327
rect 14642 7324 14648 7336
rect 14130 7296 14648 7324
rect 14130 7293 14142 7296
rect 14084 7287 14142 7293
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 15838 7324 15844 7336
rect 15751 7296 15844 7324
rect 15838 7284 15844 7296
rect 15896 7324 15902 7336
rect 16666 7324 16672 7336
rect 15896 7296 16672 7324
rect 15896 7284 15902 7296
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18104 7296 18429 7324
rect 18104 7284 18110 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 19610 7324 19616 7336
rect 19571 7296 19616 7324
rect 18417 7287 18475 7293
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 20162 7324 20168 7336
rect 20123 7296 20168 7324
rect 20162 7284 20168 7296
rect 20220 7324 20226 7336
rect 21266 7324 21272 7336
rect 20220 7296 21272 7324
rect 20220 7284 20226 7296
rect 16022 7256 16028 7268
rect 13556 7228 16028 7256
rect 16022 7216 16028 7228
rect 16080 7256 16086 7268
rect 16117 7259 16175 7265
rect 16117 7256 16129 7259
rect 16080 7228 16129 7256
rect 16080 7216 16086 7228
rect 16117 7225 16129 7228
rect 16163 7225 16175 7259
rect 16117 7219 16175 7225
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 16264 7228 16773 7256
rect 16264 7216 16270 7228
rect 16761 7225 16773 7228
rect 16807 7225 16819 7259
rect 16761 7219 16819 7225
rect 18966 7216 18972 7268
rect 19024 7256 19030 7268
rect 21192 7265 21220 7296
rect 21266 7284 21272 7296
rect 21324 7284 21330 7336
rect 21376 7324 21404 7355
rect 23934 7352 23940 7404
rect 23992 7392 23998 7404
rect 24121 7395 24179 7401
rect 24121 7392 24133 7395
rect 23992 7364 24133 7392
rect 23992 7352 23998 7364
rect 24121 7361 24133 7364
rect 24167 7361 24179 7395
rect 24302 7392 24308 7404
rect 24215 7364 24308 7392
rect 24121 7355 24179 7361
rect 24302 7352 24308 7364
rect 24360 7392 24366 7404
rect 25314 7392 25320 7404
rect 24360 7364 25320 7392
rect 24360 7352 24366 7364
rect 25314 7352 25320 7364
rect 25372 7352 25378 7404
rect 22094 7324 22100 7336
rect 21376 7296 22100 7324
rect 22094 7284 22100 7296
rect 22152 7324 22158 7336
rect 22465 7327 22523 7333
rect 22152 7296 22245 7324
rect 22152 7284 22158 7296
rect 22465 7293 22477 7327
rect 22511 7324 22523 7327
rect 22922 7324 22928 7336
rect 22511 7296 22928 7324
rect 22511 7293 22523 7296
rect 22465 7287 22523 7293
rect 22922 7284 22928 7296
rect 22980 7284 22986 7336
rect 23106 7324 23112 7336
rect 23019 7296 23112 7324
rect 23106 7284 23112 7296
rect 23164 7324 23170 7336
rect 24320 7324 24348 7352
rect 25222 7324 25228 7336
rect 23164 7296 24348 7324
rect 25183 7296 25228 7324
rect 23164 7284 23170 7296
rect 25222 7284 25228 7296
rect 25280 7324 25286 7336
rect 25777 7327 25835 7333
rect 25777 7324 25789 7327
rect 25280 7296 25789 7324
rect 25280 7284 25286 7296
rect 25777 7293 25789 7296
rect 25823 7293 25835 7327
rect 25777 7287 25835 7293
rect 20533 7259 20591 7265
rect 20533 7256 20545 7259
rect 19024 7228 20545 7256
rect 19024 7216 19030 7228
rect 20533 7225 20545 7228
rect 20579 7256 20591 7259
rect 21085 7259 21143 7265
rect 21085 7256 21097 7259
rect 20579 7228 21097 7256
rect 20579 7225 20591 7228
rect 20533 7219 20591 7225
rect 21085 7225 21097 7228
rect 21131 7225 21143 7259
rect 21085 7219 21143 7225
rect 21177 7259 21235 7265
rect 21177 7225 21189 7259
rect 21223 7225 21235 7259
rect 21177 7219 21235 7225
rect 12802 7188 12808 7200
rect 9723 7160 10456 7188
rect 12763 7160 12808 7188
rect 9723 7157 9735 7160
rect 9677 7151 9735 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 18012 7160 18061 7188
rect 18012 7148 18018 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 18049 7151 18107 7157
rect 19797 7191 19855 7197
rect 19797 7157 19809 7191
rect 19843 7188 19855 7191
rect 20346 7188 20352 7200
rect 19843 7160 20352 7188
rect 19843 7157 19855 7160
rect 19797 7151 19855 7157
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 21100 7188 21128 7219
rect 23750 7216 23756 7268
rect 23808 7256 23814 7268
rect 24029 7259 24087 7265
rect 24029 7256 24041 7259
rect 23808 7228 24041 7256
rect 23808 7216 23814 7228
rect 24029 7225 24041 7228
rect 24075 7225 24087 7259
rect 24029 7219 24087 7225
rect 21358 7188 21364 7200
rect 21100 7160 21364 7188
rect 21358 7148 21364 7160
rect 21416 7148 21422 7200
rect 22649 7191 22707 7197
rect 22649 7157 22661 7191
rect 22695 7188 22707 7191
rect 23290 7188 23296 7200
rect 22695 7160 23296 7188
rect 22695 7157 22707 7160
rect 22649 7151 22707 7157
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 23566 7148 23572 7200
rect 23624 7188 23630 7200
rect 24673 7191 24731 7197
rect 24673 7188 24685 7191
rect 23624 7160 24685 7188
rect 23624 7148 23630 7160
rect 24673 7157 24685 7160
rect 24719 7157 24731 7191
rect 25406 7188 25412 7200
rect 25367 7160 25412 7188
rect 24673 7151 24731 7157
rect 25406 7148 25412 7160
rect 25464 7148 25470 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 2409 6987 2467 6993
rect 2409 6953 2421 6987
rect 2455 6984 2467 6987
rect 2590 6984 2596 6996
rect 2455 6956 2596 6984
rect 2455 6953 2467 6956
rect 2409 6947 2467 6953
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 7006 6984 7012 6996
rect 4028 6956 7012 6984
rect 4028 6944 4034 6956
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 10962 6944 10968 6996
rect 11020 6984 11026 6996
rect 11606 6984 11612 6996
rect 11020 6956 11612 6984
rect 11020 6944 11026 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 12158 6984 12164 6996
rect 12071 6956 12164 6984
rect 12158 6944 12164 6956
rect 12216 6984 12222 6996
rect 13354 6984 13360 6996
rect 12216 6956 13360 6984
rect 12216 6944 12222 6956
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 18046 6984 18052 6996
rect 18007 6956 18052 6984
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18874 6984 18880 6996
rect 18835 6956 18880 6984
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 20254 6984 20260 6996
rect 20215 6956 20260 6984
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 22094 6984 22100 6996
rect 20763 6956 22100 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 22094 6944 22100 6956
rect 22152 6984 22158 6996
rect 22281 6987 22339 6993
rect 22281 6984 22293 6987
rect 22152 6956 22293 6984
rect 22152 6944 22158 6956
rect 22281 6953 22293 6956
rect 22327 6953 22339 6987
rect 22281 6947 22339 6953
rect 22922 6944 22928 6996
rect 22980 6984 22986 6996
rect 23201 6987 23259 6993
rect 23201 6984 23213 6987
rect 22980 6956 23213 6984
rect 22980 6944 22986 6956
rect 23201 6953 23213 6956
rect 23247 6953 23259 6987
rect 23201 6947 23259 6953
rect 5712 6919 5770 6925
rect 5712 6916 5724 6919
rect 5644 6888 5724 6916
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 2188 6820 2789 6848
rect 2188 6808 2194 6820
rect 2777 6817 2789 6820
rect 2823 6848 2835 6851
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 2823 6820 4077 6848
rect 2823 6817 2835 6820
rect 2777 6811 2835 6817
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5534 6848 5540 6860
rect 5307 6820 5540 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5534 6808 5540 6820
rect 5592 6848 5598 6860
rect 5644 6848 5672 6888
rect 5712 6885 5724 6888
rect 5758 6916 5770 6919
rect 5810 6916 5816 6928
rect 5758 6888 5816 6916
rect 5758 6885 5770 6888
rect 5712 6879 5770 6885
rect 5810 6876 5816 6888
rect 5868 6876 5874 6928
rect 5994 6876 6000 6928
rect 6052 6916 6058 6928
rect 8297 6919 8355 6925
rect 6052 6888 6868 6916
rect 6052 6876 6058 6888
rect 5592 6820 5672 6848
rect 6840 6848 6868 6888
rect 8297 6885 8309 6919
rect 8343 6916 8355 6919
rect 9858 6916 9864 6928
rect 8343 6888 9864 6916
rect 8343 6885 8355 6888
rect 8297 6879 8355 6885
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 10980 6888 13185 6916
rect 6840 6820 7972 6848
rect 5592 6808 5598 6820
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6780 2007 6783
rect 2406 6780 2412 6792
rect 1995 6752 2412 6780
rect 1995 6749 2007 6752
rect 1949 6743 2007 6749
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 2866 6780 2872 6792
rect 2827 6752 2872 6780
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3510 6780 3516 6792
rect 3099 6752 3516 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 2424 6712 2452 6740
rect 3068 6712 3096 6743
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 2424 6684 3096 6712
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 3292 6684 3924 6712
rect 3292 6672 3298 6684
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 3896 6653 3924 6684
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 7944 6721 7972 6820
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 8076 6820 8401 6848
rect 8076 6808 8082 6820
rect 8389 6817 8401 6820
rect 8435 6848 8447 6851
rect 9674 6848 9680 6860
rect 8435 6820 9680 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 9769 6851 9827 6857
rect 9769 6817 9781 6851
rect 9815 6848 9827 6851
rect 10980 6848 11008 6888
rect 13173 6885 13185 6888
rect 13219 6916 13231 6919
rect 13725 6919 13783 6925
rect 13725 6916 13737 6919
rect 13219 6888 13737 6916
rect 13219 6885 13231 6888
rect 13173 6879 13231 6885
rect 13725 6885 13737 6888
rect 13771 6885 13783 6919
rect 15102 6916 15108 6928
rect 13725 6879 13783 6885
rect 13924 6888 15108 6916
rect 11054 6857 11060 6860
rect 9815 6820 11008 6848
rect 9815 6817 9827 6820
rect 9769 6811 9827 6817
rect 11048 6811 11060 6857
rect 11112 6848 11118 6860
rect 11112 6820 11148 6848
rect 11054 6808 11060 6811
rect 11112 6808 11118 6820
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 13924 6848 13952 6888
rect 15102 6876 15108 6888
rect 15160 6876 15166 6928
rect 19334 6876 19340 6928
rect 19392 6916 19398 6928
rect 19610 6916 19616 6928
rect 19392 6888 19616 6916
rect 19392 6876 19398 6888
rect 19610 6876 19616 6888
rect 19668 6876 19674 6928
rect 24020 6919 24078 6925
rect 24020 6885 24032 6919
rect 24066 6916 24078 6919
rect 24302 6916 24308 6928
rect 24066 6888 24308 6916
rect 24066 6885 24078 6888
rect 24020 6879 24078 6885
rect 24302 6876 24308 6888
rect 24360 6876 24366 6928
rect 12308 6820 13952 6848
rect 12308 6808 12314 6820
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14274 6848 14280 6860
rect 14056 6820 14280 6848
rect 14056 6808 14062 6820
rect 14274 6808 14280 6820
rect 14332 6848 14338 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 14332 6820 15025 6848
rect 14332 6808 14338 6820
rect 15013 6817 15025 6820
rect 15059 6817 15071 6851
rect 15562 6848 15568 6860
rect 15523 6820 15568 6848
rect 15013 6811 15071 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 16114 6808 16120 6860
rect 16172 6848 16178 6860
rect 16281 6851 16339 6857
rect 16281 6848 16293 6851
rect 16172 6820 16293 6848
rect 16172 6808 16178 6820
rect 16281 6817 16293 6820
rect 16327 6817 16339 6851
rect 16281 6811 16339 6817
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 19981 6851 20039 6857
rect 19981 6848 19993 6851
rect 18196 6820 19993 6848
rect 18196 6808 18202 6820
rect 19981 6817 19993 6820
rect 20027 6848 20039 6851
rect 20070 6848 20076 6860
rect 20027 6820 20076 6848
rect 20027 6817 20039 6820
rect 19981 6811 20039 6817
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 20622 6808 20628 6860
rect 20680 6848 20686 6860
rect 21157 6851 21215 6857
rect 21157 6848 21169 6851
rect 20680 6820 21169 6848
rect 20680 6808 20686 6820
rect 21157 6817 21169 6820
rect 21203 6817 21215 6851
rect 21157 6811 21215 6817
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8036 6752 8493 6780
rect 7929 6715 7987 6721
rect 6972 6684 7880 6712
rect 6972 6672 6978 6684
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 1728 6616 3433 6644
rect 1728 6604 1734 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 3881 6647 3939 6653
rect 3881 6613 3893 6647
rect 3927 6644 3939 6647
rect 4614 6644 4620 6656
rect 3927 6616 4620 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 4614 6604 4620 6616
rect 4672 6644 4678 6656
rect 5074 6644 5080 6656
rect 4672 6616 5080 6644
rect 4672 6604 4678 6616
rect 5074 6604 5080 6616
rect 5132 6644 5138 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 5132 6616 6837 6644
rect 5132 6604 5138 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 7650 6644 7656 6656
rect 7611 6616 7656 6644
rect 6825 6607 6883 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 7852 6644 7880 6684
rect 7929 6681 7941 6715
rect 7975 6681 7987 6715
rect 7929 6675 7987 6681
rect 8036 6644 8064 6752
rect 8481 6749 8493 6752
rect 8527 6780 8539 6783
rect 9490 6780 9496 6792
rect 8527 6752 9496 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6749 10839 6783
rect 10781 6743 10839 6749
rect 8938 6644 8944 6656
rect 7852 6616 8064 6644
rect 8899 6616 8944 6644
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9306 6644 9312 6656
rect 9180 6616 9312 6644
rect 9180 6604 9186 6616
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 9732 6616 10241 6644
rect 9732 6604 9738 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10594 6644 10600 6656
rect 10555 6616 10600 6644
rect 10229 6607 10287 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10796 6644 10824 6743
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 13412 6752 13829 6780
rect 13412 6740 13418 6752
rect 13817 6749 13829 6752
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 12897 6715 12955 6721
rect 12897 6681 12909 6715
rect 12943 6712 12955 6715
rect 13924 6712 13952 6743
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 16025 6783 16083 6789
rect 16025 6780 16037 6783
rect 15896 6752 16037 6780
rect 15896 6740 15902 6752
rect 16025 6749 16037 6752
rect 16071 6749 16083 6783
rect 18966 6780 18972 6792
rect 18927 6752 18972 6780
rect 16025 6743 16083 6749
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19116 6752 19161 6780
rect 19116 6740 19122 6752
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20864 6752 20913 6780
rect 20864 6740 20870 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 23753 6783 23811 6789
rect 23753 6780 23765 6783
rect 23624 6752 23765 6780
rect 23624 6740 23630 6752
rect 23753 6749 23765 6752
rect 23799 6749 23811 6783
rect 23753 6743 23811 6749
rect 13998 6712 14004 6724
rect 12943 6684 14004 6712
rect 12943 6681 12955 6684
rect 12897 6675 12955 6681
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 11146 6644 11152 6656
rect 10796 6616 11152 6644
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 13357 6647 13415 6653
rect 13357 6613 13369 6647
rect 13403 6644 13415 6647
rect 13722 6644 13728 6656
rect 13403 6616 13728 6644
rect 13403 6613 13415 6616
rect 13357 6607 13415 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14369 6647 14427 6653
rect 14369 6644 14381 6647
rect 14148 6616 14381 6644
rect 14148 6604 14154 6616
rect 14369 6613 14381 6616
rect 14415 6613 14427 6647
rect 14369 6607 14427 6613
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 16206 6644 16212 6656
rect 15979 6616 16212 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18509 6647 18567 6653
rect 18509 6644 18521 6647
rect 18012 6616 18521 6644
rect 18012 6604 18018 6616
rect 18509 6613 18521 6616
rect 18555 6613 18567 6647
rect 19518 6644 19524 6656
rect 19479 6616 19524 6644
rect 18509 6607 18567 6613
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 22922 6644 22928 6656
rect 22883 6616 22928 6644
rect 22922 6604 22928 6616
rect 22980 6604 22986 6656
rect 23661 6647 23719 6653
rect 23661 6613 23673 6647
rect 23707 6644 23719 6647
rect 25130 6644 25136 6656
rect 23707 6616 25136 6644
rect 23707 6613 23719 6616
rect 23661 6607 23719 6613
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2130 6440 2136 6452
rect 2091 6412 2136 6440
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 2832 6412 2877 6440
rect 2832 6400 2838 6412
rect 3142 6400 3148 6452
rect 3200 6440 3206 6452
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 3200 6412 4445 6440
rect 3200 6400 3206 6412
rect 4433 6409 4445 6412
rect 4479 6409 4491 6443
rect 4433 6403 4491 6409
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5592 6412 5825 6440
rect 5592 6400 5598 6412
rect 5813 6409 5825 6412
rect 5859 6409 5871 6443
rect 5813 6403 5871 6409
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6914 6440 6920 6452
rect 6687 6412 6920 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 9490 6440 9496 6452
rect 9451 6412 9496 6440
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 12986 6440 12992 6452
rect 10744 6412 12992 6440
rect 10744 6400 10750 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13354 6440 13360 6452
rect 13315 6412 13360 6440
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 14700 6412 15117 6440
rect 14700 6400 14706 6412
rect 15105 6409 15117 6412
rect 15151 6409 15163 6443
rect 15105 6403 15163 6409
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17497 6443 17555 6449
rect 17497 6440 17509 6443
rect 17460 6412 17509 6440
rect 17460 6400 17466 6412
rect 17497 6409 17509 6412
rect 17543 6440 17555 6443
rect 17865 6443 17923 6449
rect 17865 6440 17877 6443
rect 17543 6412 17877 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17865 6409 17877 6412
rect 17911 6440 17923 6443
rect 19058 6440 19064 6452
rect 17911 6412 19064 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 20806 6440 20812 6452
rect 19260 6412 20812 6440
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6372 2559 6375
rect 2866 6372 2872 6384
rect 2547 6344 2872 6372
rect 2547 6341 2559 6344
rect 2501 6335 2559 6341
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 5442 6372 5448 6384
rect 4212 6344 5448 6372
rect 4212 6332 4218 6344
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 10502 6372 10508 6384
rect 10415 6344 10508 6372
rect 10502 6332 10508 6344
rect 10560 6372 10566 6384
rect 11330 6372 11336 6384
rect 10560 6344 11336 6372
rect 10560 6332 10566 6344
rect 11330 6332 11336 6344
rect 11388 6332 11394 6384
rect 11606 6332 11612 6384
rect 11664 6372 11670 6384
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 11664 6344 12173 6372
rect 11664 6332 11670 6344
rect 12161 6341 12173 6344
rect 12207 6341 12219 6375
rect 12161 6335 12219 6341
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3326 6304 3332 6316
rect 3283 6276 3332 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3510 6304 3516 6316
rect 3467 6276 3516 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 5074 6304 5080 6316
rect 5035 6276 5080 6304
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6236 6276 6837 6304
rect 6236 6264 6242 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 11149 6307 11207 6313
rect 11149 6304 11161 6307
rect 10192 6276 11161 6304
rect 10192 6264 10198 6276
rect 11149 6273 11161 6276
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 3142 6236 3148 6248
rect 3103 6208 3148 6236
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 4019 6208 4813 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4801 6205 4813 6208
rect 4847 6236 4859 6239
rect 7466 6236 7472 6248
rect 4847 6208 7472 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7883 6208 8125 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 8202 6236 8208 6248
rect 8159 6208 8208 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10744 6208 10977 6236
rect 10744 6196 10750 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 12176 6236 12204 6335
rect 17034 6304 17040 6316
rect 16947 6276 17040 6304
rect 17034 6264 17040 6276
rect 17092 6304 17098 6316
rect 17420 6304 17448 6400
rect 18785 6375 18843 6381
rect 18785 6341 18797 6375
rect 18831 6372 18843 6375
rect 18966 6372 18972 6384
rect 18831 6344 18972 6372
rect 18831 6341 18843 6344
rect 18785 6335 18843 6341
rect 18966 6332 18972 6344
rect 19024 6332 19030 6384
rect 17092 6276 17448 6304
rect 17092 6264 17098 6276
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12176 6208 12633 6236
rect 10965 6199 11023 6205
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 13998 6245 14004 6248
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 12860 6208 13737 6236
rect 12860 6196 12866 6208
rect 13725 6205 13737 6208
rect 13771 6205 13783 6239
rect 13992 6236 14004 6245
rect 13959 6208 14004 6236
rect 13725 6199 13783 6205
rect 13992 6199 14004 6208
rect 8386 6177 8392 6180
rect 4341 6171 4399 6177
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 7653 6171 7711 6177
rect 4387 6140 4936 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 4908 6112 4936 6140
rect 7653 6137 7665 6171
rect 7699 6168 7711 6171
rect 8380 6168 8392 6177
rect 7699 6140 8392 6168
rect 7699 6137 7711 6140
rect 7653 6131 7711 6137
rect 8380 6131 8392 6140
rect 8386 6128 8392 6131
rect 8444 6128 8450 6180
rect 11057 6171 11115 6177
rect 11057 6137 11069 6171
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 1397 6103 1455 6109
rect 1397 6069 1409 6103
rect 1443 6100 1455 6103
rect 1578 6100 1584 6112
rect 1443 6072 1584 6100
rect 1443 6069 1455 6072
rect 1397 6063 1455 6069
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 6178 6100 6184 6112
rect 4948 6072 4993 6100
rect 6139 6072 6184 6100
rect 4948 6060 4954 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7616 6072 7849 6100
rect 7616 6060 7622 6072
rect 7837 6069 7849 6072
rect 7883 6100 7895 6103
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7883 6072 7941 6100
rect 7883 6069 7895 6072
rect 7837 6063 7895 6069
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 10134 6100 10140 6112
rect 10095 6072 10140 6100
rect 7929 6063 7987 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 10870 6100 10876 6112
rect 10643 6072 10876 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11072 6100 11100 6131
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 11609 6171 11667 6177
rect 11609 6168 11621 6171
rect 11204 6140 11621 6168
rect 11204 6128 11210 6140
rect 11609 6137 11621 6140
rect 11655 6137 11667 6171
rect 13740 6168 13768 6199
rect 13998 6196 14004 6199
rect 14056 6196 14062 6248
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 16853 6239 16911 6245
rect 16853 6236 16865 6239
rect 16632 6208 16865 6236
rect 16632 6196 16638 6208
rect 16853 6205 16865 6208
rect 16899 6236 16911 6239
rect 17678 6236 17684 6248
rect 16899 6208 17684 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 18138 6236 18144 6248
rect 18099 6208 18144 6236
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 19260 6245 19288 6412
rect 20806 6400 20812 6412
rect 20864 6440 20870 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20864 6412 21189 6440
rect 20864 6400 20870 6412
rect 21177 6409 21189 6412
rect 21223 6440 21235 6443
rect 22278 6440 22284 6452
rect 21223 6412 22284 6440
rect 21223 6409 21235 6412
rect 21177 6403 21235 6409
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 22649 6307 22707 6313
rect 22649 6273 22661 6307
rect 22695 6304 22707 6307
rect 22922 6304 22928 6316
rect 22695 6276 22928 6304
rect 22695 6273 22707 6276
rect 22649 6267 22707 6273
rect 22922 6264 22928 6276
rect 22980 6304 22986 6316
rect 23382 6304 23388 6316
rect 22980 6276 23388 6304
rect 22980 6264 22986 6276
rect 23382 6264 23388 6276
rect 23440 6264 23446 6316
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 14090 6168 14096 6180
rect 13740 6140 14096 6168
rect 11609 6131 11667 6137
rect 14090 6128 14096 6140
rect 14148 6168 14154 6180
rect 15838 6168 15844 6180
rect 14148 6140 15844 6168
rect 14148 6128 14154 6140
rect 15838 6128 15844 6140
rect 15896 6128 15902 6180
rect 16298 6168 16304 6180
rect 16211 6140 16304 6168
rect 16298 6128 16304 6140
rect 16356 6168 16362 6180
rect 16761 6171 16819 6177
rect 16761 6168 16773 6171
rect 16356 6140 16773 6168
rect 16356 6128 16362 6140
rect 16761 6137 16773 6140
rect 16807 6168 16819 6171
rect 17494 6168 17500 6180
rect 16807 6140 17500 6168
rect 16807 6137 16819 6140
rect 16761 6131 16819 6137
rect 17494 6128 17500 6140
rect 17552 6128 17558 6180
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 19061 6171 19119 6177
rect 19061 6168 19073 6171
rect 17828 6140 19073 6168
rect 17828 6128 17834 6140
rect 19061 6137 19073 6140
rect 19107 6168 19119 6171
rect 19260 6168 19288 6199
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 19392 6208 19656 6236
rect 19392 6196 19398 6208
rect 19628 6180 19656 6208
rect 22278 6196 22284 6248
rect 22336 6236 22342 6248
rect 23477 6239 23535 6245
rect 23477 6236 23489 6239
rect 22336 6208 23489 6236
rect 22336 6196 22342 6208
rect 23477 6205 23489 6208
rect 23523 6236 23535 6239
rect 23566 6236 23572 6248
rect 23523 6208 23572 6236
rect 23523 6205 23535 6208
rect 23477 6199 23535 6205
rect 23566 6196 23572 6208
rect 23624 6236 23630 6248
rect 23937 6239 23995 6245
rect 23937 6236 23949 6239
rect 23624 6208 23949 6236
rect 23624 6196 23630 6208
rect 23937 6205 23949 6208
rect 23983 6236 23995 6239
rect 24121 6239 24179 6245
rect 24121 6236 24133 6239
rect 23983 6208 24133 6236
rect 23983 6205 23995 6208
rect 23937 6199 23995 6205
rect 24121 6205 24133 6208
rect 24167 6205 24179 6239
rect 24121 6199 24179 6205
rect 24388 6239 24446 6245
rect 24388 6205 24400 6239
rect 24434 6236 24446 6239
rect 24762 6236 24768 6248
rect 24434 6208 24768 6236
rect 24434 6205 24446 6208
rect 24388 6199 24446 6205
rect 24762 6196 24768 6208
rect 24820 6236 24826 6248
rect 25130 6236 25136 6248
rect 24820 6208 25136 6236
rect 24820 6196 24826 6208
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 19518 6177 19524 6180
rect 19512 6168 19524 6177
rect 19107 6140 19288 6168
rect 19479 6140 19524 6168
rect 19107 6137 19119 6140
rect 19061 6131 19119 6137
rect 19512 6131 19524 6140
rect 19518 6128 19524 6131
rect 19576 6128 19582 6180
rect 19610 6128 19616 6180
rect 19668 6128 19674 6180
rect 22373 6171 22431 6177
rect 22373 6168 22385 6171
rect 21836 6140 22385 6168
rect 21836 6112 21864 6140
rect 22373 6137 22385 6140
rect 22419 6137 22431 6171
rect 22373 6131 22431 6137
rect 11330 6100 11336 6112
rect 11072 6072 11336 6100
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 13722 6100 13728 6112
rect 12851 6072 13728 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 16393 6103 16451 6109
rect 16393 6069 16405 6103
rect 16439 6100 16451 6103
rect 16482 6100 16488 6112
rect 16439 6072 16488 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 19242 6100 19248 6112
rect 18371 6072 19248 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19978 6060 19984 6112
rect 20036 6100 20042 6112
rect 20622 6100 20628 6112
rect 20036 6072 20628 6100
rect 20036 6060 20042 6072
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 21818 6100 21824 6112
rect 21779 6072 21824 6100
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 22002 6100 22008 6112
rect 21963 6072 22008 6100
rect 22002 6060 22008 6072
rect 22060 6060 22066 6112
rect 22465 6103 22523 6109
rect 22465 6069 22477 6103
rect 22511 6100 22523 6103
rect 22554 6100 22560 6112
rect 22511 6072 22560 6100
rect 22511 6069 22523 6072
rect 22465 6063 22523 6069
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 25498 6100 25504 6112
rect 25459 6072 25504 6100
rect 25498 6060 25504 6072
rect 25556 6060 25562 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 2777 5899 2835 5905
rect 2777 5896 2789 5899
rect 2740 5868 2789 5896
rect 2740 5856 2746 5868
rect 2777 5865 2789 5868
rect 2823 5865 2835 5899
rect 2777 5859 2835 5865
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 3510 5896 3516 5908
rect 3467 5868 3516 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4488 5868 4537 5896
rect 4488 5856 4494 5868
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 5626 5896 5632 5908
rect 5587 5868 5632 5896
rect 4525 5859 4583 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 6972 5868 7481 5896
rect 6972 5856 6978 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 7469 5859 7527 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8481 5899 8539 5905
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 8846 5896 8852 5908
rect 8527 5868 8852 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 9858 5896 9864 5908
rect 9723 5868 9864 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11054 5896 11060 5908
rect 10919 5868 11060 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11238 5896 11244 5908
rect 11199 5868 11244 5896
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12529 5899 12587 5905
rect 12529 5896 12541 5899
rect 12492 5868 12541 5896
rect 12492 5856 12498 5868
rect 12529 5865 12541 5868
rect 12575 5896 12587 5899
rect 13538 5896 13544 5908
rect 12575 5868 13544 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 13998 5856 14004 5908
rect 14056 5896 14062 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 14056 5868 14105 5896
rect 14056 5856 14062 5868
rect 14093 5865 14105 5868
rect 14139 5896 14151 5899
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14139 5868 14657 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 14826 5856 14832 5908
rect 14884 5896 14890 5908
rect 15013 5899 15071 5905
rect 15013 5896 15025 5899
rect 14884 5868 15025 5896
rect 14884 5856 14890 5868
rect 15013 5865 15025 5868
rect 15059 5865 15071 5899
rect 16114 5896 16120 5908
rect 16075 5868 16120 5896
rect 15013 5859 15071 5865
rect 10134 5828 10140 5840
rect 9876 5800 10140 5828
rect 9876 5772 9904 5800
rect 10134 5788 10140 5800
rect 10192 5788 10198 5840
rect 12980 5831 13038 5837
rect 12980 5797 12992 5831
rect 13026 5828 13038 5831
rect 13170 5828 13176 5840
rect 13026 5800 13176 5828
rect 13026 5797 13038 5800
rect 12980 5791 13038 5797
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2685 5763 2743 5769
rect 2685 5760 2697 5763
rect 2648 5732 2697 5760
rect 2648 5720 2654 5732
rect 2685 5729 2697 5732
rect 2731 5729 2743 5763
rect 2685 5723 2743 5729
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4120 5732 4445 5760
rect 4120 5720 4126 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 5994 5760 6000 5772
rect 5955 5732 6000 5760
rect 4433 5723 4491 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 8478 5760 8484 5772
rect 8435 5732 8484 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 9858 5720 9864 5772
rect 9916 5720 9922 5772
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 10008 5732 10057 5760
rect 10008 5720 10014 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 11204 5732 12725 5760
rect 11204 5720 11210 5732
rect 12713 5729 12725 5732
rect 12759 5760 12771 5763
rect 12802 5760 12808 5772
rect 12759 5732 12808 5760
rect 12759 5729 12771 5732
rect 12713 5723 12771 5729
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 15028 5760 15056 5859
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 16485 5899 16543 5905
rect 16485 5865 16497 5899
rect 16531 5896 16543 5899
rect 16574 5896 16580 5908
rect 16531 5868 16580 5896
rect 16531 5865 16543 5868
rect 16485 5859 16543 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 18785 5899 18843 5905
rect 18785 5865 18797 5899
rect 18831 5896 18843 5899
rect 18874 5896 18880 5908
rect 18831 5868 18880 5896
rect 18831 5865 18843 5868
rect 18785 5859 18843 5865
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 19705 5899 19763 5905
rect 19705 5865 19717 5899
rect 19751 5896 19763 5899
rect 20070 5896 20076 5908
rect 19751 5868 20076 5896
rect 19751 5865 19763 5868
rect 19705 5859 19763 5865
rect 20070 5856 20076 5868
rect 20128 5896 20134 5908
rect 20438 5896 20444 5908
rect 20128 5868 20444 5896
rect 20128 5856 20134 5868
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 20622 5856 20628 5908
rect 20680 5896 20686 5908
rect 21637 5899 21695 5905
rect 21637 5896 21649 5899
rect 20680 5868 21649 5896
rect 20680 5856 20686 5868
rect 21637 5865 21649 5868
rect 21683 5865 21695 5899
rect 21637 5859 21695 5865
rect 24397 5899 24455 5905
rect 24397 5865 24409 5899
rect 24443 5896 24455 5899
rect 24670 5896 24676 5908
rect 24443 5868 24676 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 24946 5856 24952 5908
rect 25004 5896 25010 5908
rect 25041 5899 25099 5905
rect 25041 5896 25053 5899
rect 25004 5868 25053 5896
rect 25004 5856 25010 5868
rect 25041 5865 25053 5868
rect 25087 5865 25099 5899
rect 25041 5859 25099 5865
rect 17034 5837 17040 5840
rect 17028 5828 17040 5837
rect 16995 5800 17040 5828
rect 17028 5791 17040 5800
rect 17034 5788 17040 5791
rect 17092 5788 17098 5840
rect 22097 5831 22155 5837
rect 22097 5797 22109 5831
rect 22143 5828 22155 5831
rect 22554 5828 22560 5840
rect 22143 5800 22560 5828
rect 22143 5797 22155 5800
rect 22097 5791 22155 5797
rect 22554 5788 22560 5800
rect 22612 5828 22618 5840
rect 23474 5828 23480 5840
rect 22612 5800 23480 5828
rect 22612 5788 22618 5800
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 15289 5763 15347 5769
rect 15289 5760 15301 5763
rect 15028 5732 15301 5760
rect 15289 5729 15301 5732
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 16758 5760 16764 5772
rect 15896 5732 16764 5760
rect 15896 5720 15902 5732
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 19610 5760 19616 5772
rect 19571 5732 19616 5760
rect 19610 5720 19616 5732
rect 19668 5720 19674 5772
rect 21085 5763 21143 5769
rect 21085 5729 21097 5763
rect 21131 5760 21143 5763
rect 21726 5760 21732 5772
rect 21131 5732 21732 5760
rect 21131 5729 21143 5732
rect 21085 5723 21143 5729
rect 21726 5720 21732 5732
rect 21784 5720 21790 5772
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5760 22247 5763
rect 22278 5760 22284 5772
rect 22235 5732 22284 5760
rect 22235 5729 22247 5732
rect 22189 5723 22247 5729
rect 22278 5720 22284 5732
rect 22336 5720 22342 5772
rect 22456 5763 22514 5769
rect 22456 5729 22468 5763
rect 22502 5760 22514 5763
rect 22738 5760 22744 5772
rect 22502 5732 22744 5760
rect 22502 5729 22514 5732
rect 22456 5723 22514 5729
rect 22738 5720 22744 5732
rect 22796 5720 22802 5772
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2700 5664 2881 5692
rect 2700 5636 2728 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 2682 5584 2688 5636
rect 2740 5584 2746 5636
rect 3970 5584 3976 5636
rect 4028 5624 4034 5636
rect 4065 5627 4123 5633
rect 4065 5624 4077 5627
rect 4028 5596 4077 5624
rect 4028 5584 4034 5596
rect 4065 5593 4077 5596
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 4724 5568 4752 5655
rect 5258 5652 5264 5704
rect 5316 5692 5322 5704
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 5316 5664 6101 5692
rect 5316 5652 5322 5664
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5661 6239 5695
rect 6181 5655 6239 5661
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5661 8723 5695
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 8665 5655 8723 5661
rect 6196 5624 6224 5655
rect 5092 5596 6224 5624
rect 7929 5627 7987 5633
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2314 5556 2320 5568
rect 2275 5528 2320 5556
rect 2314 5516 2320 5528
rect 2372 5516 2378 5568
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5556 3847 5559
rect 4246 5556 4252 5568
rect 3835 5528 4252 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 5092 5565 5120 5596
rect 7929 5593 7941 5627
rect 7975 5624 7987 5627
rect 8386 5624 8392 5636
rect 7975 5596 8392 5624
rect 7975 5593 7987 5596
rect 7929 5587 7987 5593
rect 8386 5584 8392 5596
rect 8444 5624 8450 5636
rect 8680 5624 8708 5655
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10318 5692 10324 5704
rect 10279 5664 10324 5692
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 11698 5692 11704 5704
rect 11659 5664 11704 5692
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5692 19947 5695
rect 25130 5692 25136 5704
rect 19935 5664 20668 5692
rect 25091 5664 25136 5692
rect 19935 5661 19947 5664
rect 19889 5655 19947 5661
rect 9030 5624 9036 5636
rect 8444 5596 9036 5624
rect 8444 5584 8450 5596
rect 9030 5584 9036 5596
rect 9088 5624 9094 5636
rect 10336 5624 10364 5652
rect 9088 5596 10364 5624
rect 19153 5627 19211 5633
rect 9088 5584 9094 5596
rect 19153 5593 19165 5627
rect 19199 5624 19211 5627
rect 19518 5624 19524 5636
rect 19199 5596 19524 5624
rect 19199 5593 19211 5596
rect 19153 5587 19211 5593
rect 19518 5584 19524 5596
rect 19576 5624 19582 5636
rect 19904 5624 19932 5655
rect 19576 5596 19932 5624
rect 19576 5584 19582 5596
rect 20640 5568 20668 5664
rect 25130 5652 25136 5664
rect 25188 5652 25194 5704
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5692 25375 5695
rect 25498 5692 25504 5704
rect 25363 5664 25504 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 23842 5584 23848 5636
rect 23900 5624 23906 5636
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 23900 5596 24685 5624
rect 23900 5584 23906 5596
rect 24673 5593 24685 5596
rect 24719 5593 24731 5627
rect 24673 5587 24731 5593
rect 24854 5584 24860 5636
rect 24912 5624 24918 5636
rect 25332 5624 25360 5655
rect 25498 5652 25504 5664
rect 25556 5652 25562 5704
rect 24912 5596 25360 5624
rect 24912 5584 24918 5596
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 4764 5528 5089 5556
rect 4764 5516 4770 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5077 5519 5135 5525
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 6914 5556 6920 5568
rect 6875 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 11514 5556 11520 5568
rect 11475 5528 11520 5556
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 15470 5556 15476 5568
rect 15431 5528 15476 5556
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 18138 5556 18144 5568
rect 18099 5528 18144 5556
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 19245 5559 19303 5565
rect 19245 5525 19257 5559
rect 19291 5556 19303 5559
rect 19334 5556 19340 5568
rect 19291 5528 19340 5556
rect 19291 5525 19303 5528
rect 19245 5519 19303 5525
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 20622 5556 20628 5568
rect 20583 5528 20628 5556
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 21266 5556 21272 5568
rect 21227 5528 21272 5556
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 23382 5516 23388 5568
rect 23440 5556 23446 5568
rect 23569 5559 23627 5565
rect 23569 5556 23581 5559
rect 23440 5528 23581 5556
rect 23440 5516 23446 5528
rect 23569 5525 23581 5528
rect 23615 5525 23627 5559
rect 23569 5519 23627 5525
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 1670 5352 1676 5364
rect 1443 5324 1676 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3789 5355 3847 5361
rect 3789 5352 3801 5355
rect 2832 5324 2877 5352
rect 3252 5324 3801 5352
rect 2832 5312 2838 5324
rect 2038 5216 2044 5228
rect 1951 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5216 2102 5228
rect 2682 5216 2688 5228
rect 2096 5188 2688 5216
rect 2096 5176 2102 5188
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 3252 5225 3280 5324
rect 3789 5321 3801 5324
rect 3835 5352 3847 5355
rect 4062 5352 4068 5364
rect 3835 5324 4068 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 4430 5352 4436 5364
rect 4203 5324 4436 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 4430 5312 4436 5324
rect 4488 5312 4494 5364
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 8846 5352 8852 5364
rect 8628 5324 8852 5352
rect 8628 5312 8634 5324
rect 8846 5312 8852 5324
rect 8904 5352 8910 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8904 5324 9137 5352
rect 8904 5312 8910 5324
rect 9125 5321 9137 5324
rect 9171 5321 9183 5355
rect 11330 5352 11336 5364
rect 11291 5324 11336 5352
rect 9125 5315 9183 5321
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 11790 5352 11796 5364
rect 11751 5324 11796 5352
rect 11790 5312 11796 5324
rect 11848 5352 11854 5364
rect 12342 5352 12348 5364
rect 11848 5324 12348 5352
rect 11848 5312 11854 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12860 5324 13001 5352
rect 12860 5312 12866 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 13538 5352 13544 5364
rect 13499 5324 13544 5352
rect 12989 5315 13047 5321
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14148 5324 14933 5352
rect 14148 5312 14154 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 8757 5287 8815 5293
rect 8757 5284 8769 5287
rect 8536 5256 8769 5284
rect 8536 5244 8542 5256
rect 8757 5253 8769 5256
rect 8803 5253 8815 5287
rect 8757 5247 8815 5253
rect 10689 5287 10747 5293
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 10735 5256 12173 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 12161 5253 12173 5256
rect 12207 5284 12219 5287
rect 13170 5284 13176 5296
rect 12207 5256 13176 5284
rect 12207 5253 12219 5256
rect 12161 5247 12219 5253
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 5316 5188 6193 5216
rect 5316 5176 5322 5188
rect 6181 5185 6193 5188
rect 6227 5216 6239 5219
rect 6638 5216 6644 5228
rect 6227 5188 6644 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 8772 5216 8800 5247
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 13449 5219 13507 5225
rect 8772 5188 9444 5216
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1636 5120 1777 5148
rect 1636 5108 1642 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 4249 5151 4307 5157
rect 4249 5148 4261 5151
rect 4212 5120 4261 5148
rect 4212 5108 4218 5120
rect 4249 5117 4261 5120
rect 4295 5148 4307 5151
rect 6454 5148 6460 5160
rect 4295 5120 6460 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 6454 5108 6460 5120
rect 6512 5148 6518 5160
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 6512 5120 6561 5148
rect 6512 5108 6518 5120
rect 6549 5117 6561 5120
rect 6595 5148 6607 5151
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6595 5120 6837 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7081 5151 7139 5157
rect 7081 5148 7093 5151
rect 6972 5120 7093 5148
rect 6972 5108 6978 5120
rect 7081 5117 7093 5120
rect 7127 5117 7139 5151
rect 7081 5111 7139 5117
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 8996 5120 9321 5148
rect 8996 5108 9002 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9416 5148 9444 5188
rect 13449 5185 13461 5219
rect 13495 5216 13507 5219
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13495 5188 14197 5216
rect 13495 5185 13507 5188
rect 13449 5179 13507 5185
rect 14185 5185 14197 5188
rect 14231 5216 14243 5219
rect 14642 5216 14648 5228
rect 14231 5188 14648 5216
rect 14231 5185 14243 5188
rect 14185 5179 14243 5185
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 14936 5216 14964 5315
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 16816 5324 17049 5352
rect 16816 5312 16822 5324
rect 17037 5321 17049 5324
rect 17083 5352 17095 5355
rect 17770 5352 17776 5364
rect 17083 5324 17776 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17770 5312 17776 5324
rect 17828 5352 17834 5364
rect 20070 5352 20076 5364
rect 17828 5324 18092 5352
rect 20031 5324 20076 5352
rect 17828 5312 17834 5324
rect 16482 5284 16488 5296
rect 16443 5256 16488 5284
rect 16482 5244 16488 5256
rect 16540 5244 16546 5296
rect 18064 5225 18092 5324
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 21637 5355 21695 5361
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 21726 5352 21732 5364
rect 21683 5324 21732 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 24305 5355 24363 5361
rect 24305 5321 24317 5355
rect 24351 5352 24363 5355
rect 25130 5352 25136 5364
rect 24351 5324 25136 5352
rect 24351 5321 24363 5324
rect 24305 5315 24363 5321
rect 25130 5312 25136 5324
rect 25188 5352 25194 5364
rect 25685 5355 25743 5361
rect 25685 5352 25697 5355
rect 25188 5324 25697 5352
rect 25188 5312 25194 5324
rect 25685 5321 25697 5324
rect 25731 5321 25743 5355
rect 25685 5315 25743 5321
rect 19429 5287 19487 5293
rect 19429 5253 19441 5287
rect 19475 5253 19487 5287
rect 19429 5247 19487 5253
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 14936 5188 15117 5216
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5185 18107 5219
rect 19444 5216 19472 5247
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 24029 5287 24087 5293
rect 24029 5284 24041 5287
rect 19576 5256 24041 5284
rect 19576 5244 19582 5256
rect 24029 5253 24041 5256
rect 24075 5284 24087 5287
rect 24121 5287 24179 5293
rect 24121 5284 24133 5287
rect 24075 5256 24133 5284
rect 24075 5253 24087 5256
rect 24029 5247 24087 5253
rect 24121 5253 24133 5256
rect 24167 5253 24179 5287
rect 24121 5247 24179 5253
rect 24946 5244 24952 5296
rect 25004 5284 25010 5296
rect 25317 5287 25375 5293
rect 25317 5284 25329 5287
rect 25004 5256 25329 5284
rect 25004 5244 25010 5256
rect 25317 5253 25329 5256
rect 25363 5253 25375 5287
rect 25317 5247 25375 5253
rect 20622 5216 20628 5228
rect 19444 5188 20628 5216
rect 18049 5179 18107 5185
rect 20622 5176 20628 5188
rect 20680 5216 20686 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 20680 5188 21097 5216
rect 20680 5176 20686 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 23477 5219 23535 5225
rect 23477 5185 23489 5219
rect 23523 5216 23535 5219
rect 24762 5216 24768 5228
rect 23523 5188 24768 5216
rect 23523 5185 23535 5188
rect 23477 5179 23535 5185
rect 24762 5176 24768 5188
rect 24820 5216 24826 5228
rect 24857 5219 24915 5225
rect 24857 5216 24869 5219
rect 24820 5188 24869 5216
rect 24820 5176 24826 5188
rect 24857 5185 24869 5188
rect 24903 5185 24915 5219
rect 24857 5179 24915 5185
rect 10778 5148 10784 5160
rect 9416 5120 10784 5148
rect 9309 5111 9367 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12492 5120 12537 5148
rect 12492 5108 12498 5120
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 13909 5151 13967 5157
rect 13909 5148 13921 5151
rect 13872 5120 13921 5148
rect 13872 5108 13878 5120
rect 13909 5117 13921 5120
rect 13955 5117 13967 5151
rect 13909 5111 13967 5117
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14734 5148 14740 5160
rect 14047 5120 14740 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 4516 5083 4574 5089
rect 4516 5049 4528 5083
rect 4562 5080 4574 5083
rect 4706 5080 4712 5092
rect 4562 5052 4712 5080
rect 4562 5049 4574 5052
rect 4516 5043 4574 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 6932 5080 6960 5108
rect 9398 5080 9404 5092
rect 5644 5052 6960 5080
rect 8220 5052 9404 5080
rect 1486 4972 1492 5024
rect 1544 5012 1550 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1544 4984 1869 5012
rect 1544 4972 1550 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 2409 5015 2467 5021
rect 2409 5012 2421 5015
rect 2096 4984 2421 5012
rect 2096 4972 2102 4984
rect 2409 4981 2421 4984
rect 2455 5012 2467 5015
rect 2590 5012 2596 5024
rect 2455 4984 2596 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 5644 5021 5672 5052
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 5500 4984 5641 5012
rect 5500 4972 5506 4984
rect 5629 4981 5641 4984
rect 5675 4981 5687 5015
rect 5629 4975 5687 4981
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 8220 5021 8248 5052
rect 9398 5040 9404 5052
rect 9456 5080 9462 5092
rect 9554 5083 9612 5089
rect 9554 5080 9566 5083
rect 9456 5052 9566 5080
rect 9456 5040 9462 5052
rect 9554 5049 9566 5052
rect 9600 5049 9612 5083
rect 9554 5043 9612 5049
rect 12526 5040 12532 5092
rect 12584 5080 12590 5092
rect 12894 5080 12900 5092
rect 12584 5052 12900 5080
rect 12584 5040 12590 5052
rect 12894 5040 12900 5052
rect 12952 5040 12958 5092
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 14016 5080 14044 5111
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 18138 5108 18144 5160
rect 18196 5148 18202 5160
rect 18305 5151 18363 5157
rect 18305 5148 18317 5151
rect 18196 5120 18317 5148
rect 18196 5108 18202 5120
rect 18305 5117 18317 5120
rect 18351 5117 18363 5151
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 18305 5111 18363 5117
rect 20364 5120 20913 5148
rect 13688 5052 14044 5080
rect 14645 5083 14703 5089
rect 13688 5040 13694 5052
rect 14645 5049 14657 5083
rect 14691 5080 14703 5083
rect 15350 5083 15408 5089
rect 15350 5080 15362 5083
rect 14691 5052 15362 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 15350 5049 15362 5052
rect 15396 5080 15408 5083
rect 15838 5080 15844 5092
rect 15396 5052 15844 5080
rect 15396 5049 15408 5052
rect 15350 5043 15408 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 17494 5080 17500 5092
rect 17407 5052 17500 5080
rect 17494 5040 17500 5052
rect 17552 5080 17558 5092
rect 18156 5080 18184 5108
rect 17552 5052 18184 5080
rect 17552 5040 17558 5052
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 6972 4984 8217 5012
rect 6972 4972 6978 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 8205 4975 8263 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 20254 4972 20260 5024
rect 20312 5012 20318 5024
rect 20364 5021 20392 5120
rect 20901 5117 20913 5120
rect 20947 5148 20959 5151
rect 21818 5148 21824 5160
rect 20947 5120 21824 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 22462 5148 22468 5160
rect 22423 5120 22468 5148
rect 22462 5108 22468 5120
rect 22520 5108 22526 5160
rect 24029 5151 24087 5157
rect 24029 5117 24041 5151
rect 24075 5148 24087 5151
rect 24673 5151 24731 5157
rect 24673 5148 24685 5151
rect 24075 5120 24685 5148
rect 24075 5117 24087 5120
rect 24029 5111 24087 5117
rect 24673 5117 24685 5120
rect 24719 5117 24731 5151
rect 24673 5111 24731 5117
rect 20806 5040 20812 5092
rect 20864 5080 20870 5092
rect 20993 5083 21051 5089
rect 20993 5080 21005 5083
rect 20864 5052 21005 5080
rect 20864 5040 20870 5052
rect 20993 5049 21005 5052
rect 21039 5049 21051 5083
rect 20993 5043 21051 5049
rect 22738 5040 22744 5092
rect 22796 5080 22802 5092
rect 23109 5083 23167 5089
rect 23109 5080 23121 5083
rect 22796 5052 23121 5080
rect 22796 5040 22802 5052
rect 23109 5049 23121 5052
rect 23155 5080 23167 5083
rect 24854 5080 24860 5092
rect 23155 5052 24860 5080
rect 23155 5049 23167 5052
rect 23109 5043 23167 5049
rect 24854 5040 24860 5052
rect 24912 5040 24918 5092
rect 20349 5015 20407 5021
rect 20349 5012 20361 5015
rect 20312 4984 20361 5012
rect 20312 4972 20318 4984
rect 20349 4981 20361 4984
rect 20395 4981 20407 5015
rect 20530 5012 20536 5024
rect 20491 4984 20536 5012
rect 20349 4975 20407 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 22278 5012 22284 5024
rect 22239 4984 22284 5012
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 22649 5015 22707 5021
rect 22649 4981 22661 5015
rect 22695 5012 22707 5015
rect 23198 5012 23204 5024
rect 22695 4984 23204 5012
rect 22695 4981 22707 4984
rect 22649 4975 22707 4981
rect 23198 4972 23204 4984
rect 23256 4972 23262 5024
rect 24670 4972 24676 5024
rect 24728 5012 24734 5024
rect 24765 5015 24823 5021
rect 24765 5012 24777 5015
rect 24728 4984 24777 5012
rect 24728 4972 24734 4984
rect 24765 4981 24777 4984
rect 24811 4981 24823 5015
rect 24765 4975 24823 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1486 4768 1492 4820
rect 1544 4808 1550 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1544 4780 1593 4808
rect 1544 4768 1550 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1581 4771 1639 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 2409 4811 2467 4817
rect 2409 4808 2421 4811
rect 2372 4780 2421 4808
rect 2372 4768 2378 4780
rect 2409 4777 2421 4780
rect 2455 4808 2467 4811
rect 3697 4811 3755 4817
rect 3697 4808 3709 4811
rect 2455 4780 3709 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 3697 4777 3709 4780
rect 3743 4777 3755 4811
rect 3697 4771 3755 4777
rect 4801 4811 4859 4817
rect 4801 4777 4813 4811
rect 4847 4777 4859 4811
rect 5166 4808 5172 4820
rect 5127 4780 5172 4808
rect 4801 4771 4859 4777
rect 4816 4740 4844 4771
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6730 4768 6736 4820
rect 6788 4808 6794 4820
rect 6825 4811 6883 4817
rect 6825 4808 6837 4811
rect 6788 4780 6837 4808
rect 6788 4768 6794 4780
rect 6825 4777 6837 4780
rect 6871 4777 6883 4811
rect 6825 4771 6883 4777
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8352 4780 8401 4808
rect 8352 4768 8358 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 9030 4808 9036 4820
rect 8991 4780 9036 4808
rect 8389 4771 8447 4777
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 9950 4808 9956 4820
rect 9911 4780 9956 4808
rect 9950 4768 9956 4780
rect 10008 4808 10014 4820
rect 12529 4811 12587 4817
rect 10008 4780 12480 4808
rect 10008 4768 10014 4780
rect 11238 4740 11244 4752
rect 4816 4712 6684 4740
rect 6656 4684 6684 4712
rect 10060 4712 11244 4740
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4672 2375 4675
rect 4246 4672 4252 4684
rect 2363 4644 4252 4672
rect 2363 4641 2375 4644
rect 2317 4635 2375 4641
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6696 4644 6745 4672
rect 6696 4632 6702 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 6733 4635 6791 4641
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 8297 4675 8355 4681
rect 8297 4672 8309 4675
rect 8260 4644 8309 4672
rect 8260 4632 8266 4644
rect 8297 4641 8309 4644
rect 8343 4672 8355 4675
rect 9122 4672 9128 4684
rect 8343 4644 9128 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 10060 4681 10088 4712
rect 11238 4700 11244 4712
rect 11296 4700 11302 4752
rect 11416 4743 11474 4749
rect 11416 4709 11428 4743
rect 11462 4740 11474 4743
rect 11606 4740 11612 4752
rect 11462 4712 11612 4740
rect 11462 4709 11474 4712
rect 11416 4703 11474 4709
rect 11606 4700 11612 4712
rect 11664 4740 11670 4752
rect 12158 4740 12164 4752
rect 11664 4712 12164 4740
rect 11664 4700 11670 4712
rect 12158 4700 12164 4712
rect 12216 4700 12222 4752
rect 12452 4740 12480 4780
rect 12529 4777 12541 4811
rect 12575 4808 12587 4811
rect 12710 4808 12716 4820
rect 12575 4780 12716 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 13998 4808 14004 4820
rect 13587 4780 14004 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14550 4768 14556 4820
rect 14608 4808 14614 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 14608 4780 15301 4808
rect 14608 4768 14614 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 16853 4811 16911 4817
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 17126 4808 17132 4820
rect 16899 4780 17132 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 17862 4808 17868 4820
rect 17276 4780 17868 4808
rect 17276 4768 17282 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 19058 4808 19064 4820
rect 19019 4780 19064 4808
rect 19058 4768 19064 4780
rect 19116 4768 19122 4820
rect 19150 4768 19156 4820
rect 19208 4808 19214 4820
rect 19245 4811 19303 4817
rect 19245 4808 19257 4811
rect 19208 4780 19257 4808
rect 19208 4768 19214 4780
rect 19245 4777 19257 4780
rect 19291 4777 19303 4811
rect 19245 4771 19303 4777
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19613 4811 19671 4817
rect 19613 4808 19625 4811
rect 19392 4780 19625 4808
rect 19392 4768 19398 4780
rect 19613 4777 19625 4780
rect 19659 4777 19671 4811
rect 19613 4771 19671 4777
rect 19705 4811 19763 4817
rect 19705 4777 19717 4811
rect 19751 4808 19763 4811
rect 20530 4808 20536 4820
rect 19751 4780 20536 4808
rect 19751 4777 19763 4780
rect 19705 4771 19763 4777
rect 12618 4740 12624 4752
rect 12452 4712 12624 4740
rect 12618 4700 12624 4712
rect 12676 4740 12682 4752
rect 13814 4740 13820 4752
rect 12676 4712 13820 4740
rect 12676 4700 12682 4712
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 14016 4740 14044 4768
rect 14016 4712 14136 4740
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4641 10103 4675
rect 11146 4672 11152 4684
rect 11107 4644 11152 4672
rect 10045 4635 10103 4641
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 14001 4675 14059 4681
rect 14001 4672 14013 4675
rect 13964 4644 14013 4672
rect 13964 4632 13970 4644
rect 14001 4641 14013 4644
rect 14047 4641 14059 4675
rect 14108 4672 14136 4712
rect 16574 4700 16580 4752
rect 16632 4740 16638 4752
rect 17313 4743 17371 4749
rect 17313 4740 17325 4743
rect 16632 4712 17325 4740
rect 16632 4700 16638 4712
rect 17313 4709 17325 4712
rect 17359 4740 17371 4743
rect 17402 4740 17408 4752
rect 17359 4712 17408 4740
rect 17359 4709 17371 4712
rect 17313 4703 17371 4709
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 19518 4700 19524 4752
rect 19576 4740 19582 4752
rect 19720 4740 19748 4771
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 21453 4811 21511 4817
rect 21453 4777 21465 4811
rect 21499 4808 21511 4811
rect 22002 4808 22008 4820
rect 21499 4780 22008 4808
rect 21499 4777 21511 4780
rect 21453 4771 21511 4777
rect 22002 4768 22008 4780
rect 22060 4768 22066 4820
rect 22462 4808 22468 4820
rect 22423 4780 22468 4808
rect 22462 4768 22468 4780
rect 22520 4768 22526 4820
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 19576 4712 19748 4740
rect 21361 4743 21419 4749
rect 19576 4700 19582 4712
rect 21361 4709 21373 4743
rect 21407 4740 21419 4743
rect 21634 4740 21640 4752
rect 21407 4712 21640 4740
rect 21407 4709 21419 4712
rect 21361 4703 21419 4709
rect 21634 4700 21640 4712
rect 21692 4700 21698 4752
rect 14826 4672 14832 4684
rect 14108 4644 14228 4672
rect 14001 4635 14059 4641
rect 2590 4604 2596 4616
rect 2503 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4604 2654 4616
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 2648 4576 3341 4604
rect 2648 4564 2654 4576
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 5442 4604 5448 4616
rect 5403 4576 5448 4604
rect 3329 4567 3387 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 8478 4604 8484 4616
rect 6972 4576 7017 4604
rect 8439 4576 8484 4604
rect 6972 4564 6978 4576
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 14200 4613 14228 4644
rect 14292 4644 14832 4672
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13136 4576 14105 4604
rect 13136 4564 13142 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 4706 4536 4712 4548
rect 4619 4508 4712 4536
rect 4706 4496 4712 4508
rect 4764 4536 4770 4548
rect 4764 4508 6316 4536
rect 4764 4496 4770 4508
rect 6288 4480 6316 4508
rect 6454 4496 6460 4548
rect 6512 4536 6518 4548
rect 7558 4536 7564 4548
rect 6512 4508 7564 4536
rect 6512 4496 6518 4508
rect 7558 4496 7564 4508
rect 7616 4536 7622 4548
rect 7653 4539 7711 4545
rect 7653 4536 7665 4539
rect 7616 4508 7665 4536
rect 7616 4496 7622 4508
rect 7653 4505 7665 4508
rect 7699 4536 7711 4539
rect 8938 4536 8944 4548
rect 7699 4508 8944 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 8938 4496 8944 4508
rect 8996 4536 9002 4548
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 8996 4508 9321 4536
rect 8996 4496 9002 4508
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 9309 4499 9367 4505
rect 10229 4539 10287 4545
rect 10229 4505 10241 4539
rect 10275 4536 10287 4539
rect 10962 4536 10968 4548
rect 10275 4508 10968 4536
rect 10275 4505 10287 4508
rect 10229 4499 10287 4505
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 13630 4536 13636 4548
rect 13591 4508 13636 4536
rect 13630 4496 13636 4508
rect 13688 4496 13694 4548
rect 13814 4496 13820 4548
rect 13872 4536 13878 4548
rect 14292 4536 14320 4644
rect 14826 4632 14832 4644
rect 14884 4672 14890 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 14884 4644 15669 4672
rect 14884 4632 14890 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16761 4675 16819 4681
rect 16761 4641 16773 4675
rect 16807 4672 16819 4675
rect 17034 4672 17040 4684
rect 16807 4644 17040 4672
rect 16807 4641 16819 4644
rect 16761 4635 16819 4641
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 19426 4632 19432 4684
rect 19484 4672 19490 4684
rect 20533 4675 20591 4681
rect 20533 4672 20545 4675
rect 19484 4644 20545 4672
rect 19484 4632 19490 4644
rect 20533 4641 20545 4644
rect 20579 4672 20591 4675
rect 20806 4672 20812 4684
rect 20579 4644 20812 4672
rect 20579 4641 20591 4644
rect 20533 4635 20591 4641
rect 20806 4632 20812 4644
rect 20864 4632 20870 4684
rect 22824 4675 22882 4681
rect 22824 4641 22836 4675
rect 22870 4672 22882 4675
rect 23382 4672 23388 4684
rect 22870 4644 23388 4672
rect 22870 4641 22882 4644
rect 22824 4635 22882 4641
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 25038 4672 25044 4684
rect 24999 4644 25044 4672
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4573 15807 4607
rect 15930 4604 15936 4616
rect 15843 4576 15936 4604
rect 15749 4567 15807 4573
rect 15010 4536 15016 4548
rect 13872 4508 14320 4536
rect 14971 4508 15016 4536
rect 13872 4496 13878 4508
rect 15010 4496 15016 4508
rect 15068 4536 15074 4548
rect 15764 4536 15792 4567
rect 15930 4564 15936 4576
rect 15988 4604 15994 4616
rect 16301 4607 16359 4613
rect 16301 4604 16313 4607
rect 15988 4576 16313 4604
rect 15988 4564 15994 4576
rect 16301 4573 16313 4576
rect 16347 4573 16359 4607
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 16301 4567 16359 4573
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 19794 4604 19800 4616
rect 19755 4576 19800 4604
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 21637 4607 21695 4613
rect 21637 4573 21649 4607
rect 21683 4604 21695 4607
rect 22094 4604 22100 4616
rect 21683 4576 22100 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 22094 4564 22100 4576
rect 22152 4564 22158 4616
rect 22278 4564 22284 4616
rect 22336 4604 22342 4616
rect 22557 4607 22615 4613
rect 22557 4604 22569 4607
rect 22336 4576 22569 4604
rect 22336 4564 22342 4576
rect 22557 4573 22569 4576
rect 22603 4573 22615 4607
rect 22557 4567 22615 4573
rect 15068 4508 15792 4536
rect 18325 4539 18383 4545
rect 15068 4496 15074 4508
rect 18325 4505 18337 4539
rect 18371 4536 18383 4539
rect 18966 4536 18972 4548
rect 18371 4508 18972 4536
rect 18371 4505 18383 4508
rect 18325 4499 18383 4505
rect 18966 4496 18972 4508
rect 19024 4496 19030 4548
rect 20993 4539 21051 4545
rect 20993 4505 21005 4539
rect 21039 4536 21051 4539
rect 21542 4536 21548 4548
rect 21039 4508 21548 4536
rect 21039 4505 21051 4508
rect 20993 4499 21051 4505
rect 21542 4496 21548 4508
rect 21600 4496 21606 4548
rect 2682 4428 2688 4480
rect 2740 4468 2746 4480
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 2740 4440 2973 4468
rect 2740 4428 2746 4440
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 2961 4431 3019 4437
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 4212 4440 4261 4468
rect 4212 4428 4218 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 5813 4471 5871 4477
rect 5813 4468 5825 4471
rect 5408 4440 5825 4468
rect 5408 4428 5414 4440
rect 5813 4437 5825 4440
rect 5859 4468 5871 4471
rect 5994 4468 6000 4480
rect 5859 4440 6000 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6270 4468 6276 4480
rect 6231 4440 6276 4468
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 7926 4468 7932 4480
rect 7887 4440 7932 4468
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 10689 4471 10747 4477
rect 10689 4437 10701 4471
rect 10735 4468 10747 4471
rect 10778 4468 10784 4480
rect 10735 4440 10784 4468
rect 10735 4437 10747 4440
rect 10689 4431 10747 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 13170 4468 13176 4480
rect 13131 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 17954 4468 17960 4480
rect 17915 4440 17960 4468
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 18690 4468 18696 4480
rect 18651 4440 18696 4468
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 22572 4468 22600 4567
rect 22830 4468 22836 4480
rect 22572 4440 22836 4468
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 23842 4428 23848 4480
rect 23900 4468 23906 4480
rect 23937 4471 23995 4477
rect 23937 4468 23949 4471
rect 23900 4440 23949 4468
rect 23900 4428 23906 4440
rect 23937 4437 23949 4440
rect 23983 4437 23995 4471
rect 23937 4431 23995 4437
rect 25225 4471 25283 4477
rect 25225 4437 25237 4471
rect 25271 4468 25283 4471
rect 27062 4468 27068 4480
rect 25271 4440 27068 4468
rect 25271 4437 25283 4440
rect 25225 4431 25283 4437
rect 27062 4428 27068 4440
rect 27120 4428 27126 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 5169 4267 5227 4273
rect 5169 4233 5181 4267
rect 5215 4264 5227 4267
rect 6457 4267 6515 4273
rect 5215 4236 6408 4264
rect 5215 4233 5227 4236
rect 5169 4227 5227 4233
rect 2038 4196 2044 4208
rect 1320 4168 2044 4196
rect 290 4088 296 4140
rect 348 4128 354 4140
rect 1320 4128 1348 4168
rect 2038 4156 2044 4168
rect 2096 4156 2102 4208
rect 4525 4199 4583 4205
rect 4525 4165 4537 4199
rect 4571 4196 4583 4199
rect 4893 4199 4951 4205
rect 4893 4196 4905 4199
rect 4571 4168 4905 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 4893 4165 4905 4168
rect 4939 4196 4951 4199
rect 5442 4196 5448 4208
rect 4939 4168 5448 4196
rect 4939 4165 4951 4168
rect 4893 4159 4951 4165
rect 5442 4156 5448 4168
rect 5500 4196 5506 4208
rect 6380 4196 6408 4236
rect 6457 4233 6469 4267
rect 6503 4264 6515 4267
rect 6914 4264 6920 4276
rect 6503 4236 6920 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 6914 4224 6920 4236
rect 6972 4224 6978 4276
rect 11146 4264 11152 4276
rect 11107 4236 11152 4264
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11606 4264 11612 4276
rect 11567 4236 11612 4264
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 12805 4267 12863 4273
rect 12805 4233 12817 4267
rect 12851 4264 12863 4267
rect 12851 4236 13860 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 6730 4196 6736 4208
rect 5500 4168 5764 4196
rect 6380 4168 6736 4196
rect 5500 4156 5506 4168
rect 5736 4137 5764 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 13170 4156 13176 4208
rect 13228 4196 13234 4208
rect 13832 4196 13860 4236
rect 13906 4224 13912 4276
rect 13964 4264 13970 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 13964 4236 14105 4264
rect 13964 4224 13970 4236
rect 14093 4233 14105 4236
rect 14139 4233 14151 4267
rect 14093 4227 14151 4233
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 15657 4267 15715 4273
rect 15657 4264 15669 4267
rect 14240 4236 15669 4264
rect 14240 4224 14246 4236
rect 15657 4233 15669 4236
rect 15703 4264 15715 4267
rect 15933 4267 15991 4273
rect 15933 4264 15945 4267
rect 15703 4236 15945 4264
rect 15703 4233 15715 4236
rect 15657 4227 15715 4233
rect 15933 4233 15945 4236
rect 15979 4233 15991 4267
rect 16206 4264 16212 4276
rect 16167 4236 16212 4264
rect 15933 4227 15991 4233
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 17313 4267 17371 4273
rect 17313 4233 17325 4267
rect 17359 4264 17371 4267
rect 17494 4264 17500 4276
rect 17359 4236 17500 4264
rect 17359 4233 17371 4236
rect 17313 4227 17371 4233
rect 17494 4224 17500 4236
rect 17552 4224 17558 4276
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 18233 4267 18291 4273
rect 18233 4264 18245 4267
rect 18012 4236 18245 4264
rect 18012 4224 18018 4236
rect 18233 4233 18245 4236
rect 18279 4233 18291 4267
rect 18233 4227 18291 4233
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19794 4264 19800 4276
rect 19383 4236 19800 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19794 4224 19800 4236
rect 19852 4224 19858 4276
rect 21634 4224 21640 4276
rect 21692 4264 21698 4276
rect 21729 4267 21787 4273
rect 21729 4264 21741 4267
rect 21692 4236 21741 4264
rect 21692 4224 21698 4236
rect 21729 4233 21741 4236
rect 21775 4233 21787 4267
rect 23382 4264 23388 4276
rect 23343 4236 23388 4264
rect 21729 4227 21787 4233
rect 23382 4224 23388 4236
rect 23440 4224 23446 4276
rect 25038 4224 25044 4276
rect 25096 4264 25102 4276
rect 25869 4267 25927 4273
rect 25869 4264 25881 4267
rect 25096 4236 25881 4264
rect 25096 4224 25102 4236
rect 25869 4233 25881 4236
rect 25915 4233 25927 4267
rect 25869 4227 25927 4233
rect 16942 4196 16948 4208
rect 13228 4168 13676 4196
rect 13832 4168 16948 4196
rect 13228 4156 13234 4168
rect 348 4100 1348 4128
rect 5721 4131 5779 4137
rect 348 4088 354 4100
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 5721 4091 5779 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7616 4100 7665 4128
rect 7616 4088 7622 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1872 4032 2053 4060
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 1872 3933 1900 4032
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 2308 4063 2366 4069
rect 2308 4029 2320 4063
rect 2354 4060 2366 4063
rect 2590 4060 2596 4072
rect 2354 4032 2596 4060
rect 2354 4029 2366 4032
rect 2308 4023 2366 4029
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 6178 4060 6184 4072
rect 5675 4032 6184 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 7668 4060 7696 4091
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10008 4100 10701 4128
rect 10008 4088 10014 4100
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 12124 4100 12173 4128
rect 12124 4088 12130 4100
rect 12161 4097 12173 4100
rect 12207 4128 12219 4131
rect 13446 4128 13452 4140
rect 12207 4100 13452 4128
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 13648 4137 13676 4168
rect 16942 4156 16948 4168
rect 17000 4196 17006 4208
rect 17773 4199 17831 4205
rect 17773 4196 17785 4199
rect 17000 4168 17785 4196
rect 17000 4156 17006 4168
rect 17773 4165 17785 4168
rect 17819 4196 17831 4199
rect 17819 4168 18644 4196
rect 17819 4165 17831 4168
rect 17773 4159 17831 4165
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 14792 4100 15209 4128
rect 14792 4088 14798 4100
rect 15197 4097 15209 4100
rect 15243 4097 15255 4131
rect 15197 4091 15255 4097
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 16448 4100 16773 4128
rect 16448 4088 16454 4100
rect 16761 4097 16773 4100
rect 16807 4097 16819 4131
rect 16761 4091 16819 4097
rect 8294 4060 8300 4072
rect 7668 4032 8300 4060
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 10778 4060 10784 4072
rect 10551 4032 10784 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 12894 4060 12900 4072
rect 12855 4032 12900 4060
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 14553 4063 14611 4069
rect 14553 4029 14565 4063
rect 14599 4060 14611 4063
rect 15105 4063 15163 4069
rect 15105 4060 15117 4063
rect 14599 4032 15117 4060
rect 14599 4029 14611 4032
rect 14553 4023 14611 4029
rect 15105 4029 15117 4032
rect 15151 4060 15163 4063
rect 15286 4060 15292 4072
rect 15151 4032 15292 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4060 16175 4063
rect 16206 4060 16212 4072
rect 16163 4032 16212 4060
rect 16163 4029 16175 4032
rect 16117 4023 16175 4029
rect 16206 4020 16212 4032
rect 16264 4060 16270 4072
rect 16577 4063 16635 4069
rect 16577 4060 16589 4063
rect 16264 4032 16589 4060
rect 16264 4020 16270 4032
rect 16577 4029 16589 4032
rect 16623 4060 16635 4063
rect 16850 4060 16856 4072
rect 16623 4032 16856 4060
rect 16623 4029 16635 4032
rect 16577 4023 16635 4029
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 18616 4069 18644 4168
rect 24578 4156 24584 4208
rect 24636 4196 24642 4208
rect 24636 4168 24716 4196
rect 24636 4156 24642 4168
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18748 4100 18797 4128
rect 18748 4088 18754 4100
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 20622 4128 20628 4140
rect 19935 4100 20628 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 20622 4088 20628 4100
rect 20680 4128 20686 4140
rect 24688 4137 24716 4168
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 20680 4100 21281 4128
rect 20680 4088 20686 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 24673 4131 24731 4137
rect 24673 4097 24685 4131
rect 24719 4128 24731 4131
rect 25133 4131 25191 4137
rect 25133 4128 25145 4131
rect 24719 4100 25145 4128
rect 24719 4097 24731 4100
rect 24673 4091 24731 4097
rect 25133 4097 25145 4100
rect 25179 4128 25191 4131
rect 25498 4128 25504 4140
rect 25179 4100 25504 4128
rect 25179 4097 25191 4100
rect 25133 4091 25191 4097
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4029 18659 4063
rect 18601 4023 18659 4029
rect 20441 4063 20499 4069
rect 20441 4029 20453 4063
rect 20487 4060 20499 4063
rect 21085 4063 21143 4069
rect 21085 4060 21097 4063
rect 20487 4032 21097 4060
rect 20487 4029 20499 4032
rect 20441 4023 20499 4029
rect 21085 4029 21097 4032
rect 21131 4029 21143 4063
rect 21085 4023 21143 4029
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22646 4060 22652 4072
rect 22511 4032 22652 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 22646 4020 22652 4032
rect 22704 4020 22710 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 23952 4032 24501 4060
rect 7926 4001 7932 4004
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 7920 3992 7932 4001
rect 7239 3964 7932 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 7920 3955 7932 3964
rect 7926 3952 7932 3955
rect 7984 3952 7990 4004
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 12912 3992 12940 4020
rect 13449 3995 13507 4001
rect 13449 3992 13461 3995
rect 9723 3964 10640 3992
rect 12912 3964 13461 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1636 3896 1869 3924
rect 1636 3884 1642 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 2924 3896 3433 3924
rect 2924 3884 2930 3896
rect 3421 3893 3433 3896
rect 3467 3924 3479 3927
rect 4062 3924 4068 3936
rect 3467 3896 4068 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6546 3924 6552 3936
rect 5592 3896 6552 3924
rect 5592 3884 5598 3896
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 9030 3924 9036 3936
rect 8991 3896 9036 3924
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10134 3924 10140 3936
rect 10095 3896 10140 3924
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10612 3933 10640 3964
rect 13449 3961 13461 3964
rect 13495 3961 13507 3995
rect 13449 3955 13507 3961
rect 15933 3995 15991 4001
rect 15933 3961 15945 3995
rect 15979 3992 15991 3995
rect 16666 3992 16672 4004
rect 15979 3964 16672 3992
rect 15979 3961 15991 3964
rect 15933 3955 15991 3961
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 20257 3995 20315 4001
rect 20257 3961 20269 3995
rect 20303 3992 20315 3995
rect 20303 3964 21220 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 21192 3936 21220 3964
rect 22094 3952 22100 4004
rect 22152 3992 22158 4004
rect 22189 3995 22247 4001
rect 22189 3992 22201 3995
rect 22152 3964 22201 3992
rect 22152 3952 22158 3964
rect 22189 3961 22201 3964
rect 22235 3992 22247 3995
rect 23842 3992 23848 4004
rect 22235 3964 23848 3992
rect 22235 3961 22247 3964
rect 22189 3955 22247 3961
rect 23842 3952 23848 3964
rect 23900 3952 23906 4004
rect 23952 3936 23980 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24489 4023 24547 4029
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 24581 3995 24639 4001
rect 24581 3992 24593 3995
rect 24268 3964 24593 3992
rect 24268 3952 24274 3964
rect 24581 3961 24593 3964
rect 24627 3992 24639 3995
rect 25501 3995 25559 4001
rect 25501 3992 25513 3995
rect 24627 3964 25513 3992
rect 24627 3961 24639 3964
rect 24581 3955 24639 3961
rect 25501 3961 25513 3964
rect 25547 3961 25559 3995
rect 25501 3955 25559 3961
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 10686 3924 10692 3936
rect 10643 3896 10692 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 11112 3896 12817 3924
rect 11112 3884 11118 3896
rect 12805 3893 12817 3896
rect 12851 3893 12863 3927
rect 13078 3924 13084 3936
rect 13039 3896 13084 3924
rect 12805 3887 12863 3893
rect 13078 3884 13084 3896
rect 13136 3884 13142 3936
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 13228 3896 13553 3924
rect 13228 3884 13234 3896
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 14642 3924 14648 3936
rect 14603 3896 14648 3924
rect 13541 3887 13599 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 15010 3924 15016 3936
rect 14971 3896 15016 3924
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 18693 3927 18751 3933
rect 18693 3893 18705 3927
rect 18739 3924 18751 3927
rect 18966 3924 18972 3936
rect 18739 3896 18972 3924
rect 18739 3893 18751 3896
rect 18693 3887 18751 3893
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 19484 3896 20453 3924
rect 19484 3884 19490 3896
rect 20441 3893 20453 3896
rect 20487 3924 20499 3927
rect 20533 3927 20591 3933
rect 20533 3924 20545 3927
rect 20487 3896 20545 3924
rect 20487 3893 20499 3896
rect 20441 3887 20499 3893
rect 20533 3893 20545 3896
rect 20579 3893 20591 3927
rect 20714 3924 20720 3936
rect 20675 3896 20720 3924
rect 20533 3887 20591 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 21174 3884 21180 3936
rect 21232 3924 21238 3936
rect 22646 3924 22652 3936
rect 21232 3896 21277 3924
rect 22607 3896 22652 3924
rect 21232 3884 21238 3896
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 22830 3884 22836 3936
rect 22888 3924 22894 3936
rect 23109 3927 23167 3933
rect 23109 3924 23121 3927
rect 22888 3896 23121 3924
rect 22888 3884 22894 3896
rect 23109 3893 23121 3896
rect 23155 3924 23167 3927
rect 23566 3924 23572 3936
rect 23155 3896 23572 3924
rect 23155 3893 23167 3896
rect 23109 3887 23167 3893
rect 23566 3884 23572 3896
rect 23624 3884 23630 3936
rect 23934 3924 23940 3936
rect 23895 3896 23940 3924
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 24118 3924 24124 3936
rect 24079 3896 24124 3924
rect 24118 3884 24124 3896
rect 24176 3884 24182 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2038 3720 2044 3732
rect 1999 3692 2044 3720
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2498 3720 2504 3732
rect 2459 3692 2504 3720
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2958 3720 2964 3732
rect 2648 3692 2964 3720
rect 2648 3680 2654 3692
rect 2958 3680 2964 3692
rect 3016 3720 3022 3732
rect 3053 3723 3111 3729
rect 3053 3720 3065 3723
rect 3016 3692 3065 3720
rect 3016 3680 3022 3692
rect 3053 3689 3065 3692
rect 3099 3720 3111 3723
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3099 3692 3433 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 6236 3692 6561 3720
rect 6236 3680 6242 3692
rect 6549 3689 6561 3692
rect 6595 3689 6607 3723
rect 6549 3683 6607 3689
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7834 3720 7840 3732
rect 7340 3692 7840 3720
rect 7340 3680 7346 3692
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 8478 3720 8484 3732
rect 8435 3692 8484 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 4310 3655 4368 3661
rect 4310 3652 4322 3655
rect 4120 3624 4322 3652
rect 4120 3612 4126 3624
rect 4310 3621 4322 3624
rect 4356 3621 4368 3655
rect 4310 3615 4368 3621
rect 7009 3655 7067 3661
rect 7009 3621 7021 3655
rect 7055 3652 7067 3655
rect 7558 3652 7564 3664
rect 7055 3624 7564 3652
rect 7055 3621 7067 3624
rect 7009 3615 7067 3621
rect 7558 3612 7564 3624
rect 7616 3652 7622 3664
rect 7742 3652 7748 3664
rect 7616 3624 7748 3652
rect 7616 3612 7622 3624
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 1946 3544 1952 3596
rect 2004 3584 2010 3596
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 2004 3556 2421 3584
rect 2004 3544 2010 3556
rect 2409 3553 2421 3556
rect 2455 3584 2467 3587
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 2455 3556 6193 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 6181 3553 6193 3556
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6604 3556 6929 3584
rect 6604 3544 6610 3556
rect 6917 3553 6929 3556
rect 6963 3553 6975 3587
rect 6917 3547 6975 3553
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7929 3587 7987 3593
rect 7929 3584 7941 3587
rect 7156 3556 7941 3584
rect 7156 3544 7162 3556
rect 7929 3553 7941 3556
rect 7975 3584 7987 3587
rect 8202 3584 8208 3596
rect 7975 3556 8208 3584
rect 7975 3553 7987 3556
rect 7929 3547 7987 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2866 3516 2872 3528
rect 2731 3488 2872 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 4062 3516 4068 3528
rect 4023 3488 4068 3516
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3516 7251 3519
rect 8404 3516 8432 3683
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 9306 3720 9312 3732
rect 8619 3692 9312 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 10321 3723 10379 3729
rect 10321 3720 10333 3723
rect 10100 3692 10333 3720
rect 10100 3680 10106 3692
rect 10321 3689 10333 3692
rect 10367 3689 10379 3723
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10321 3683 10379 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11146 3720 11152 3732
rect 10888 3692 11152 3720
rect 8662 3612 8668 3664
rect 8720 3652 8726 3664
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8720 3624 9045 3652
rect 8720 3612 8726 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9033 3615 9091 3621
rect 9048 3584 9076 3615
rect 9582 3584 9588 3596
rect 9048 3556 9588 3584
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 9769 3587 9827 3593
rect 9769 3553 9781 3587
rect 9815 3584 9827 3587
rect 10060 3584 10088 3680
rect 10888 3593 10916 3692
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 12250 3720 12256 3732
rect 12211 3692 12256 3720
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 12400 3692 13093 3720
rect 12400 3680 12406 3692
rect 13081 3689 13093 3692
rect 13127 3720 13139 3723
rect 13170 3720 13176 3732
rect 13127 3692 13176 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13354 3720 13360 3732
rect 13315 3692 13360 3720
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13504 3692 13737 3720
rect 13504 3680 13510 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14976 3692 15025 3720
rect 14976 3680 14982 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15286 3720 15292 3732
rect 15247 3692 15292 3720
rect 15013 3683 15071 3689
rect 15286 3680 15292 3692
rect 15344 3680 15350 3732
rect 15562 3680 15568 3732
rect 15620 3720 15626 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 15620 3692 15669 3720
rect 15620 3680 15626 3692
rect 15657 3689 15669 3692
rect 15703 3689 15715 3723
rect 16390 3720 16396 3732
rect 16351 3692 16396 3720
rect 15657 3683 15715 3689
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 16761 3723 16819 3729
rect 16761 3689 16773 3723
rect 16807 3720 16819 3723
rect 17218 3720 17224 3732
rect 16807 3692 17224 3720
rect 16807 3689 16819 3692
rect 16761 3683 16819 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17402 3720 17408 3732
rect 17363 3692 17408 3720
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18509 3723 18567 3729
rect 18509 3720 18521 3723
rect 18012 3692 18521 3720
rect 18012 3680 18018 3692
rect 18509 3689 18521 3692
rect 18555 3689 18567 3723
rect 18509 3683 18567 3689
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 19061 3723 19119 3729
rect 19061 3720 19073 3723
rect 18748 3692 19073 3720
rect 18748 3680 18754 3692
rect 19061 3689 19073 3692
rect 19107 3689 19119 3723
rect 19061 3683 19119 3689
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 20257 3723 20315 3729
rect 20257 3720 20269 3723
rect 19392 3692 20269 3720
rect 19392 3680 19398 3692
rect 20257 3689 20269 3692
rect 20303 3689 20315 3723
rect 20898 3720 20904 3732
rect 20859 3692 20904 3720
rect 20257 3683 20315 3689
rect 20898 3680 20904 3692
rect 20956 3680 20962 3732
rect 21082 3680 21088 3732
rect 21140 3720 21146 3732
rect 21269 3723 21327 3729
rect 21269 3720 21281 3723
rect 21140 3692 21281 3720
rect 21140 3680 21146 3692
rect 21269 3689 21281 3692
rect 21315 3689 21327 3723
rect 21910 3720 21916 3732
rect 21871 3692 21916 3720
rect 21269 3683 21327 3689
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22186 3680 22192 3732
rect 22244 3720 22250 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 22244 3692 22293 3720
rect 22244 3680 22250 3692
rect 22281 3689 22293 3692
rect 22327 3689 22339 3723
rect 22281 3683 22339 3689
rect 14642 3612 14648 3664
rect 14700 3652 14706 3664
rect 15749 3655 15807 3661
rect 15749 3652 15761 3655
rect 14700 3624 15761 3652
rect 14700 3612 14706 3624
rect 15749 3621 15761 3624
rect 15795 3621 15807 3655
rect 15749 3615 15807 3621
rect 17310 3612 17316 3664
rect 17368 3652 17374 3664
rect 18417 3655 18475 3661
rect 18417 3652 18429 3655
rect 17368 3624 18429 3652
rect 17368 3612 17374 3624
rect 18417 3621 18429 3624
rect 18463 3621 18475 3655
rect 19518 3652 19524 3664
rect 19479 3624 19524 3652
rect 18417 3615 18475 3621
rect 19518 3612 19524 3624
rect 19576 3612 19582 3664
rect 20717 3655 20775 3661
rect 20717 3621 20729 3655
rect 20763 3652 20775 3655
rect 20806 3652 20812 3664
rect 20763 3624 20812 3652
rect 20763 3621 20775 3624
rect 20717 3615 20775 3621
rect 20806 3612 20812 3624
rect 20864 3612 20870 3664
rect 21174 3612 21180 3664
rect 21232 3652 21238 3664
rect 21358 3652 21364 3664
rect 21232 3624 21364 3652
rect 21232 3612 21238 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 9815 3556 10088 3584
rect 10873 3587 10931 3593
rect 9815 3553 9827 3556
rect 9769 3547 9827 3553
rect 10873 3553 10885 3587
rect 10919 3553 10931 3587
rect 10873 3547 10931 3553
rect 11140 3587 11198 3593
rect 11140 3553 11152 3587
rect 11186 3584 11198 3587
rect 11514 3584 11520 3596
rect 11186 3556 11520 3584
rect 11186 3553 11198 3556
rect 11140 3547 11198 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 16850 3584 16856 3596
rect 16811 3556 16856 3584
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3584 19763 3587
rect 21928 3584 21956 3680
rect 19751 3556 21956 3584
rect 22296 3584 22324 3683
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 23017 3723 23075 3729
rect 23017 3720 23029 3723
rect 22796 3692 23029 3720
rect 22796 3680 22802 3692
rect 23017 3689 23029 3692
rect 23063 3689 23075 3723
rect 23017 3683 23075 3689
rect 23842 3661 23848 3664
rect 23836 3652 23848 3661
rect 23803 3624 23848 3652
rect 23836 3615 23848 3624
rect 23842 3612 23848 3615
rect 23900 3612 23906 3664
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22296 3556 22477 3584
rect 19751 3553 19763 3556
rect 19705 3547 19763 3553
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 22465 3547 22523 3553
rect 13814 3516 13820 3528
rect 7239 3488 8432 3516
rect 13775 3488 13820 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 5445 3451 5503 3457
rect 5445 3417 5457 3451
rect 5491 3448 5503 3451
rect 6270 3448 6276 3460
rect 5491 3420 6276 3448
rect 5491 3417 5503 3420
rect 5445 3411 5503 3417
rect 6270 3408 6276 3420
rect 6328 3448 6334 3460
rect 6457 3451 6515 3457
rect 6457 3448 6469 3451
rect 6328 3420 6469 3448
rect 6328 3408 6334 3420
rect 6457 3417 6469 3420
rect 6503 3448 6515 3451
rect 7208 3448 7236 3479
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 15838 3516 15844 3528
rect 15799 3488 15844 3516
rect 13909 3479 13967 3485
rect 9401 3451 9459 3457
rect 9401 3448 9413 3451
rect 6503 3420 7236 3448
rect 7300 3420 9413 3448
rect 6503 3417 6515 3420
rect 6457 3411 6515 3417
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 3881 3383 3939 3389
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 4338 3380 4344 3392
rect 3927 3352 4344 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 6086 3380 6092 3392
rect 6047 3352 6092 3380
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6181 3383 6239 3389
rect 6181 3349 6193 3383
rect 6227 3380 6239 3383
rect 7300 3380 7328 3420
rect 9401 3417 9413 3420
rect 9447 3417 9459 3451
rect 9401 3411 9459 3417
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 13924 3448 13952 3479
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18564 3488 18613 3516
rect 18564 3476 18570 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21358 3516 21364 3528
rect 20772 3488 21364 3516
rect 20772 3476 20778 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 23566 3516 23572 3528
rect 21508 3488 21553 3516
rect 23527 3488 23572 3516
rect 21508 3476 21514 3488
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 13596 3420 13952 3448
rect 13596 3408 13602 3420
rect 15010 3408 15016 3460
rect 15068 3408 15074 3460
rect 17957 3451 18015 3457
rect 17957 3417 17969 3451
rect 18003 3448 18015 3451
rect 18138 3448 18144 3460
rect 18003 3420 18144 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 18138 3408 18144 3420
rect 18196 3408 18202 3460
rect 22646 3448 22652 3460
rect 22607 3420 22652 3448
rect 22646 3408 22652 3420
rect 22704 3408 22710 3460
rect 6227 3352 7328 3380
rect 6227 3349 6239 3352
rect 6181 3343 6239 3349
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 7524 3352 7573 3380
rect 7524 3340 7530 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 9950 3380 9956 3392
rect 9911 3352 9956 3380
rect 7561 3343 7619 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14645 3383 14703 3389
rect 14645 3380 14657 3383
rect 14608 3352 14657 3380
rect 14608 3340 14614 3352
rect 14645 3349 14657 3352
rect 14691 3380 14703 3383
rect 15028 3380 15056 3408
rect 17034 3380 17040 3392
rect 14691 3352 15056 3380
rect 16995 3352 17040 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 18049 3383 18107 3389
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 18782 3380 18788 3392
rect 18095 3352 18788 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 19886 3380 19892 3392
rect 19847 3352 19892 3380
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 23477 3383 23535 3389
rect 23477 3349 23489 3383
rect 23523 3380 23535 3383
rect 24762 3380 24768 3392
rect 23523 3352 24768 3380
rect 23523 3349 23535 3352
rect 23477 3343 23535 3349
rect 24762 3340 24768 3352
rect 24820 3380 24826 3392
rect 24949 3383 25007 3389
rect 24949 3380 24961 3383
rect 24820 3352 24961 3380
rect 24820 3340 24826 3352
rect 24949 3349 24961 3352
rect 24995 3349 25007 3383
rect 24949 3343 25007 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3418 3136 3424 3188
rect 3476 3176 3482 3188
rect 3476 3148 5212 3176
rect 3476 3136 3482 3148
rect 5184 3108 5212 3148
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 6144 3148 6837 3176
rect 6144 3136 6150 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7248 3148 7849 3176
rect 7248 3136 7254 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 8665 3179 8723 3185
rect 8665 3176 8677 3179
rect 8352 3148 8677 3176
rect 8352 3136 8358 3148
rect 8665 3145 8677 3148
rect 8711 3145 8723 3179
rect 8665 3139 8723 3145
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11146 3176 11152 3188
rect 11011 3148 11152 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 7208 3108 7236 3136
rect 5184 3080 7236 3108
rect 6270 3040 6276 3052
rect 6183 3012 6276 3040
rect 6270 3000 6276 3012
rect 6328 3040 6334 3052
rect 7282 3040 7288 3052
rect 6328 3012 7288 3040
rect 6328 3000 6334 3012
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 8680 3040 8708 3139
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13538 3176 13544 3188
rect 12492 3148 12537 3176
rect 13499 3148 13544 3176
rect 12492 3136 12498 3148
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 14090 3136 14096 3188
rect 14148 3176 14154 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14148 3148 14473 3176
rect 14148 3136 14154 3148
rect 14461 3145 14473 3148
rect 14507 3176 14519 3179
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14507 3148 14565 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 15896 3148 16129 3176
rect 15896 3136 15902 3148
rect 16117 3145 16129 3148
rect 16163 3176 16175 3179
rect 17037 3179 17095 3185
rect 17037 3176 17049 3179
rect 16163 3148 17049 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 17037 3145 17049 3148
rect 17083 3145 17095 3179
rect 17037 3139 17095 3145
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17368 3148 17417 3176
rect 17368 3136 17374 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17405 3139 17463 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18690 3136 18696 3188
rect 18748 3176 18754 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 18748 3148 19441 3176
rect 18748 3136 18754 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 19429 3139 19487 3145
rect 20165 3179 20223 3185
rect 20165 3145 20177 3179
rect 20211 3176 20223 3179
rect 20990 3176 20996 3188
rect 20211 3148 20996 3176
rect 20211 3145 20223 3148
rect 20165 3139 20223 3145
rect 20990 3136 20996 3148
rect 21048 3136 21054 3188
rect 21542 3136 21548 3188
rect 21600 3176 21606 3188
rect 22554 3176 22560 3188
rect 21600 3148 22560 3176
rect 21600 3136 21606 3148
rect 22554 3136 22560 3148
rect 22612 3136 22618 3188
rect 23109 3179 23167 3185
rect 23109 3145 23121 3179
rect 23155 3176 23167 3179
rect 23842 3176 23848 3188
rect 23155 3148 23848 3176
rect 23155 3145 23167 3148
rect 23109 3139 23167 3145
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 25498 3176 25504 3188
rect 25459 3148 25504 3176
rect 25498 3136 25504 3148
rect 25556 3136 25562 3188
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 11885 3111 11943 3117
rect 11885 3108 11897 3111
rect 11848 3080 11897 3108
rect 11848 3068 11854 3080
rect 11885 3077 11897 3080
rect 11931 3108 11943 3111
rect 11974 3108 11980 3120
rect 11931 3080 11980 3108
rect 11931 3077 11943 3080
rect 11885 3071 11943 3077
rect 11974 3068 11980 3080
rect 12032 3068 12038 3120
rect 12342 3068 12348 3120
rect 12400 3108 12406 3120
rect 12400 3080 13124 3108
rect 12400 3068 12406 3080
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 8680 3012 8861 3040
rect 7377 3003 7435 3009
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 11330 3040 11336 3052
rect 11291 3012 11336 3040
rect 8849 3003 8907 3009
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2972 1642 2984
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 1636 2944 3709 2972
rect 1636 2932 1642 2944
rect 3697 2941 3709 2944
rect 3743 2972 3755 2975
rect 3878 2972 3884 2984
rect 3743 2944 3884 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 3878 2932 3884 2944
rect 3936 2972 3942 2984
rect 4062 2972 4068 2984
rect 3936 2944 4068 2972
rect 3936 2932 3942 2944
rect 4062 2932 4068 2944
rect 4120 2972 4126 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4120 2944 4261 2972
rect 4120 2932 4126 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 4338 2932 4344 2984
rect 4396 2972 4402 2984
rect 4505 2975 4563 2981
rect 4505 2972 4517 2975
rect 4396 2944 4517 2972
rect 4396 2932 4402 2944
rect 4505 2941 4517 2944
rect 4551 2972 4563 2975
rect 5626 2972 5632 2984
rect 4551 2944 5632 2972
rect 4551 2941 4563 2944
rect 4505 2935 4563 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 7190 2972 7196 2984
rect 7151 2944 7196 2972
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 1670 2864 1676 2916
rect 1728 2904 1734 2916
rect 1848 2907 1906 2913
rect 1848 2904 1860 2907
rect 1728 2876 1860 2904
rect 1728 2864 1734 2876
rect 1848 2873 1860 2876
rect 1894 2904 1906 2907
rect 2682 2904 2688 2916
rect 1894 2876 2688 2904
rect 1894 2873 1906 2876
rect 1848 2867 1906 2873
rect 2682 2864 2688 2876
rect 2740 2904 2746 2916
rect 7392 2904 7420 3003
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 12894 3040 12900 3052
rect 12855 3012 12900 3040
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 13096 3049 13124 3080
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13556 3040 13584 3136
rect 13127 3012 13584 3040
rect 14277 3043 14335 3049
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 14277 3009 14289 3043
rect 14323 3040 14335 3043
rect 17788 3040 17816 3136
rect 26050 3108 26056 3120
rect 26011 3080 26056 3108
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 18046 3040 18052 3052
rect 14323 3012 14872 3040
rect 17788 3012 18052 3040
rect 14323 3009 14335 3012
rect 14277 3003 14335 3009
rect 14844 2984 14872 3012
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 8662 2932 8668 2984
rect 8720 2972 8726 2984
rect 9105 2975 9163 2981
rect 9105 2972 9117 2975
rect 8720 2944 9117 2972
rect 8720 2932 8726 2944
rect 9105 2941 9117 2944
rect 9151 2941 9163 2975
rect 9105 2935 9163 2941
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 10134 2972 10140 2984
rect 9732 2944 10140 2972
rect 9732 2932 9738 2944
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 12158 2972 12164 2984
rect 12119 2944 12164 2972
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12584 2944 12817 2972
rect 12584 2932 12590 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 14734 2972 14740 2984
rect 14507 2944 14740 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 15010 2981 15016 2984
rect 14993 2975 15016 2981
rect 14993 2972 15005 2975
rect 14884 2944 15005 2972
rect 14884 2932 14890 2944
rect 14993 2941 15005 2944
rect 15068 2972 15074 2984
rect 15068 2944 15141 2972
rect 14993 2935 15016 2941
rect 15010 2932 15016 2935
rect 15068 2932 15074 2944
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 15620 2944 16681 2972
rect 15620 2932 15626 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 20898 2981 20904 2984
rect 18305 2975 18363 2981
rect 18305 2972 18317 2975
rect 18196 2944 18317 2972
rect 18196 2932 18202 2944
rect 18305 2941 18317 2944
rect 18351 2941 18363 2975
rect 18305 2935 18363 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 20625 2975 20683 2981
rect 20625 2972 20637 2975
rect 20579 2944 20637 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 20625 2941 20637 2944
rect 20671 2941 20683 2975
rect 20892 2972 20904 2981
rect 20859 2944 20904 2972
rect 20625 2935 20683 2941
rect 20892 2935 20904 2944
rect 7466 2904 7472 2916
rect 2740 2876 7472 2904
rect 2740 2864 2746 2876
rect 5644 2845 5672 2876
rect 7466 2864 7472 2876
rect 7524 2864 7530 2916
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 8297 2907 8355 2913
rect 8297 2904 8309 2907
rect 7616 2876 8309 2904
rect 7616 2864 7622 2876
rect 8297 2873 8309 2876
rect 8343 2904 8355 2907
rect 8343 2876 14504 2904
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 5629 2839 5687 2845
rect 5629 2805 5641 2839
rect 5675 2805 5687 2839
rect 6546 2836 6552 2848
rect 6507 2808 6552 2836
rect 5629 2799 5687 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 9916 2808 10241 2836
rect 9916 2796 9922 2808
rect 10229 2805 10241 2808
rect 10275 2836 10287 2839
rect 10686 2836 10692 2848
rect 10275 2808 10692 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 13814 2836 13820 2848
rect 11664 2808 13820 2836
rect 11664 2796 11670 2808
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14476 2836 14504 2876
rect 17218 2836 17224 2848
rect 14476 2808 17224 2836
rect 17218 2796 17224 2808
rect 17276 2796 17282 2848
rect 20640 2836 20668 2935
rect 20898 2932 20904 2935
rect 20956 2932 20962 2984
rect 22094 2932 22100 2984
rect 22152 2972 22158 2984
rect 23385 2975 23443 2981
rect 23385 2972 23397 2975
rect 22152 2944 23397 2972
rect 22152 2932 22158 2944
rect 23385 2941 23397 2944
rect 23431 2972 23443 2975
rect 23566 2972 23572 2984
rect 23431 2944 23572 2972
rect 23431 2941 23443 2944
rect 23385 2935 23443 2941
rect 23566 2932 23572 2944
rect 23624 2972 23630 2984
rect 23937 2975 23995 2981
rect 23937 2972 23949 2975
rect 23624 2944 23949 2972
rect 23624 2932 23630 2944
rect 23937 2941 23949 2944
rect 23983 2972 23995 2975
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 23983 2944 24133 2972
rect 23983 2941 23995 2944
rect 23937 2935 23995 2941
rect 24121 2941 24133 2944
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 24388 2975 24446 2981
rect 24388 2941 24400 2975
rect 24434 2972 24446 2975
rect 24762 2972 24768 2984
rect 24434 2944 24768 2972
rect 24434 2941 24446 2944
rect 24388 2935 24446 2941
rect 24762 2932 24768 2944
rect 24820 2932 24826 2984
rect 23750 2864 23756 2916
rect 23808 2904 23814 2916
rect 23808 2876 24164 2904
rect 23808 2864 23814 2876
rect 24136 2848 24164 2876
rect 20806 2836 20812 2848
rect 20640 2808 20812 2836
rect 20806 2796 20812 2808
rect 20864 2796 20870 2848
rect 22002 2836 22008 2848
rect 21963 2808 22008 2836
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 22554 2836 22560 2848
rect 22515 2808 22560 2836
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 24118 2796 24124 2848
rect 24176 2796 24182 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 1946 2632 1952 2644
rect 1903 2604 1952 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3878 2632 3884 2644
rect 3839 2604 3884 2632
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5684 2604 5733 2632
rect 5684 2592 5690 2604
rect 5721 2601 5733 2604
rect 5767 2632 5779 2635
rect 6362 2632 6368 2644
rect 5767 2604 6368 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2601 6975 2635
rect 6917 2595 6975 2601
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 9674 2632 9680 2644
rect 8527 2604 9680 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 1762 2524 1768 2576
rect 1820 2564 1826 2576
rect 2225 2567 2283 2573
rect 2225 2564 2237 2567
rect 1820 2536 2237 2564
rect 1820 2524 1826 2536
rect 2225 2533 2237 2536
rect 2271 2533 2283 2567
rect 2225 2527 2283 2533
rect 3896 2496 3924 2592
rect 4246 2524 4252 2576
rect 4304 2564 4310 2576
rect 6932 2564 6960 2595
rect 4304 2536 6960 2564
rect 4304 2524 4310 2536
rect 4614 2505 4620 2508
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 3896 2468 4353 2496
rect 4341 2465 4353 2468
rect 4387 2465 4399 2499
rect 4608 2496 4620 2505
rect 4341 2459 4399 2465
rect 4448 2468 4620 2496
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 2958 2428 2964 2440
rect 2547 2400 2964 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 4448 2428 4476 2468
rect 4608 2459 4620 2468
rect 4614 2456 4620 2459
rect 4672 2456 4678 2508
rect 6362 2496 6368 2508
rect 6275 2468 6368 2496
rect 6362 2456 6368 2468
rect 6420 2496 6426 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6420 2468 7297 2496
rect 6420 2456 6426 2468
rect 7285 2465 7297 2468
rect 7331 2496 7343 2499
rect 7558 2496 7564 2508
rect 7331 2468 7564 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 8588 2505 8616 2604
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 11606 2632 11612 2644
rect 9815 2604 11612 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 11992 2604 14013 2632
rect 10965 2567 11023 2573
rect 10965 2533 10977 2567
rect 11011 2564 11023 2567
rect 11514 2564 11520 2576
rect 11011 2536 11520 2564
rect 11011 2533 11023 2536
rect 10965 2527 11023 2533
rect 11514 2524 11520 2536
rect 11572 2564 11578 2576
rect 11992 2564 12020 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 14001 2595 14059 2601
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 15197 2635 15255 2641
rect 15197 2632 15209 2635
rect 14792 2604 15209 2632
rect 14792 2592 14798 2604
rect 15197 2601 15209 2604
rect 15243 2601 15255 2635
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 15197 2595 15255 2601
rect 11572 2536 12020 2564
rect 12069 2567 12127 2573
rect 11572 2524 11578 2536
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12710 2564 12716 2576
rect 12115 2536 12716 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 12710 2524 12716 2536
rect 12768 2564 12774 2576
rect 12866 2567 12924 2573
rect 12866 2564 12878 2567
rect 12768 2536 12878 2564
rect 12768 2524 12774 2536
rect 12866 2533 12878 2536
rect 12912 2533 12924 2567
rect 12866 2527 12924 2533
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2465 8631 2499
rect 8573 2459 8631 2465
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 10042 2496 10048 2508
rect 9631 2468 10048 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 3559 2400 4476 2428
rect 6733 2431 6791 2437
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7374 2428 7380 2440
rect 6779 2400 7380 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7524 2400 7941 2428
rect 7524 2388 7530 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 9600 2428 9628 2459
rect 10042 2456 10048 2468
rect 10100 2496 10106 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 10100 2468 10149 2496
rect 10100 2456 10106 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10686 2496 10692 2508
rect 10137 2459 10195 2465
rect 10428 2468 10692 2496
rect 10226 2428 10232 2440
rect 8168 2400 9628 2428
rect 10139 2400 10232 2428
rect 8168 2388 8174 2400
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10428 2437 10456 2468
rect 10686 2456 10692 2468
rect 10744 2496 10750 2508
rect 11241 2499 11299 2505
rect 11241 2496 11253 2499
rect 10744 2468 11253 2496
rect 10744 2456 10750 2468
rect 11241 2465 11253 2468
rect 11287 2465 11299 2499
rect 11241 2459 11299 2465
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11790 2496 11796 2508
rect 11471 2468 11796 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 15212 2496 15240 2595
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18506 2632 18512 2644
rect 18419 2604 18512 2632
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15212 2468 15485 2496
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15729 2499 15787 2505
rect 15729 2496 15741 2499
rect 15473 2459 15531 2465
rect 15580 2468 15741 2496
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 11204 2400 12357 2428
rect 11204 2388 11210 2400
rect 12345 2397 12357 2400
rect 12391 2428 12403 2431
rect 12621 2431 12679 2437
rect 12621 2428 12633 2431
rect 12391 2400 12633 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12621 2397 12633 2400
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15580 2428 15608 2468
rect 15729 2465 15741 2468
rect 15775 2496 15787 2499
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 15775 2468 17693 2496
rect 15775 2465 15787 2468
rect 15729 2459 15787 2465
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 18064 2496 18092 2592
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18064 2468 18337 2496
rect 17681 2459 17739 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 14967 2400 15608 2428
rect 17696 2428 17724 2459
rect 18432 2428 18460 2604
rect 18506 2592 18512 2604
rect 18564 2632 18570 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 18564 2604 19717 2632
rect 18564 2592 18570 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 20806 2592 20812 2644
rect 20864 2632 20870 2644
rect 20993 2635 21051 2641
rect 20993 2632 21005 2635
rect 20864 2604 21005 2632
rect 20864 2592 20870 2604
rect 20993 2601 21005 2604
rect 21039 2632 21051 2635
rect 21910 2632 21916 2644
rect 21039 2604 21916 2632
rect 21039 2601 21051 2604
rect 20993 2595 21051 2601
rect 18592 2567 18650 2573
rect 18592 2533 18604 2567
rect 18638 2564 18650 2567
rect 18690 2564 18696 2576
rect 18638 2536 18696 2564
rect 18638 2533 18650 2536
rect 18592 2527 18650 2533
rect 18690 2524 18696 2536
rect 18748 2524 18754 2576
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 20714 2564 20720 2576
rect 20671 2536 20720 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 20714 2524 20720 2536
rect 20772 2524 20778 2576
rect 21192 2505 21220 2604
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 22554 2632 22560 2644
rect 22515 2604 22560 2632
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 24210 2632 24216 2644
rect 24171 2604 24216 2632
rect 24210 2592 24216 2604
rect 24268 2592 24274 2644
rect 21450 2573 21456 2576
rect 21444 2564 21456 2573
rect 21411 2536 21456 2564
rect 21444 2527 21456 2536
rect 21450 2524 21456 2527
rect 21508 2524 21514 2576
rect 21177 2499 21235 2505
rect 21177 2465 21189 2499
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 23750 2456 23756 2508
rect 23808 2496 23814 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 23808 2468 24593 2496
rect 23808 2456 23814 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 17696 2400 18460 2428
rect 23477 2431 23535 2437
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 23477 2397 23489 2431
rect 23523 2428 23535 2431
rect 24670 2428 24676 2440
rect 23523 2400 24676 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 24820 2400 25237 2428
rect 24820 2388 24826 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 9122 2360 9128 2372
rect 9083 2332 9128 2360
rect 9122 2320 9128 2332
rect 9180 2360 9186 2372
rect 10244 2360 10272 2388
rect 9180 2332 10272 2360
rect 9180 2320 9186 2332
rect 8754 2292 8760 2304
rect 8715 2264 8760 2292
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 23750 2292 23756 2304
rect 23711 2264 23756 2292
rect 23750 2252 23756 2264
rect 23808 2252 23814 2304
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24762 2292 24768 2304
rect 24084 2264 24768 2292
rect 24084 2252 24090 2264
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 19426 620 19432 672
rect 19484 660 19490 672
rect 19484 632 21312 660
rect 19484 620 19490 632
rect 21284 604 21312 632
rect 4338 552 4344 604
rect 4396 592 4402 604
rect 5258 592 5264 604
rect 4396 564 5264 592
rect 4396 552 4402 564
rect 5258 552 5264 564
rect 5316 552 5322 604
rect 8202 552 8208 604
rect 8260 592 8266 604
rect 9582 592 9588 604
rect 8260 564 9588 592
rect 8260 552 8266 564
rect 9582 552 9588 564
rect 9640 552 9646 604
rect 20162 552 20168 604
rect 20220 592 20226 604
rect 20622 592 20628 604
rect 20220 564 20628 592
rect 20220 552 20226 564
rect 20622 552 20628 564
rect 20680 552 20686 604
rect 21266 552 21272 604
rect 21324 552 21330 604
<< via1 >>
rect 14096 26256 14148 26308
rect 24768 26256 24820 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 24676 23128 24728 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 23664 22559 23716 22568
rect 23664 22525 23673 22559
rect 23673 22525 23707 22559
rect 23707 22525 23716 22559
rect 23664 22516 23716 22525
rect 1400 22380 1452 22432
rect 2688 22380 2740 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 24676 21972 24728 22024
rect 24768 21947 24820 21956
rect 24768 21913 24777 21947
rect 24777 21913 24811 21947
rect 24811 21913 24820 21947
rect 24768 21904 24820 21913
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 24584 21335 24636 21344
rect 24584 21301 24593 21335
rect 24593 21301 24627 21335
rect 24627 21301 24636 21335
rect 24584 21292 24636 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 24216 20952 24268 21004
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 2688 20587 2740 20596
rect 2688 20553 2697 20587
rect 2697 20553 2731 20587
rect 2731 20553 2740 20587
rect 2688 20544 2740 20553
rect 13452 20383 13504 20392
rect 13452 20349 13461 20383
rect 13461 20349 13495 20383
rect 13495 20349 13504 20383
rect 13452 20340 13504 20349
rect 13728 20383 13780 20392
rect 13728 20349 13762 20383
rect 13762 20349 13780 20383
rect 13728 20340 13780 20349
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 3056 20247 3108 20256
rect 3056 20213 3065 20247
rect 3065 20213 3099 20247
rect 3099 20213 3108 20247
rect 3056 20204 3108 20213
rect 14648 20204 14700 20256
rect 24216 20204 24268 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1492 20000 1544 20052
rect 2044 20000 2096 20052
rect 2412 19864 2464 19916
rect 2596 19864 2648 19916
rect 13452 19703 13504 19712
rect 13452 19669 13461 19703
rect 13461 19669 13495 19703
rect 13495 19669 13504 19703
rect 13452 19660 13504 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1860 19320 1912 19372
rect 3332 19320 3384 19372
rect 1676 19252 1728 19304
rect 13820 19184 13872 19236
rect 1400 19116 1452 19168
rect 2412 19116 2464 19168
rect 2596 19159 2648 19168
rect 2596 19125 2605 19159
rect 2605 19125 2639 19159
rect 2639 19125 2648 19159
rect 2596 19116 2648 19125
rect 13452 19116 13504 19168
rect 14832 19159 14884 19168
rect 14832 19125 14841 19159
rect 14841 19125 14875 19159
rect 14875 19125 14884 19159
rect 14832 19116 14884 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 12348 18955 12400 18964
rect 12348 18921 12357 18955
rect 12357 18921 12391 18955
rect 12391 18921 12400 18955
rect 12348 18912 12400 18921
rect 12900 18776 12952 18828
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 12440 18708 12492 18760
rect 14832 18776 14884 18828
rect 13912 18751 13964 18760
rect 12256 18640 12308 18692
rect 13912 18717 13921 18751
rect 13921 18717 13955 18751
rect 13955 18717 13964 18751
rect 13912 18708 13964 18717
rect 10968 18572 11020 18624
rect 13820 18572 13872 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 12440 18368 12492 18420
rect 9680 18300 9732 18352
rect 12256 18343 12308 18352
rect 12256 18309 12265 18343
rect 12265 18309 12299 18343
rect 12299 18309 12308 18343
rect 12256 18300 12308 18309
rect 10968 18275 11020 18284
rect 10968 18241 10977 18275
rect 10977 18241 11011 18275
rect 11011 18241 11020 18275
rect 10968 18232 11020 18241
rect 10048 18096 10100 18148
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 9772 18028 9824 18080
rect 11428 18028 11480 18080
rect 12716 18139 12768 18148
rect 12716 18105 12750 18139
rect 12750 18105 12768 18139
rect 12716 18096 12768 18105
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1768 17824 1820 17876
rect 9588 17824 9640 17876
rect 11336 17824 11388 17876
rect 12900 17824 12952 17876
rect 14648 17867 14700 17876
rect 14648 17833 14657 17867
rect 14657 17833 14691 17867
rect 14691 17833 14700 17867
rect 14648 17824 14700 17833
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 12716 17756 12768 17808
rect 2320 17688 2372 17740
rect 10324 17688 10376 17740
rect 11888 17688 11940 17740
rect 13544 17688 13596 17740
rect 13912 17731 13964 17740
rect 13912 17697 13921 17731
rect 13921 17697 13955 17731
rect 13955 17697 13964 17731
rect 13912 17688 13964 17697
rect 24676 17688 24728 17740
rect 14004 17663 14056 17672
rect 10048 17484 10100 17536
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 14004 17629 14013 17663
rect 14013 17629 14047 17663
rect 14047 17629 14056 17663
rect 14004 17620 14056 17629
rect 13820 17552 13872 17604
rect 24584 17552 24636 17604
rect 24768 17552 24820 17604
rect 11428 17484 11480 17536
rect 13360 17527 13412 17536
rect 13360 17493 13369 17527
rect 13369 17493 13403 17527
rect 13403 17493 13412 17527
rect 13360 17484 13412 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1492 17280 1544 17332
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 10324 17323 10376 17332
rect 10324 17289 10333 17323
rect 10333 17289 10367 17323
rect 10367 17289 10376 17323
rect 10324 17280 10376 17289
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 24768 17323 24820 17332
rect 12440 17280 12492 17289
rect 24768 17289 24777 17323
rect 24777 17289 24811 17323
rect 24811 17289 24820 17323
rect 24768 17280 24820 17289
rect 11428 17212 11480 17264
rect 13452 17212 13504 17264
rect 8300 17144 8352 17196
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 12532 17144 12584 17196
rect 13360 17144 13412 17196
rect 14648 17187 14700 17196
rect 14648 17153 14657 17187
rect 14657 17153 14691 17187
rect 14691 17153 14700 17187
rect 14648 17144 14700 17153
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 10876 17076 10928 17128
rect 13084 17076 13136 17128
rect 14004 17076 14056 17128
rect 10600 17051 10652 17060
rect 10600 17017 10609 17051
rect 10609 17017 10643 17051
rect 10643 17017 10652 17051
rect 11244 17051 11296 17060
rect 10600 17008 10652 17017
rect 11244 17017 11253 17051
rect 11253 17017 11287 17051
rect 11287 17017 11296 17051
rect 11244 17008 11296 17017
rect 2044 16983 2096 16992
rect 2044 16949 2053 16983
rect 2053 16949 2087 16983
rect 2087 16949 2096 16983
rect 2044 16940 2096 16949
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 9312 16940 9364 16992
rect 10876 16940 10928 16992
rect 11980 16940 12032 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 13820 16940 13872 16992
rect 23388 17076 23440 17128
rect 14832 17008 14884 17060
rect 15476 16940 15528 16992
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 9312 16779 9364 16788
rect 9312 16745 9321 16779
rect 9321 16745 9355 16779
rect 9355 16745 9364 16779
rect 9312 16736 9364 16745
rect 11336 16736 11388 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12532 16779 12584 16788
rect 12532 16745 12541 16779
rect 12541 16745 12575 16779
rect 12575 16745 12584 16779
rect 12532 16736 12584 16745
rect 13544 16779 13596 16788
rect 13544 16745 13553 16779
rect 13553 16745 13587 16779
rect 13587 16745 13596 16779
rect 13544 16736 13596 16745
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 14648 16736 14700 16788
rect 10692 16668 10744 16720
rect 10876 16668 10928 16720
rect 12900 16711 12952 16720
rect 12900 16677 12909 16711
rect 12909 16677 12943 16711
rect 12943 16677 12952 16711
rect 12900 16668 12952 16677
rect 13084 16668 13136 16720
rect 14004 16711 14056 16720
rect 14004 16677 14013 16711
rect 14013 16677 14047 16711
rect 14047 16677 14056 16711
rect 14004 16668 14056 16677
rect 1492 16600 1544 16652
rect 11336 16600 11388 16652
rect 24400 16736 24452 16788
rect 24768 16779 24820 16788
rect 24768 16745 24777 16779
rect 24777 16745 24811 16779
rect 24811 16745 24820 16779
rect 24768 16736 24820 16745
rect 13360 16532 13412 16584
rect 23848 16600 23900 16652
rect 24124 16600 24176 16652
rect 14648 16532 14700 16584
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 9404 16396 9456 16448
rect 13636 16439 13688 16448
rect 13636 16405 13645 16439
rect 13645 16405 13679 16439
rect 13679 16405 13688 16439
rect 13636 16396 13688 16405
rect 15476 16396 15528 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2320 16192 2372 16244
rect 9312 16192 9364 16244
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 11428 16235 11480 16244
rect 11428 16201 11437 16235
rect 11437 16201 11471 16235
rect 11471 16201 11480 16235
rect 11428 16192 11480 16201
rect 13360 16192 13412 16244
rect 14004 16192 14056 16244
rect 24124 16192 24176 16244
rect 2964 16056 3016 16108
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 23848 16167 23900 16176
rect 23848 16133 23857 16167
rect 23857 16133 23891 16167
rect 23891 16133 23900 16167
rect 23848 16124 23900 16133
rect 13636 16056 13688 16108
rect 1492 15920 1544 15972
rect 9404 15988 9456 16040
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 2688 15920 2740 15972
rect 2780 15920 2832 15972
rect 7564 15920 7616 15972
rect 10876 15920 10928 15972
rect 14648 15920 14700 15972
rect 15476 15988 15528 16040
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 1860 15852 1912 15904
rect 8576 15895 8628 15904
rect 8576 15861 8585 15895
rect 8585 15861 8619 15895
rect 8619 15861 8628 15895
rect 8576 15852 8628 15861
rect 9680 15852 9732 15904
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 14556 15852 14608 15904
rect 15292 15920 15344 15972
rect 15936 15852 15988 15904
rect 17776 15852 17828 15904
rect 23020 15852 23072 15904
rect 24952 15852 25004 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1400 15648 1452 15700
rect 8392 15648 8444 15700
rect 9220 15648 9272 15700
rect 10692 15648 10744 15700
rect 11428 15648 11480 15700
rect 13636 15648 13688 15700
rect 13728 15648 13780 15700
rect 15660 15691 15712 15700
rect 15660 15657 15669 15691
rect 15669 15657 15703 15691
rect 15703 15657 15712 15691
rect 15660 15648 15712 15657
rect 16028 15648 16080 15700
rect 24676 15648 24728 15700
rect 1676 15512 1728 15564
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 2688 15444 2740 15496
rect 6736 15444 6788 15496
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 10324 15512 10376 15564
rect 13820 15580 13872 15632
rect 14832 15580 14884 15632
rect 15844 15580 15896 15632
rect 11428 15512 11480 15564
rect 12992 15512 13044 15564
rect 8484 15444 8536 15496
rect 15476 15512 15528 15564
rect 17316 15512 17368 15564
rect 18236 15512 18288 15564
rect 19340 15512 19392 15564
rect 23572 15555 23624 15564
rect 23572 15521 23581 15555
rect 23581 15521 23615 15555
rect 23615 15521 23624 15555
rect 23572 15512 23624 15521
rect 23940 15512 23992 15564
rect 14648 15444 14700 15496
rect 22284 15444 22336 15496
rect 8668 15376 8720 15428
rect 13636 15419 13688 15428
rect 13636 15385 13645 15419
rect 13645 15385 13679 15419
rect 13679 15385 13688 15419
rect 13636 15376 13688 15385
rect 2688 15308 2740 15360
rect 4252 15351 4304 15360
rect 4252 15317 4261 15351
rect 4261 15317 4295 15351
rect 4295 15317 4304 15351
rect 4252 15308 4304 15317
rect 9588 15308 9640 15360
rect 11704 15308 11756 15360
rect 16488 15308 16540 15360
rect 16764 15351 16816 15360
rect 16764 15317 16773 15351
rect 16773 15317 16807 15351
rect 16807 15317 16816 15351
rect 16764 15308 16816 15317
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 17040 15308 17092 15317
rect 18328 15308 18380 15360
rect 19432 15308 19484 15360
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 2688 15104 2740 15156
rect 2780 15147 2832 15156
rect 2780 15113 2789 15147
rect 2789 15113 2823 15147
rect 2823 15113 2832 15147
rect 2780 15104 2832 15113
rect 7104 15147 7156 15156
rect 7104 15113 7113 15147
rect 7113 15113 7147 15147
rect 7147 15113 7156 15147
rect 7104 15104 7156 15113
rect 8208 15104 8260 15156
rect 9772 15104 9824 15156
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 10876 15104 10928 15156
rect 12992 15147 13044 15156
rect 12992 15113 13001 15147
rect 13001 15113 13035 15147
rect 13035 15113 13044 15147
rect 12992 15104 13044 15113
rect 13820 15104 13872 15156
rect 16028 15104 16080 15156
rect 24768 15147 24820 15156
rect 24768 15113 24777 15147
rect 24777 15113 24811 15147
rect 24811 15113 24820 15147
rect 24768 15104 24820 15113
rect 10692 15036 10744 15088
rect 5724 14968 5776 15020
rect 6828 14968 6880 15020
rect 22928 15036 22980 15088
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 11612 14968 11664 15020
rect 16672 14968 16724 15020
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 3148 14764 3200 14816
rect 6736 14832 6788 14884
rect 7012 14832 7064 14884
rect 9496 14900 9548 14952
rect 12348 14900 12400 14952
rect 12992 14900 13044 14952
rect 8024 14832 8076 14884
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 8484 14764 8536 14816
rect 9864 14764 9916 14816
rect 11336 14764 11388 14816
rect 11428 14764 11480 14816
rect 12348 14764 12400 14816
rect 13452 14764 13504 14816
rect 14556 14900 14608 14952
rect 16304 14900 16356 14952
rect 18512 14900 18564 14952
rect 19340 14900 19392 14952
rect 24400 14943 24452 14952
rect 13912 14832 13964 14884
rect 15936 14832 15988 14884
rect 17224 14832 17276 14884
rect 18788 14832 18840 14884
rect 13820 14764 13872 14816
rect 16396 14764 16448 14816
rect 17316 14807 17368 14816
rect 17316 14773 17325 14807
rect 17325 14773 17359 14807
rect 17359 14773 17368 14807
rect 17316 14764 17368 14773
rect 17408 14764 17460 14816
rect 18236 14764 18288 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 20168 14764 20220 14816
rect 24400 14909 24409 14943
rect 24409 14909 24443 14943
rect 24443 14909 24452 14943
rect 24400 14900 24452 14909
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 23204 14764 23256 14816
rect 23572 14764 23624 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 2596 14560 2648 14612
rect 4252 14560 4304 14612
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 8392 14603 8444 14612
rect 8392 14569 8401 14603
rect 8401 14569 8435 14603
rect 8435 14569 8444 14603
rect 8392 14560 8444 14569
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 11612 14603 11664 14612
rect 11612 14569 11621 14603
rect 11621 14569 11655 14603
rect 11655 14569 11664 14603
rect 11612 14560 11664 14569
rect 13728 14560 13780 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 17316 14560 17368 14612
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 22744 14560 22796 14612
rect 24124 14560 24176 14612
rect 2412 14424 2464 14476
rect 2320 14356 2372 14408
rect 2596 14288 2648 14340
rect 5724 14492 5776 14544
rect 15660 14535 15712 14544
rect 15660 14501 15669 14535
rect 15669 14501 15703 14535
rect 15703 14501 15712 14535
rect 15660 14492 15712 14501
rect 15752 14535 15804 14544
rect 15752 14501 15761 14535
rect 15761 14501 15795 14535
rect 15795 14501 15804 14535
rect 16304 14535 16356 14544
rect 15752 14492 15804 14501
rect 16304 14501 16313 14535
rect 16313 14501 16347 14535
rect 16347 14501 16356 14535
rect 16304 14492 16356 14501
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 9772 14424 9824 14476
rect 9956 14467 10008 14476
rect 9956 14433 9990 14467
rect 9990 14433 10008 14467
rect 9956 14424 10008 14433
rect 11980 14424 12032 14476
rect 14648 14424 14700 14476
rect 16120 14424 16172 14476
rect 19064 14424 19116 14476
rect 19524 14467 19576 14476
rect 19524 14433 19533 14467
rect 19533 14433 19567 14467
rect 19567 14433 19576 14467
rect 19524 14424 19576 14433
rect 21456 14424 21508 14476
rect 21548 14424 21600 14476
rect 22560 14467 22612 14476
rect 22560 14433 22569 14467
rect 22569 14433 22603 14467
rect 22603 14433 22612 14467
rect 22560 14424 22612 14433
rect 24124 14424 24176 14476
rect 24676 14424 24728 14476
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 4160 14288 4212 14340
rect 12440 14356 12492 14408
rect 12992 14356 13044 14408
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 17316 14399 17368 14408
rect 3424 14263 3476 14272
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 15844 14288 15896 14340
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 16856 14331 16908 14340
rect 16856 14297 16865 14331
rect 16865 14297 16899 14331
rect 16899 14297 16908 14331
rect 16856 14288 16908 14297
rect 6000 14220 6052 14272
rect 7472 14220 7524 14272
rect 11428 14220 11480 14272
rect 11704 14220 11756 14272
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 17868 14220 17920 14272
rect 18420 14220 18472 14272
rect 20536 14220 20588 14272
rect 21732 14220 21784 14272
rect 22376 14220 22428 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1952 14016 2004 14068
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 4436 14016 4488 14068
rect 5540 14016 5592 14068
rect 8024 14016 8076 14068
rect 8576 14016 8628 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 10784 14016 10836 14068
rect 11704 14059 11756 14068
rect 11704 14025 11713 14059
rect 11713 14025 11747 14059
rect 11747 14025 11756 14059
rect 11704 14016 11756 14025
rect 12992 14059 13044 14068
rect 12992 14025 13001 14059
rect 13001 14025 13035 14059
rect 13035 14025 13044 14059
rect 12992 14016 13044 14025
rect 15936 14016 15988 14068
rect 17316 14059 17368 14068
rect 17316 14025 17325 14059
rect 17325 14025 17359 14059
rect 17359 14025 17368 14059
rect 17316 14016 17368 14025
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 22560 14016 22612 14068
rect 2228 13948 2280 14000
rect 4160 13991 4212 14000
rect 4160 13957 4169 13991
rect 4169 13957 4203 13991
rect 4203 13957 4212 13991
rect 4160 13948 4212 13957
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 3240 13880 3292 13932
rect 6000 13948 6052 14000
rect 7012 13948 7064 14000
rect 10692 13948 10744 14000
rect 16120 13991 16172 14000
rect 16120 13957 16129 13991
rect 16129 13957 16163 13991
rect 16163 13957 16172 13991
rect 16120 13948 16172 13957
rect 16304 13991 16356 14000
rect 16304 13957 16313 13991
rect 16313 13957 16347 13991
rect 16347 13957 16356 13991
rect 16304 13948 16356 13957
rect 17868 13948 17920 14000
rect 15108 13880 15160 13932
rect 15660 13880 15712 13932
rect 16764 13923 16816 13932
rect 16764 13889 16773 13923
rect 16773 13889 16807 13923
rect 16807 13889 16816 13923
rect 16764 13880 16816 13889
rect 17500 13880 17552 13932
rect 22100 13948 22152 14000
rect 24768 13991 24820 14000
rect 24768 13957 24777 13991
rect 24777 13957 24811 13991
rect 24811 13957 24820 13991
rect 24768 13948 24820 13957
rect 4528 13855 4580 13864
rect 3792 13744 3844 13796
rect 4528 13821 4551 13855
rect 4551 13821 4580 13855
rect 4528 13812 4580 13821
rect 5632 13744 5684 13796
rect 7472 13744 7524 13796
rect 8116 13744 8168 13796
rect 9956 13812 10008 13864
rect 11704 13812 11756 13864
rect 11980 13812 12032 13864
rect 10784 13744 10836 13796
rect 13820 13855 13872 13864
rect 13820 13821 13854 13855
rect 13854 13821 13872 13855
rect 13820 13812 13872 13821
rect 14740 13812 14792 13864
rect 17592 13812 17644 13864
rect 19248 13880 19300 13932
rect 19524 13880 19576 13932
rect 23848 13880 23900 13932
rect 19616 13855 19668 13864
rect 19616 13821 19625 13855
rect 19625 13821 19659 13855
rect 19659 13821 19668 13855
rect 19616 13812 19668 13821
rect 20904 13855 20956 13864
rect 20904 13821 20913 13855
rect 20913 13821 20947 13855
rect 20947 13821 20956 13855
rect 20904 13812 20956 13821
rect 23296 13812 23348 13864
rect 24124 13812 24176 13864
rect 16304 13744 16356 13796
rect 12440 13676 12492 13728
rect 13452 13719 13504 13728
rect 13452 13685 13461 13719
rect 13461 13685 13495 13719
rect 13495 13685 13504 13719
rect 13452 13676 13504 13685
rect 14832 13676 14884 13728
rect 18052 13719 18104 13728
rect 18052 13685 18061 13719
rect 18061 13685 18095 13719
rect 18095 13685 18104 13719
rect 18052 13676 18104 13685
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 22468 13676 22520 13728
rect 24400 13719 24452 13728
rect 24400 13685 24409 13719
rect 24409 13685 24443 13719
rect 24443 13685 24452 13719
rect 24400 13676 24452 13685
rect 24676 13676 24728 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2504 13472 2556 13524
rect 2688 13515 2740 13524
rect 2688 13481 2697 13515
rect 2697 13481 2731 13515
rect 2731 13481 2740 13515
rect 2688 13472 2740 13481
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 11520 13472 11572 13524
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 15108 13515 15160 13524
rect 15108 13481 15117 13515
rect 15117 13481 15151 13515
rect 15151 13481 15160 13515
rect 15108 13472 15160 13481
rect 15752 13472 15804 13524
rect 17868 13472 17920 13524
rect 18236 13472 18288 13524
rect 18512 13472 18564 13524
rect 20076 13515 20128 13524
rect 20076 13481 20085 13515
rect 20085 13481 20119 13515
rect 20119 13481 20128 13515
rect 20076 13472 20128 13481
rect 24400 13472 24452 13524
rect 24768 13515 24820 13524
rect 24768 13481 24777 13515
rect 24777 13481 24811 13515
rect 24811 13481 24820 13515
rect 24768 13472 24820 13481
rect 7472 13404 7524 13456
rect 8024 13447 8076 13456
rect 8024 13413 8033 13447
rect 8033 13413 8067 13447
rect 8067 13413 8076 13447
rect 8024 13404 8076 13413
rect 13820 13404 13872 13456
rect 14648 13447 14700 13456
rect 14648 13413 14657 13447
rect 14657 13413 14691 13447
rect 14691 13413 14700 13447
rect 14648 13404 14700 13413
rect 1952 13336 2004 13388
rect 2228 13336 2280 13388
rect 4160 13336 4212 13388
rect 4528 13379 4580 13388
rect 4528 13345 4562 13379
rect 4562 13345 4580 13379
rect 4528 13336 4580 13345
rect 8208 13336 8260 13388
rect 10784 13336 10836 13388
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 14004 13379 14056 13388
rect 14004 13345 14013 13379
rect 14013 13345 14047 13379
rect 14047 13345 14056 13379
rect 14004 13336 14056 13345
rect 14556 13336 14608 13388
rect 16948 13336 17000 13388
rect 18972 13336 19024 13388
rect 23480 13336 23532 13388
rect 24676 13336 24728 13388
rect 2688 13268 2740 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 8576 13268 8628 13320
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 11796 13268 11848 13320
rect 14832 13268 14884 13320
rect 15844 13268 15896 13320
rect 18604 13268 18656 13320
rect 1400 13200 1452 13252
rect 9956 13200 10008 13252
rect 15752 13200 15804 13252
rect 3516 13175 3568 13184
rect 3516 13141 3525 13175
rect 3525 13141 3559 13175
rect 3559 13141 3568 13175
rect 3516 13132 3568 13141
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 17500 13132 17552 13184
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 21180 13268 21232 13320
rect 22560 13311 22612 13320
rect 22560 13277 22569 13311
rect 22569 13277 22603 13311
rect 22603 13277 22612 13311
rect 22560 13268 22612 13277
rect 18512 13132 18564 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 4252 12971 4304 12980
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 7748 12928 7800 12980
rect 8024 12928 8076 12980
rect 8208 12971 8260 12980
rect 8208 12937 8217 12971
rect 8217 12937 8251 12971
rect 8251 12937 8260 12971
rect 8208 12928 8260 12937
rect 11520 12928 11572 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 14004 12928 14056 12980
rect 15752 12928 15804 12980
rect 16304 12971 16356 12980
rect 16304 12937 16313 12971
rect 16313 12937 16347 12971
rect 16347 12937 16356 12971
rect 16304 12928 16356 12937
rect 23480 12928 23532 12980
rect 23940 12928 23992 12980
rect 3516 12792 3568 12844
rect 8116 12860 8168 12912
rect 10784 12903 10836 12912
rect 10784 12869 10793 12903
rect 10793 12869 10827 12903
rect 10827 12869 10836 12903
rect 10784 12860 10836 12869
rect 11336 12860 11388 12912
rect 1860 12724 1912 12776
rect 3792 12792 3844 12844
rect 4528 12792 4580 12844
rect 5172 12792 5224 12844
rect 8392 12792 8444 12844
rect 8668 12792 8720 12844
rect 9864 12792 9916 12844
rect 12348 12792 12400 12844
rect 13912 12792 13964 12844
rect 14832 12792 14884 12844
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 5080 12767 5132 12776
rect 4620 12724 4672 12733
rect 5080 12733 5089 12767
rect 5089 12733 5123 12767
rect 5123 12733 5132 12767
rect 5080 12724 5132 12733
rect 8576 12767 8628 12776
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 10692 12724 10744 12776
rect 3424 12656 3476 12708
rect 4252 12656 4304 12708
rect 4804 12656 4856 12708
rect 8760 12656 8812 12708
rect 11612 12656 11664 12708
rect 13084 12724 13136 12776
rect 13636 12724 13688 12776
rect 14096 12724 14148 12776
rect 16488 12724 16540 12776
rect 16580 12724 16632 12776
rect 17408 12724 17460 12776
rect 18512 12792 18564 12844
rect 20076 12835 20128 12844
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 20076 12792 20128 12801
rect 20260 12724 20312 12776
rect 12624 12656 12676 12708
rect 13360 12656 13412 12708
rect 15292 12656 15344 12708
rect 18512 12699 18564 12708
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 19524 12699 19576 12708
rect 18512 12656 18564 12665
rect 2964 12588 3016 12640
rect 9956 12588 10008 12640
rect 10692 12588 10744 12640
rect 11244 12588 11296 12640
rect 12256 12631 12308 12640
rect 12256 12597 12265 12631
rect 12265 12597 12299 12631
rect 12299 12597 12308 12631
rect 12256 12588 12308 12597
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 15384 12588 15436 12640
rect 15844 12631 15896 12640
rect 15844 12597 15853 12631
rect 15853 12597 15887 12631
rect 15887 12597 15896 12631
rect 15844 12588 15896 12597
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 19524 12665 19533 12699
rect 19533 12665 19567 12699
rect 19567 12665 19576 12699
rect 24676 12860 24728 12912
rect 24676 12724 24728 12776
rect 19524 12656 19576 12665
rect 21364 12588 21416 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2320 12384 2372 12436
rect 2596 12384 2648 12436
rect 4436 12384 4488 12436
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 13912 12384 13964 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 16028 12384 16080 12436
rect 16580 12427 16632 12436
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 18052 12384 18104 12436
rect 18696 12384 18748 12436
rect 20260 12427 20312 12436
rect 20260 12393 20269 12427
rect 20269 12393 20303 12427
rect 20303 12393 20312 12427
rect 20260 12384 20312 12393
rect 24032 12384 24084 12436
rect 2872 12316 2924 12368
rect 3332 12316 3384 12368
rect 6184 12316 6236 12368
rect 11520 12316 11572 12368
rect 2688 12248 2740 12300
rect 3424 12248 3476 12300
rect 6092 12248 6144 12300
rect 6368 12248 6420 12300
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 5080 12223 5132 12232
rect 2964 12180 3016 12189
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 3332 12112 3384 12164
rect 4252 12112 4304 12164
rect 7932 12180 7984 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 9680 12180 9732 12232
rect 12072 12248 12124 12300
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 13820 12316 13872 12368
rect 18880 12316 18932 12368
rect 19248 12316 19300 12368
rect 14188 12248 14240 12300
rect 17500 12248 17552 12300
rect 19064 12291 19116 12300
rect 19064 12257 19073 12291
rect 19073 12257 19107 12291
rect 19107 12257 19116 12291
rect 19064 12248 19116 12257
rect 20720 12248 20772 12300
rect 22284 12316 22336 12368
rect 22008 12248 22060 12300
rect 24216 12248 24268 12300
rect 13084 12180 13136 12232
rect 7472 12112 7524 12164
rect 9864 12155 9916 12164
rect 9864 12121 9873 12155
rect 9873 12121 9907 12155
rect 9907 12121 9916 12155
rect 9864 12112 9916 12121
rect 11520 12112 11572 12164
rect 13912 12180 13964 12232
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 15844 12180 15896 12232
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 16764 12180 16816 12189
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 3240 12044 3292 12096
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 6276 12087 6328 12096
rect 6276 12053 6285 12087
rect 6285 12053 6319 12087
rect 6319 12053 6328 12087
rect 6276 12044 6328 12053
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 17960 12044 18012 12096
rect 18604 12044 18656 12096
rect 21272 12180 21324 12232
rect 19064 12044 19116 12096
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 20996 12044 21048 12096
rect 21916 12044 21968 12096
rect 23940 12087 23992 12096
rect 23940 12053 23949 12087
rect 23949 12053 23983 12087
rect 23983 12053 23992 12087
rect 23940 12044 23992 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2872 11840 2924 11892
rect 3424 11840 3476 11892
rect 5080 11840 5132 11892
rect 7012 11840 7064 11892
rect 2320 11704 2372 11756
rect 8392 11840 8444 11892
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 9680 11840 9732 11849
rect 10784 11883 10836 11892
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 9680 11704 9732 11756
rect 4344 11636 4396 11688
rect 7380 11636 7432 11688
rect 7840 11636 7892 11688
rect 10140 11636 10192 11688
rect 12348 11840 12400 11892
rect 13544 11840 13596 11892
rect 16120 11883 16172 11892
rect 16120 11849 16129 11883
rect 16129 11849 16163 11883
rect 16163 11849 16172 11883
rect 16120 11840 16172 11849
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 21732 11840 21784 11892
rect 22008 11840 22060 11892
rect 22284 11840 22336 11892
rect 24032 11840 24084 11892
rect 14740 11772 14792 11824
rect 19064 11772 19116 11824
rect 20996 11772 21048 11824
rect 16028 11704 16080 11756
rect 12532 11636 12584 11688
rect 13452 11636 13504 11688
rect 13912 11679 13964 11688
rect 13912 11645 13946 11679
rect 13946 11645 13964 11679
rect 3976 11568 4028 11620
rect 6092 11568 6144 11620
rect 11520 11568 11572 11620
rect 11980 11568 12032 11620
rect 13912 11636 13964 11645
rect 14648 11636 14700 11688
rect 17960 11704 18012 11756
rect 17868 11636 17920 11688
rect 20720 11636 20772 11688
rect 14280 11568 14332 11620
rect 19524 11568 19576 11620
rect 20352 11568 20404 11620
rect 23940 11611 23992 11620
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 2320 11500 2372 11552
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 8300 11500 8352 11552
rect 9956 11543 10008 11552
rect 9956 11509 9965 11543
rect 9965 11509 9999 11543
rect 9999 11509 10008 11543
rect 9956 11500 10008 11509
rect 10048 11500 10100 11552
rect 12440 11500 12492 11552
rect 12624 11500 12676 11552
rect 14096 11500 14148 11552
rect 15016 11543 15068 11552
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 15476 11500 15528 11552
rect 16396 11500 16448 11552
rect 16764 11500 16816 11552
rect 17868 11500 17920 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 20076 11500 20128 11552
rect 20812 11500 20864 11552
rect 21088 11500 21140 11552
rect 21824 11543 21876 11552
rect 21824 11509 21833 11543
rect 21833 11509 21867 11543
rect 21867 11509 21876 11543
rect 21824 11500 21876 11509
rect 22284 11543 22336 11552
rect 22284 11509 22293 11543
rect 22293 11509 22327 11543
rect 22327 11509 22336 11543
rect 22284 11500 22336 11509
rect 23480 11500 23532 11552
rect 23940 11577 23974 11611
rect 23974 11577 23992 11611
rect 23940 11568 23992 11577
rect 24032 11568 24084 11620
rect 24584 11500 24636 11552
rect 25044 11543 25096 11552
rect 25044 11509 25053 11543
rect 25053 11509 25087 11543
rect 25087 11509 25096 11543
rect 25044 11500 25096 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2228 11296 2280 11348
rect 2688 11296 2740 11348
rect 2780 11296 2832 11348
rect 4344 11296 4396 11348
rect 6644 11296 6696 11348
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 13084 11339 13136 11348
rect 13084 11305 13093 11339
rect 13093 11305 13127 11339
rect 13127 11305 13136 11339
rect 13084 11296 13136 11305
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 14648 11339 14700 11348
rect 13176 11296 13228 11305
rect 14648 11305 14657 11339
rect 14657 11305 14691 11339
rect 14691 11305 14700 11339
rect 14648 11296 14700 11305
rect 16488 11296 16540 11348
rect 16856 11296 16908 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 21088 11296 21140 11348
rect 22560 11296 22612 11348
rect 2872 11228 2924 11280
rect 6276 11228 6328 11280
rect 7012 11228 7064 11280
rect 7656 11271 7708 11280
rect 7656 11237 7665 11271
rect 7665 11237 7699 11271
rect 7699 11237 7708 11271
rect 7656 11228 7708 11237
rect 8024 11228 8076 11280
rect 8392 11228 8444 11280
rect 11612 11228 11664 11280
rect 12440 11228 12492 11280
rect 18512 11228 18564 11280
rect 18972 11228 19024 11280
rect 20444 11228 20496 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 3608 11160 3660 11212
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 6552 11160 6604 11212
rect 7564 11160 7616 11212
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 10968 11203 11020 11212
rect 10968 11169 11002 11203
rect 11002 11169 11020 11203
rect 10968 11160 11020 11169
rect 2320 11092 2372 11144
rect 4620 11135 4672 11144
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 2596 11024 2648 11076
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 6184 11092 6236 11144
rect 6460 11092 6512 11144
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 2412 10956 2464 11008
rect 3148 11024 3200 11076
rect 3976 11024 4028 11076
rect 5540 11024 5592 11076
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 5080 10999 5132 11008
rect 5080 10965 5089 10999
rect 5089 10965 5123 10999
rect 5123 10965 5132 10999
rect 5080 10956 5132 10965
rect 6000 10956 6052 11008
rect 11336 10956 11388 11008
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 13176 11160 13228 11212
rect 13728 11160 13780 11212
rect 15016 11160 15068 11212
rect 16120 11160 16172 11212
rect 19616 11203 19668 11212
rect 19616 11169 19625 11203
rect 19625 11169 19659 11203
rect 19659 11169 19668 11203
rect 19616 11160 19668 11169
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 19984 11160 20036 11212
rect 13912 11092 13964 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 15292 11135 15344 11144
rect 14280 11092 14332 11101
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 18512 11092 18564 11144
rect 20076 11092 20128 11144
rect 20720 11092 20772 11144
rect 21916 11024 21968 11076
rect 22744 11228 22796 11280
rect 24860 11296 24912 11348
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 23480 11228 23532 11280
rect 22560 11160 22612 11212
rect 23572 11160 23624 11212
rect 23848 11160 23900 11212
rect 24584 11160 24636 11212
rect 24952 11203 25004 11212
rect 24952 11169 24961 11203
rect 24961 11169 24995 11203
rect 24995 11169 25004 11203
rect 24952 11160 25004 11169
rect 22744 11092 22796 11144
rect 23940 11135 23992 11144
rect 23940 11101 23949 11135
rect 23949 11101 23983 11135
rect 23983 11101 23992 11135
rect 23940 11092 23992 11101
rect 24216 11024 24268 11076
rect 16856 10956 16908 11008
rect 18604 10956 18656 11008
rect 19524 10956 19576 11008
rect 20720 10956 20772 11008
rect 23388 10999 23440 11008
rect 23388 10965 23397 10999
rect 23397 10965 23431 10999
rect 23431 10965 23440 10999
rect 23388 10956 23440 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2136 10752 2188 10804
rect 4620 10795 4672 10804
rect 4620 10761 4629 10795
rect 4629 10761 4663 10795
rect 4663 10761 4672 10795
rect 4620 10752 4672 10761
rect 4896 10752 4948 10804
rect 7104 10752 7156 10804
rect 8024 10752 8076 10804
rect 10692 10752 10744 10804
rect 12532 10752 12584 10804
rect 13176 10752 13228 10804
rect 13912 10752 13964 10804
rect 15292 10752 15344 10804
rect 7196 10727 7248 10736
rect 7196 10693 7205 10727
rect 7205 10693 7239 10727
rect 7239 10693 7248 10727
rect 7196 10684 7248 10693
rect 9496 10684 9548 10736
rect 11612 10684 11664 10736
rect 12900 10684 12952 10736
rect 5080 10616 5132 10668
rect 6000 10616 6052 10668
rect 6460 10616 6512 10668
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 11428 10616 11480 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 16764 10752 16816 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 19248 10752 19300 10804
rect 19616 10752 19668 10804
rect 21456 10752 21508 10804
rect 22652 10795 22704 10804
rect 22652 10761 22661 10795
rect 22661 10761 22695 10795
rect 22695 10761 22704 10795
rect 22652 10752 22704 10761
rect 24952 10795 25004 10804
rect 24952 10761 24961 10795
rect 24961 10761 24995 10795
rect 24995 10761 25004 10795
rect 24952 10752 25004 10761
rect 25504 10752 25556 10804
rect 12256 10616 12308 10625
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 21916 10684 21968 10736
rect 23664 10684 23716 10736
rect 4436 10548 4488 10600
rect 8208 10548 8260 10600
rect 3424 10480 3476 10532
rect 5356 10480 5408 10532
rect 6184 10523 6236 10532
rect 6184 10489 6193 10523
rect 6193 10489 6227 10523
rect 6227 10489 6236 10523
rect 6184 10480 6236 10489
rect 8116 10480 8168 10532
rect 1676 10412 1728 10464
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 9680 10412 9732 10464
rect 11152 10480 11204 10532
rect 12532 10548 12584 10600
rect 12716 10548 12768 10600
rect 15752 10591 15804 10600
rect 15752 10557 15786 10591
rect 15786 10557 15804 10591
rect 15752 10548 15804 10557
rect 16488 10548 16540 10600
rect 18144 10591 18196 10600
rect 18144 10557 18153 10591
rect 18153 10557 18187 10591
rect 18187 10557 18196 10591
rect 18144 10548 18196 10557
rect 20720 10548 20772 10600
rect 22192 10548 22244 10600
rect 23480 10548 23532 10600
rect 25044 10616 25096 10668
rect 24676 10548 24728 10600
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25228 10548 25280 10557
rect 20628 10480 20680 10532
rect 21824 10480 21876 10532
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 12532 10412 12584 10464
rect 13728 10412 13780 10464
rect 14372 10412 14424 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 17408 10455 17460 10464
rect 14464 10412 14516 10421
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 17868 10455 17920 10464
rect 17868 10421 17877 10455
rect 17877 10421 17911 10455
rect 17911 10421 17920 10455
rect 17868 10412 17920 10421
rect 18144 10412 18196 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 22008 10455 22060 10464
rect 22008 10421 22017 10455
rect 22017 10421 22051 10455
rect 22051 10421 22060 10455
rect 22008 10412 22060 10421
rect 22468 10412 22520 10464
rect 22652 10412 22704 10464
rect 23664 10455 23716 10464
rect 23664 10421 23673 10455
rect 23673 10421 23707 10455
rect 23707 10421 23716 10455
rect 23664 10412 23716 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10208 1912 10260
rect 2320 10208 2372 10260
rect 2596 10208 2648 10260
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 7380 10208 7432 10260
rect 8300 10208 8352 10260
rect 8484 10208 8536 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 10692 10208 10744 10260
rect 10968 10251 11020 10260
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 16120 10251 16172 10260
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 17316 10208 17368 10260
rect 18236 10251 18288 10260
rect 18236 10217 18245 10251
rect 18245 10217 18279 10251
rect 18279 10217 18288 10251
rect 18236 10208 18288 10217
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 19340 10208 19392 10260
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 20720 10208 20772 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 22284 10208 22336 10260
rect 23388 10208 23440 10260
rect 25044 10208 25096 10260
rect 2504 10140 2556 10192
rect 6276 10140 6328 10192
rect 12256 10140 12308 10192
rect 13544 10140 13596 10192
rect 17776 10140 17828 10192
rect 1584 10072 1636 10124
rect 3884 10072 3936 10124
rect 4160 10072 4212 10124
rect 6460 10072 6512 10124
rect 7932 10115 7984 10124
rect 7932 10081 7941 10115
rect 7941 10081 7975 10115
rect 7975 10081 7984 10115
rect 7932 10072 7984 10081
rect 8116 10072 8168 10124
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 11060 10072 11112 10124
rect 16948 10072 17000 10124
rect 19984 10140 20036 10192
rect 22744 10183 22796 10192
rect 22744 10149 22753 10183
rect 22753 10149 22787 10183
rect 22787 10149 22796 10183
rect 22744 10140 22796 10149
rect 23572 10140 23624 10192
rect 19800 10115 19852 10124
rect 19800 10081 19809 10115
rect 19809 10081 19843 10115
rect 19843 10081 19852 10115
rect 19800 10072 19852 10081
rect 21824 10072 21876 10124
rect 23020 10072 23072 10124
rect 2596 10004 2648 10056
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 2964 10004 3016 10056
rect 3608 10004 3660 10056
rect 4436 10004 4488 10056
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 13360 10047 13412 10056
rect 3424 9936 3476 9988
rect 7104 9979 7156 9988
rect 2320 9911 2372 9920
rect 2320 9877 2329 9911
rect 2329 9877 2363 9911
rect 2363 9877 2372 9911
rect 2320 9868 2372 9877
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 7104 9945 7113 9979
rect 7113 9945 7147 9979
rect 7147 9945 7156 9979
rect 7104 9936 7156 9945
rect 8944 9979 8996 9988
rect 8944 9945 8953 9979
rect 8953 9945 8987 9979
rect 8987 9945 8996 9979
rect 8944 9936 8996 9945
rect 10968 9936 11020 9988
rect 11152 9979 11204 9988
rect 11152 9945 11161 9979
rect 11161 9945 11195 9979
rect 11195 9945 11204 9979
rect 11152 9936 11204 9945
rect 11520 9936 11572 9988
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 14832 10004 14884 10056
rect 17408 10004 17460 10056
rect 19524 10004 19576 10056
rect 21088 10004 21140 10056
rect 19984 9979 20036 9988
rect 19984 9945 19993 9979
rect 19993 9945 20027 9979
rect 20027 9945 20036 9979
rect 19984 9936 20036 9945
rect 22008 10004 22060 10056
rect 23112 10004 23164 10056
rect 5172 9868 5224 9920
rect 6460 9911 6512 9920
rect 6460 9877 6469 9911
rect 6469 9877 6503 9911
rect 6503 9877 6512 9911
rect 6460 9868 6512 9877
rect 10600 9911 10652 9920
rect 10600 9877 10609 9911
rect 10609 9877 10643 9911
rect 10643 9877 10652 9911
rect 10600 9868 10652 9877
rect 12808 9868 12860 9920
rect 13728 9868 13780 9920
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 16580 9911 16632 9920
rect 16580 9877 16589 9911
rect 16589 9877 16623 9911
rect 16623 9877 16632 9911
rect 16580 9868 16632 9877
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 20076 9868 20128 9920
rect 20352 9868 20404 9920
rect 24676 9868 24728 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1584 9707 1636 9716
rect 1584 9673 1593 9707
rect 1593 9673 1627 9707
rect 1627 9673 1636 9707
rect 1584 9664 1636 9673
rect 2320 9664 2372 9716
rect 6000 9664 6052 9716
rect 9680 9664 9732 9716
rect 9864 9664 9916 9716
rect 10692 9664 10744 9716
rect 11060 9664 11112 9716
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 4160 9596 4212 9648
rect 4344 9639 4396 9648
rect 4344 9605 4353 9639
rect 4353 9605 4387 9639
rect 4387 9605 4396 9639
rect 4344 9596 4396 9605
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 9312 9639 9364 9648
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 2044 9367 2096 9376
rect 2044 9333 2053 9367
rect 2053 9333 2087 9367
rect 2087 9333 2096 9367
rect 2044 9324 2096 9333
rect 3240 9324 3292 9376
rect 3516 9324 3568 9376
rect 5172 9528 5224 9580
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 11336 9596 11388 9648
rect 12256 9596 12308 9648
rect 5448 9460 5500 9512
rect 7656 9460 7708 9512
rect 10692 9528 10744 9580
rect 11428 9528 11480 9580
rect 13360 9664 13412 9716
rect 13176 9596 13228 9648
rect 17316 9664 17368 9716
rect 9036 9460 9088 9512
rect 9864 9460 9916 9512
rect 10876 9460 10928 9512
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 8576 9392 8628 9444
rect 11336 9392 11388 9444
rect 12808 9435 12860 9444
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 4160 9324 4212 9376
rect 6000 9324 6052 9376
rect 6368 9324 6420 9376
rect 7012 9324 7064 9376
rect 7932 9324 7984 9376
rect 10784 9324 10836 9376
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 13728 9528 13780 9580
rect 14556 9528 14608 9580
rect 15016 9571 15068 9580
rect 15016 9537 15025 9571
rect 15025 9537 15059 9571
rect 15059 9537 15068 9571
rect 15016 9528 15068 9537
rect 14832 9503 14884 9512
rect 14832 9469 14841 9503
rect 14841 9469 14875 9503
rect 14875 9469 14884 9503
rect 14832 9460 14884 9469
rect 15660 9596 15712 9648
rect 16120 9528 16172 9580
rect 16488 9460 16540 9512
rect 17960 9460 18012 9512
rect 18236 9664 18288 9716
rect 19524 9664 19576 9716
rect 20352 9707 20404 9716
rect 20352 9673 20361 9707
rect 20361 9673 20395 9707
rect 20395 9673 20404 9707
rect 20352 9664 20404 9673
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 21272 9664 21324 9716
rect 23020 9664 23072 9716
rect 23204 9596 23256 9648
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 22284 9528 22336 9580
rect 23112 9528 23164 9580
rect 24676 9528 24728 9580
rect 18144 9460 18196 9512
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 20720 9460 20772 9512
rect 23664 9460 23716 9512
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 16304 9392 16356 9444
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 16120 9324 16172 9376
rect 16948 9324 17000 9376
rect 19248 9324 19300 9376
rect 20996 9324 21048 9376
rect 24952 9324 25004 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2504 9120 2556 9172
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 7104 9163 7156 9172
rect 2780 9120 2832 9129
rect 7104 9129 7113 9163
rect 7113 9129 7147 9163
rect 7147 9129 7156 9163
rect 7104 9120 7156 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 8024 9120 8076 9172
rect 8300 9120 8352 9172
rect 11428 9120 11480 9172
rect 14832 9120 14884 9172
rect 15016 9163 15068 9172
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 15292 9120 15344 9172
rect 17040 9120 17092 9172
rect 17408 9120 17460 9172
rect 2964 9052 3016 9104
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 2872 8984 2924 8993
rect 4160 8984 4212 9036
rect 4344 9027 4396 9036
rect 4344 8993 4378 9027
rect 4378 8993 4396 9027
rect 4344 8984 4396 8993
rect 10048 9052 10100 9104
rect 1952 8916 2004 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 6552 8916 6604 8968
rect 9312 8984 9364 9036
rect 10600 9027 10652 9036
rect 10600 8993 10634 9027
rect 10634 8993 10652 9027
rect 10600 8984 10652 8993
rect 10876 9052 10928 9104
rect 12256 8984 12308 9036
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 8576 8916 8628 8968
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 12164 8916 12216 8968
rect 13728 8984 13780 9036
rect 15476 9052 15528 9104
rect 15844 8984 15896 9036
rect 18604 9120 18656 9172
rect 21364 9163 21416 9172
rect 21364 9129 21373 9163
rect 21373 9129 21407 9163
rect 21407 9129 21416 9163
rect 21364 9120 21416 9129
rect 22376 9163 22428 9172
rect 22376 9129 22385 9163
rect 22385 9129 22419 9163
rect 22419 9129 22428 9163
rect 22376 9120 22428 9129
rect 22836 9163 22888 9172
rect 22836 9129 22845 9163
rect 22845 9129 22879 9163
rect 22879 9129 22888 9163
rect 22836 9120 22888 9129
rect 23112 9120 23164 9172
rect 23664 9163 23716 9172
rect 23664 9129 23673 9163
rect 23673 9129 23707 9163
rect 23707 9129 23716 9163
rect 23664 9120 23716 9129
rect 18512 9095 18564 9104
rect 18512 9061 18521 9095
rect 18521 9061 18555 9095
rect 18555 9061 18564 9095
rect 18512 9052 18564 9061
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 2596 8780 2648 8832
rect 3976 8848 4028 8900
rect 13084 8848 13136 8900
rect 14740 8916 14792 8968
rect 17868 8916 17920 8968
rect 18328 8916 18380 8968
rect 20168 9052 20220 9104
rect 21272 9095 21324 9104
rect 21272 9061 21281 9095
rect 21281 9061 21315 9095
rect 21315 9061 21324 9095
rect 21272 9052 21324 9061
rect 24952 9052 25004 9104
rect 19432 8984 19484 9036
rect 22652 9027 22704 9036
rect 22652 8993 22661 9027
rect 22661 8993 22695 9027
rect 22695 8993 22704 9027
rect 22652 8984 22704 8993
rect 23020 8984 23072 9036
rect 19248 8916 19300 8968
rect 21180 8916 21232 8968
rect 19524 8848 19576 8900
rect 4068 8780 4120 8832
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 6276 8780 6328 8832
rect 6736 8823 6788 8832
rect 6736 8789 6745 8823
rect 6745 8789 6779 8823
rect 6779 8789 6788 8823
rect 6736 8780 6788 8789
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 10140 8780 10192 8832
rect 10692 8780 10744 8832
rect 12348 8780 12400 8832
rect 13728 8780 13780 8832
rect 13820 8823 13872 8832
rect 13820 8789 13829 8823
rect 13829 8789 13863 8823
rect 13863 8789 13872 8823
rect 13820 8780 13872 8789
rect 18328 8780 18380 8832
rect 19984 8780 20036 8832
rect 20720 8823 20772 8832
rect 20720 8789 20729 8823
rect 20729 8789 20763 8823
rect 20763 8789 20772 8823
rect 20720 8780 20772 8789
rect 25136 8823 25188 8832
rect 25136 8789 25145 8823
rect 25145 8789 25179 8823
rect 25179 8789 25188 8823
rect 25136 8780 25188 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2504 8576 2556 8628
rect 4344 8576 4396 8628
rect 7564 8576 7616 8628
rect 3240 8508 3292 8560
rect 5448 8440 5500 8492
rect 6460 8440 6512 8492
rect 6736 8440 6788 8492
rect 10600 8576 10652 8628
rect 13084 8576 13136 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18236 8576 18288 8628
rect 20168 8619 20220 8628
rect 20168 8585 20177 8619
rect 20177 8585 20211 8619
rect 20211 8585 20220 8619
rect 20168 8576 20220 8585
rect 21364 8576 21416 8628
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 25136 8576 25188 8628
rect 25688 8619 25740 8628
rect 25688 8585 25697 8619
rect 25697 8585 25731 8619
rect 25731 8585 25740 8619
rect 25688 8576 25740 8585
rect 16120 8508 16172 8560
rect 22008 8551 22060 8560
rect 22008 8517 22017 8551
rect 22017 8517 22051 8551
rect 22051 8517 22060 8551
rect 22008 8508 22060 8517
rect 10324 8440 10376 8492
rect 11152 8440 11204 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 11520 8440 11572 8492
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 5264 8372 5316 8424
rect 8024 8372 8076 8424
rect 2320 8304 2372 8356
rect 4252 8347 4304 8356
rect 4252 8313 4261 8347
rect 4261 8313 4295 8347
rect 4295 8313 4304 8347
rect 4252 8304 4304 8313
rect 6552 8347 6604 8356
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 7104 8304 7156 8356
rect 8300 8304 8352 8356
rect 8576 8304 8628 8356
rect 9312 8372 9364 8424
rect 24216 8440 24268 8492
rect 24584 8483 24636 8492
rect 24584 8449 24593 8483
rect 24593 8449 24627 8483
rect 24627 8449 24636 8483
rect 24584 8440 24636 8449
rect 12348 8372 12400 8424
rect 12164 8347 12216 8356
rect 12164 8313 12173 8347
rect 12173 8313 12207 8347
rect 12207 8313 12216 8347
rect 12164 8304 12216 8313
rect 3056 8236 3108 8288
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 8116 8236 8168 8245
rect 12532 8372 12584 8424
rect 14740 8372 14792 8424
rect 17960 8372 18012 8424
rect 20628 8415 20680 8424
rect 20628 8381 20637 8415
rect 20637 8381 20671 8415
rect 20671 8381 20680 8415
rect 20628 8372 20680 8381
rect 25504 8415 25556 8424
rect 25504 8381 25513 8415
rect 25513 8381 25547 8415
rect 25547 8381 25556 8415
rect 25504 8372 25556 8381
rect 15292 8304 15344 8356
rect 16580 8304 16632 8356
rect 17868 8304 17920 8356
rect 18328 8347 18380 8356
rect 18328 8313 18362 8347
rect 18362 8313 18380 8347
rect 18328 8304 18380 8313
rect 19248 8304 19300 8356
rect 20720 8304 20772 8356
rect 22652 8347 22704 8356
rect 15476 8236 15528 8288
rect 22652 8313 22661 8347
rect 22661 8313 22695 8347
rect 22695 8313 22704 8347
rect 22652 8304 22704 8313
rect 23480 8347 23532 8356
rect 23480 8313 23489 8347
rect 23489 8313 23523 8347
rect 23523 8313 23532 8347
rect 23480 8304 23532 8313
rect 22284 8236 22336 8288
rect 23940 8279 23992 8288
rect 23940 8245 23949 8279
rect 23949 8245 23983 8279
rect 23983 8245 23992 8279
rect 23940 8236 23992 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 8032 1452 8084
rect 2872 8032 2924 8084
rect 4712 8032 4764 8084
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 7472 8032 7524 8084
rect 8760 8032 8812 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 13176 8075 13228 8084
rect 13176 8041 13185 8075
rect 13185 8041 13219 8075
rect 13219 8041 13228 8075
rect 13176 8032 13228 8041
rect 13268 8032 13320 8084
rect 13728 8032 13780 8084
rect 14740 8032 14792 8084
rect 16580 8032 16632 8084
rect 17040 8032 17092 8084
rect 17776 8032 17828 8084
rect 17960 8032 18012 8084
rect 18512 8032 18564 8084
rect 18788 8032 18840 8084
rect 19524 8032 19576 8084
rect 20628 8032 20680 8084
rect 20812 8032 20864 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 23940 8032 23992 8084
rect 2688 7964 2740 8016
rect 3056 7964 3108 8016
rect 8668 7964 8720 8016
rect 10140 8007 10192 8016
rect 10140 7973 10149 8007
rect 10149 7973 10183 8007
rect 10183 7973 10192 8007
rect 10140 7964 10192 7973
rect 11428 8007 11480 8016
rect 11428 7973 11462 8007
rect 11462 7973 11480 8007
rect 11428 7964 11480 7973
rect 24584 7964 24636 8016
rect 2596 7939 2648 7948
rect 2596 7905 2605 7939
rect 2605 7905 2639 7939
rect 2639 7905 2648 7939
rect 2596 7896 2648 7905
rect 4160 7896 4212 7948
rect 6184 7939 6236 7948
rect 6184 7905 6193 7939
rect 6193 7905 6227 7939
rect 6227 7905 6236 7939
rect 6184 7896 6236 7905
rect 6460 7896 6512 7948
rect 6644 7896 6696 7948
rect 8024 7939 8076 7948
rect 8024 7905 8033 7939
rect 8033 7905 8067 7939
rect 8067 7905 8076 7939
rect 8024 7896 8076 7905
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 4620 7871 4672 7880
rect 2320 7760 2372 7812
rect 2504 7760 2556 7812
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 3332 7760 3384 7812
rect 3884 7760 3936 7812
rect 7748 7828 7800 7880
rect 12624 7896 12676 7948
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 14556 7896 14608 7948
rect 16028 7896 16080 7948
rect 16672 7896 16724 7948
rect 17960 7896 18012 7948
rect 19248 7896 19300 7948
rect 21180 7939 21232 7948
rect 21180 7905 21214 7939
rect 21214 7905 21232 7939
rect 21180 7896 21232 7905
rect 11152 7871 11204 7880
rect 6920 7760 6972 7812
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 14188 7871 14240 7880
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 10140 7760 10192 7812
rect 18144 7828 18196 7880
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 19800 7871 19852 7880
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 20720 7828 20772 7880
rect 20812 7828 20864 7880
rect 18328 7760 18380 7812
rect 1400 7692 1452 7744
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 7656 7735 7708 7744
rect 7656 7701 7665 7735
rect 7665 7701 7699 7735
rect 7699 7701 7708 7735
rect 7656 7692 7708 7701
rect 9864 7735 9916 7744
rect 9864 7701 9873 7735
rect 9873 7701 9907 7735
rect 9907 7701 9916 7735
rect 9864 7692 9916 7701
rect 12992 7692 13044 7744
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 14740 7692 14792 7744
rect 22836 7735 22888 7744
rect 22836 7701 22845 7735
rect 22845 7701 22879 7735
rect 22879 7701 22888 7735
rect 22836 7692 22888 7701
rect 23480 7692 23532 7744
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2136 7488 2188 7540
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 4712 7488 4764 7540
rect 3976 7420 4028 7472
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 9680 7488 9732 7540
rect 11152 7488 11204 7540
rect 11428 7488 11480 7540
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 14188 7488 14240 7540
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 16672 7488 16724 7540
rect 17592 7488 17644 7540
rect 6460 7420 6512 7472
rect 8024 7420 8076 7472
rect 9312 7463 9364 7472
rect 9312 7429 9321 7463
rect 9321 7429 9355 7463
rect 9355 7429 9364 7463
rect 9312 7420 9364 7429
rect 5816 7352 5868 7361
rect 10140 7352 10192 7404
rect 13176 7352 13228 7404
rect 15476 7420 15528 7472
rect 16396 7420 16448 7472
rect 17040 7352 17092 7404
rect 19708 7488 19760 7540
rect 20260 7488 20312 7540
rect 20812 7488 20864 7540
rect 23572 7488 23624 7540
rect 25136 7531 25188 7540
rect 25136 7497 25145 7531
rect 25145 7497 25179 7531
rect 25179 7497 25188 7531
rect 25136 7488 25188 7497
rect 19800 7420 19852 7472
rect 23756 7420 23808 7472
rect 19248 7352 19300 7404
rect 21180 7352 21232 7404
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 6000 7284 6052 7336
rect 6184 7284 6236 7336
rect 3240 7216 3292 7268
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 5540 7148 5592 7200
rect 6920 7284 6972 7336
rect 9680 7284 9732 7336
rect 8300 7148 8352 7200
rect 9312 7148 9364 7200
rect 13084 7216 13136 7268
rect 14648 7284 14700 7336
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 16672 7327 16724 7336
rect 15844 7284 15896 7293
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 18052 7284 18104 7336
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 20168 7327 20220 7336
rect 20168 7293 20177 7327
rect 20177 7293 20211 7327
rect 20211 7293 20220 7327
rect 20168 7284 20220 7293
rect 16028 7216 16080 7268
rect 16212 7216 16264 7268
rect 18972 7216 19024 7268
rect 21272 7284 21324 7336
rect 23940 7352 23992 7404
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 25320 7352 25372 7404
rect 22100 7327 22152 7336
rect 22100 7293 22109 7327
rect 22109 7293 22143 7327
rect 22143 7293 22152 7327
rect 22100 7284 22152 7293
rect 22928 7284 22980 7336
rect 23112 7327 23164 7336
rect 23112 7293 23121 7327
rect 23121 7293 23155 7327
rect 23155 7293 23164 7327
rect 25228 7327 25280 7336
rect 23112 7284 23164 7293
rect 25228 7293 25237 7327
rect 25237 7293 25271 7327
rect 25271 7293 25280 7327
rect 25228 7284 25280 7293
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 17960 7148 18012 7200
rect 20352 7148 20404 7200
rect 23756 7216 23808 7268
rect 21364 7148 21416 7200
rect 23296 7148 23348 7200
rect 23572 7148 23624 7200
rect 25412 7191 25464 7200
rect 25412 7157 25421 7191
rect 25421 7157 25455 7191
rect 25455 7157 25464 7191
rect 25412 7148 25464 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 2596 6944 2648 6996
rect 3976 6944 4028 6996
rect 7012 6944 7064 6996
rect 10968 6944 11020 6996
rect 11612 6944 11664 6996
rect 12164 6987 12216 6996
rect 12164 6953 12173 6987
rect 12173 6953 12207 6987
rect 12207 6953 12216 6987
rect 12164 6944 12216 6953
rect 13360 6944 13412 6996
rect 18052 6987 18104 6996
rect 18052 6953 18061 6987
rect 18061 6953 18095 6987
rect 18095 6953 18104 6987
rect 18052 6944 18104 6953
rect 18880 6987 18932 6996
rect 18880 6953 18889 6987
rect 18889 6953 18923 6987
rect 18923 6953 18932 6987
rect 18880 6944 18932 6953
rect 20260 6987 20312 6996
rect 20260 6953 20269 6987
rect 20269 6953 20303 6987
rect 20303 6953 20312 6987
rect 20260 6944 20312 6953
rect 22100 6944 22152 6996
rect 22928 6944 22980 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 2136 6808 2188 6860
rect 5540 6808 5592 6860
rect 5816 6876 5868 6928
rect 6000 6876 6052 6928
rect 9864 6876 9916 6928
rect 2412 6740 2464 6792
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 3516 6740 3568 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 3240 6672 3292 6724
rect 1676 6604 1728 6656
rect 6920 6672 6972 6724
rect 8024 6808 8076 6860
rect 9680 6808 9732 6860
rect 11060 6851 11112 6860
rect 11060 6817 11094 6851
rect 11094 6817 11112 6851
rect 11060 6808 11112 6817
rect 12256 6808 12308 6860
rect 15108 6876 15160 6928
rect 19340 6876 19392 6928
rect 19616 6876 19668 6928
rect 24308 6876 24360 6928
rect 14004 6808 14056 6860
rect 14280 6808 14332 6860
rect 15568 6851 15620 6860
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 16120 6808 16172 6860
rect 18144 6808 18196 6860
rect 20076 6808 20128 6860
rect 20628 6808 20680 6860
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 4620 6604 4672 6613
rect 5080 6604 5132 6656
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 9496 6740 9548 6792
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 9128 6604 9180 6656
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 9680 6604 9732 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 13360 6740 13412 6792
rect 15844 6740 15896 6792
rect 18972 6783 19024 6792
rect 18972 6749 18981 6783
rect 18981 6749 19015 6783
rect 19015 6749 19024 6783
rect 18972 6740 19024 6749
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 20812 6740 20864 6792
rect 23572 6740 23624 6792
rect 14004 6672 14056 6724
rect 11152 6604 11204 6656
rect 13728 6604 13780 6656
rect 14096 6604 14148 6656
rect 16212 6604 16264 6656
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 17960 6604 18012 6656
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 22928 6647 22980 6656
rect 22928 6613 22937 6647
rect 22937 6613 22971 6647
rect 22971 6613 22980 6647
rect 22928 6604 22980 6613
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2136 6443 2188 6452
rect 2136 6409 2145 6443
rect 2145 6409 2179 6443
rect 2179 6409 2188 6443
rect 2136 6400 2188 6409
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 3148 6400 3200 6452
rect 5540 6400 5592 6452
rect 6920 6400 6972 6452
rect 9496 6443 9548 6452
rect 9496 6409 9505 6443
rect 9505 6409 9539 6443
rect 9539 6409 9548 6443
rect 9496 6400 9548 6409
rect 10692 6400 10744 6452
rect 12992 6400 13044 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 14648 6400 14700 6452
rect 17408 6400 17460 6452
rect 19064 6400 19116 6452
rect 2872 6332 2924 6384
rect 4160 6332 4212 6384
rect 5448 6375 5500 6384
rect 5448 6341 5457 6375
rect 5457 6341 5491 6375
rect 5491 6341 5500 6375
rect 5448 6332 5500 6341
rect 10508 6375 10560 6384
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 10508 6332 10560 6341
rect 11336 6332 11388 6384
rect 11612 6332 11664 6384
rect 3332 6264 3384 6316
rect 3516 6264 3568 6316
rect 5080 6307 5132 6316
rect 5080 6273 5089 6307
rect 5089 6273 5123 6307
rect 5123 6273 5132 6307
rect 5080 6264 5132 6273
rect 6184 6264 6236 6316
rect 10140 6264 10192 6316
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 7472 6196 7524 6248
rect 8208 6196 8260 6248
rect 10692 6196 10744 6248
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 18972 6332 19024 6384
rect 17040 6264 17092 6273
rect 12808 6196 12860 6248
rect 14004 6239 14056 6248
rect 14004 6205 14038 6239
rect 14038 6205 14056 6239
rect 8392 6171 8444 6180
rect 8392 6137 8426 6171
rect 8426 6137 8444 6171
rect 8392 6128 8444 6137
rect 1584 6060 1636 6112
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 6184 6103 6236 6112
rect 4896 6060 4948 6069
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 7564 6060 7616 6112
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 10876 6060 10928 6112
rect 11152 6128 11204 6180
rect 14004 6196 14056 6205
rect 16580 6196 16632 6248
rect 17684 6196 17736 6248
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 20812 6400 20864 6452
rect 22284 6400 22336 6452
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 22928 6264 22980 6316
rect 23388 6264 23440 6316
rect 14096 6128 14148 6180
rect 15844 6171 15896 6180
rect 15844 6137 15853 6171
rect 15853 6137 15887 6171
rect 15887 6137 15896 6171
rect 15844 6128 15896 6137
rect 16304 6171 16356 6180
rect 16304 6137 16313 6171
rect 16313 6137 16347 6171
rect 16347 6137 16356 6171
rect 16304 6128 16356 6137
rect 17500 6128 17552 6180
rect 17776 6128 17828 6180
rect 19340 6196 19392 6248
rect 22284 6196 22336 6248
rect 23572 6196 23624 6248
rect 24768 6196 24820 6248
rect 25136 6196 25188 6248
rect 19524 6171 19576 6180
rect 19524 6137 19558 6171
rect 19558 6137 19576 6171
rect 19524 6128 19576 6137
rect 19616 6128 19668 6180
rect 11336 6060 11388 6112
rect 13728 6060 13780 6112
rect 16488 6060 16540 6112
rect 19248 6060 19300 6112
rect 19984 6060 20036 6112
rect 20628 6103 20680 6112
rect 20628 6069 20637 6103
rect 20637 6069 20671 6103
rect 20671 6069 20680 6103
rect 20628 6060 20680 6069
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 22008 6103 22060 6112
rect 22008 6069 22017 6103
rect 22017 6069 22051 6103
rect 22051 6069 22060 6103
rect 22008 6060 22060 6069
rect 22560 6060 22612 6112
rect 25504 6103 25556 6112
rect 25504 6069 25513 6103
rect 25513 6069 25547 6103
rect 25547 6069 25556 6103
rect 25504 6060 25556 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 2688 5856 2740 5908
rect 3516 5856 3568 5908
rect 4436 5856 4488 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 6920 5856 6972 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 8852 5856 8904 5908
rect 9864 5856 9916 5908
rect 11060 5856 11112 5908
rect 11244 5899 11296 5908
rect 11244 5865 11253 5899
rect 11253 5865 11287 5899
rect 11287 5865 11296 5899
rect 11244 5856 11296 5865
rect 12440 5856 12492 5908
rect 13544 5856 13596 5908
rect 14004 5856 14056 5908
rect 14832 5856 14884 5908
rect 16120 5899 16172 5908
rect 10140 5788 10192 5840
rect 13176 5788 13228 5840
rect 2596 5720 2648 5772
rect 4068 5720 4120 5772
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 8484 5720 8536 5772
rect 9864 5720 9916 5772
rect 9956 5720 10008 5772
rect 11152 5720 11204 5772
rect 12808 5720 12860 5772
rect 16120 5865 16129 5899
rect 16129 5865 16163 5899
rect 16163 5865 16172 5899
rect 16120 5856 16172 5865
rect 16580 5856 16632 5908
rect 18880 5856 18932 5908
rect 20076 5856 20128 5908
rect 20444 5856 20496 5908
rect 20628 5856 20680 5908
rect 24676 5856 24728 5908
rect 24952 5856 25004 5908
rect 17040 5831 17092 5840
rect 17040 5797 17074 5831
rect 17074 5797 17092 5831
rect 17040 5788 17092 5797
rect 22560 5788 22612 5840
rect 23480 5788 23532 5840
rect 15844 5720 15896 5772
rect 16764 5763 16816 5772
rect 16764 5729 16773 5763
rect 16773 5729 16807 5763
rect 16807 5729 16816 5763
rect 16764 5720 16816 5729
rect 19616 5763 19668 5772
rect 19616 5729 19625 5763
rect 19625 5729 19659 5763
rect 19659 5729 19668 5763
rect 19616 5720 19668 5729
rect 21732 5720 21784 5772
rect 22284 5720 22336 5772
rect 22744 5720 22796 5772
rect 2688 5584 2740 5636
rect 3976 5584 4028 5636
rect 5264 5652 5316 5704
rect 10140 5695 10192 5704
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 2320 5559 2372 5568
rect 2320 5525 2329 5559
rect 2329 5525 2363 5559
rect 2363 5525 2372 5559
rect 2320 5516 2372 5525
rect 4252 5516 4304 5568
rect 4712 5516 4764 5568
rect 8392 5584 8444 5636
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 25136 5695 25188 5704
rect 9036 5584 9088 5636
rect 19524 5584 19576 5636
rect 25136 5661 25145 5695
rect 25145 5661 25179 5695
rect 25179 5661 25188 5695
rect 25136 5652 25188 5661
rect 23848 5584 23900 5636
rect 24860 5584 24912 5636
rect 25504 5652 25556 5704
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 11520 5516 11572 5525
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 19340 5516 19392 5568
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 21272 5559 21324 5568
rect 21272 5525 21281 5559
rect 21281 5525 21315 5559
rect 21315 5525 21324 5559
rect 21272 5516 21324 5525
rect 23388 5516 23440 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1676 5312 1728 5364
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2688 5176 2740 5228
rect 4068 5312 4120 5364
rect 4436 5312 4488 5364
rect 8576 5312 8628 5364
rect 8852 5312 8904 5364
rect 11336 5355 11388 5364
rect 11336 5321 11345 5355
rect 11345 5321 11379 5355
rect 11379 5321 11388 5355
rect 11336 5312 11388 5321
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 12348 5312 12400 5364
rect 12808 5312 12860 5364
rect 13544 5355 13596 5364
rect 13544 5321 13553 5355
rect 13553 5321 13587 5355
rect 13587 5321 13596 5355
rect 13544 5312 13596 5321
rect 14096 5312 14148 5364
rect 8484 5244 8536 5296
rect 5264 5176 5316 5228
rect 6644 5176 6696 5228
rect 13176 5244 13228 5296
rect 1584 5108 1636 5160
rect 4160 5108 4212 5160
rect 6460 5108 6512 5160
rect 6920 5108 6972 5160
rect 8944 5108 8996 5160
rect 14648 5176 14700 5228
rect 16764 5312 16816 5364
rect 17776 5355 17828 5364
rect 17776 5321 17785 5355
rect 17785 5321 17819 5355
rect 17819 5321 17828 5355
rect 20076 5355 20128 5364
rect 17776 5312 17828 5321
rect 16488 5287 16540 5296
rect 16488 5253 16497 5287
rect 16497 5253 16531 5287
rect 16531 5253 16540 5287
rect 16488 5244 16540 5253
rect 20076 5321 20085 5355
rect 20085 5321 20119 5355
rect 20119 5321 20128 5355
rect 20076 5312 20128 5321
rect 21732 5312 21784 5364
rect 25136 5312 25188 5364
rect 19524 5244 19576 5296
rect 24952 5244 25004 5296
rect 20628 5176 20680 5228
rect 24768 5176 24820 5228
rect 10784 5108 10836 5160
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 13820 5108 13872 5160
rect 4712 5040 4764 5092
rect 1492 4972 1544 5024
rect 2044 4972 2096 5024
rect 2596 4972 2648 5024
rect 5448 4972 5500 5024
rect 6920 4972 6972 5024
rect 9404 5040 9456 5092
rect 12532 5040 12584 5092
rect 12900 5040 12952 5092
rect 13636 5040 13688 5092
rect 14740 5108 14792 5160
rect 18144 5108 18196 5160
rect 15844 5040 15896 5092
rect 17500 5083 17552 5092
rect 17500 5049 17509 5083
rect 17509 5049 17543 5083
rect 17543 5049 17552 5083
rect 17500 5040 17552 5049
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 20260 4972 20312 5024
rect 21824 5108 21876 5160
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 20812 5040 20864 5092
rect 22744 5040 22796 5092
rect 24860 5040 24912 5092
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 22284 5015 22336 5024
rect 22284 4981 22293 5015
rect 22293 4981 22327 5015
rect 22327 4981 22336 5015
rect 22284 4972 22336 4981
rect 23204 4972 23256 5024
rect 24676 4972 24728 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1492 4768 1544 4820
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 2320 4768 2372 4820
rect 5172 4811 5224 4820
rect 5172 4777 5181 4811
rect 5181 4777 5215 4811
rect 5215 4777 5224 4811
rect 5172 4768 5224 4777
rect 5356 4768 5408 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 6736 4768 6788 4820
rect 8300 4768 8352 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 4252 4632 4304 4684
rect 6644 4632 6696 4684
rect 8208 4632 8260 4684
rect 9128 4632 9180 4684
rect 11244 4700 11296 4752
rect 11612 4700 11664 4752
rect 12164 4700 12216 4752
rect 12716 4768 12768 4820
rect 14004 4768 14056 4820
rect 14556 4768 14608 4820
rect 17132 4768 17184 4820
rect 17224 4811 17276 4820
rect 17224 4777 17233 4811
rect 17233 4777 17267 4811
rect 17267 4777 17276 4811
rect 17224 4768 17276 4777
rect 17868 4768 17920 4820
rect 19064 4811 19116 4820
rect 19064 4777 19073 4811
rect 19073 4777 19107 4811
rect 19107 4777 19116 4811
rect 19064 4768 19116 4777
rect 19156 4768 19208 4820
rect 19340 4768 19392 4820
rect 12624 4700 12676 4752
rect 13820 4700 13872 4752
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 13912 4632 13964 4684
rect 16580 4700 16632 4752
rect 17408 4700 17460 4752
rect 19524 4700 19576 4752
rect 20536 4768 20588 4820
rect 22008 4811 22060 4820
rect 22008 4777 22017 4811
rect 22017 4777 22051 4811
rect 22051 4777 22060 4811
rect 22008 4768 22060 4777
rect 22468 4811 22520 4820
rect 22468 4777 22477 4811
rect 22477 4777 22511 4811
rect 22511 4777 22520 4811
rect 22468 4768 22520 4777
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 21640 4700 21692 4752
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 8484 4607 8536 4616
rect 6920 4564 6972 4573
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 13084 4564 13136 4616
rect 4712 4539 4764 4548
rect 4712 4505 4721 4539
rect 4721 4505 4755 4539
rect 4755 4505 4764 4539
rect 4712 4496 4764 4505
rect 6460 4496 6512 4548
rect 7564 4496 7616 4548
rect 8944 4496 8996 4548
rect 10968 4496 11020 4548
rect 13636 4539 13688 4548
rect 13636 4505 13645 4539
rect 13645 4505 13679 4539
rect 13679 4505 13688 4539
rect 13636 4496 13688 4505
rect 13820 4496 13872 4548
rect 14832 4632 14884 4684
rect 17040 4632 17092 4684
rect 19432 4632 19484 4684
rect 20812 4632 20864 4684
rect 23388 4632 23440 4684
rect 25044 4675 25096 4684
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 15936 4607 15988 4616
rect 15016 4539 15068 4548
rect 15016 4505 15025 4539
rect 15025 4505 15059 4539
rect 15059 4505 15068 4539
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 22100 4564 22152 4616
rect 22284 4564 22336 4616
rect 15016 4496 15068 4505
rect 18972 4496 19024 4548
rect 21548 4496 21600 4548
rect 2688 4428 2740 4480
rect 4160 4428 4212 4480
rect 5356 4428 5408 4480
rect 6000 4428 6052 4480
rect 6276 4471 6328 4480
rect 6276 4437 6285 4471
rect 6285 4437 6319 4471
rect 6319 4437 6328 4471
rect 6276 4428 6328 4437
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 10784 4428 10836 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 17960 4428 18012 4437
rect 18696 4471 18748 4480
rect 18696 4437 18705 4471
rect 18705 4437 18739 4471
rect 18739 4437 18748 4471
rect 18696 4428 18748 4437
rect 22836 4428 22888 4480
rect 23848 4428 23900 4480
rect 27068 4428 27120 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 296 4088 348 4140
rect 2044 4156 2096 4208
rect 5448 4156 5500 4208
rect 6920 4224 6972 4276
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 11612 4267 11664 4276
rect 11612 4233 11621 4267
rect 11621 4233 11655 4267
rect 11655 4233 11664 4267
rect 11612 4224 11664 4233
rect 6736 4156 6788 4208
rect 13176 4156 13228 4208
rect 13912 4224 13964 4276
rect 14188 4224 14240 4276
rect 16212 4267 16264 4276
rect 16212 4233 16221 4267
rect 16221 4233 16255 4267
rect 16255 4233 16264 4267
rect 16212 4224 16264 4233
rect 17500 4224 17552 4276
rect 17960 4224 18012 4276
rect 19800 4224 19852 4276
rect 21640 4224 21692 4276
rect 23388 4267 23440 4276
rect 23388 4233 23397 4267
rect 23397 4233 23431 4267
rect 23431 4233 23440 4267
rect 23388 4224 23440 4233
rect 25044 4224 25096 4276
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 7564 4088 7616 4140
rect 1584 3884 1636 3936
rect 2596 4020 2648 4072
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 6184 4020 6236 4072
rect 9956 4088 10008 4140
rect 12072 4088 12124 4140
rect 13452 4088 13504 4140
rect 16948 4156 17000 4208
rect 14740 4088 14792 4140
rect 16396 4088 16448 4140
rect 8300 4020 8352 4072
rect 10784 4020 10836 4072
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 15292 4020 15344 4072
rect 16212 4020 16264 4072
rect 16856 4020 16908 4072
rect 24584 4156 24636 4208
rect 18696 4088 18748 4140
rect 20628 4088 20680 4140
rect 25504 4088 25556 4140
rect 22652 4020 22704 4072
rect 7932 3995 7984 4004
rect 7932 3961 7966 3995
rect 7966 3961 7984 3995
rect 7932 3952 7984 3961
rect 2872 3884 2924 3936
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 5540 3884 5592 3936
rect 6552 3884 6604 3936
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10140 3927 10192 3936
rect 10140 3893 10149 3927
rect 10149 3893 10183 3927
rect 10183 3893 10192 3927
rect 10140 3884 10192 3893
rect 16672 3995 16724 4004
rect 16672 3961 16681 3995
rect 16681 3961 16715 3995
rect 16715 3961 16724 3995
rect 16672 3952 16724 3961
rect 22100 3952 22152 4004
rect 23848 3952 23900 4004
rect 24216 3952 24268 4004
rect 10692 3884 10744 3936
rect 11060 3884 11112 3936
rect 13084 3927 13136 3936
rect 13084 3893 13093 3927
rect 13093 3893 13127 3927
rect 13127 3893 13136 3927
rect 13084 3884 13136 3893
rect 13176 3884 13228 3936
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 14648 3884 14700 3893
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 18972 3884 19024 3936
rect 19432 3884 19484 3936
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 22652 3927 22704 3936
rect 21180 3884 21232 3893
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 22836 3884 22888 3936
rect 23572 3884 23624 3936
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 24124 3927 24176 3936
rect 24124 3893 24133 3927
rect 24133 3893 24167 3927
rect 24167 3893 24176 3927
rect 24124 3884 24176 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2044 3723 2096 3732
rect 2044 3689 2053 3723
rect 2053 3689 2087 3723
rect 2087 3689 2096 3723
rect 2044 3680 2096 3689
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 2596 3680 2648 3732
rect 2964 3680 3016 3732
rect 6184 3680 6236 3732
rect 7288 3680 7340 3732
rect 7840 3680 7892 3732
rect 4068 3612 4120 3664
rect 7564 3612 7616 3664
rect 7748 3612 7800 3664
rect 1952 3544 2004 3596
rect 6552 3544 6604 3596
rect 7104 3544 7156 3596
rect 8208 3544 8260 3596
rect 2872 3476 2924 3528
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 8484 3680 8536 3732
rect 9312 3680 9364 3732
rect 10048 3680 10100 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 8668 3612 8720 3664
rect 9588 3544 9640 3596
rect 11152 3680 11204 3732
rect 12256 3723 12308 3732
rect 12256 3689 12265 3723
rect 12265 3689 12299 3723
rect 12299 3689 12308 3723
rect 12256 3680 12308 3689
rect 12348 3680 12400 3732
rect 13176 3680 13228 3732
rect 13360 3723 13412 3732
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 13452 3680 13504 3732
rect 14924 3680 14976 3732
rect 15292 3723 15344 3732
rect 15292 3689 15301 3723
rect 15301 3689 15335 3723
rect 15335 3689 15344 3723
rect 15292 3680 15344 3689
rect 15568 3680 15620 3732
rect 16396 3723 16448 3732
rect 16396 3689 16405 3723
rect 16405 3689 16439 3723
rect 16439 3689 16448 3723
rect 16396 3680 16448 3689
rect 17224 3680 17276 3732
rect 17408 3723 17460 3732
rect 17408 3689 17417 3723
rect 17417 3689 17451 3723
rect 17451 3689 17460 3723
rect 17408 3680 17460 3689
rect 17960 3680 18012 3732
rect 18696 3680 18748 3732
rect 19340 3680 19392 3732
rect 20904 3723 20956 3732
rect 20904 3689 20913 3723
rect 20913 3689 20947 3723
rect 20947 3689 20956 3723
rect 20904 3680 20956 3689
rect 21088 3680 21140 3732
rect 21916 3723 21968 3732
rect 21916 3689 21925 3723
rect 21925 3689 21959 3723
rect 21959 3689 21968 3723
rect 21916 3680 21968 3689
rect 22192 3680 22244 3732
rect 14648 3612 14700 3664
rect 17316 3612 17368 3664
rect 19524 3655 19576 3664
rect 19524 3621 19533 3655
rect 19533 3621 19567 3655
rect 19567 3621 19576 3655
rect 19524 3612 19576 3621
rect 20812 3612 20864 3664
rect 21180 3612 21232 3664
rect 21364 3612 21416 3664
rect 11520 3544 11572 3596
rect 16856 3587 16908 3596
rect 16856 3553 16865 3587
rect 16865 3553 16899 3587
rect 16899 3553 16908 3587
rect 16856 3544 16908 3553
rect 22744 3680 22796 3732
rect 23848 3655 23900 3664
rect 23848 3621 23882 3655
rect 23882 3621 23900 3655
rect 23848 3612 23900 3621
rect 13820 3519 13872 3528
rect 6276 3408 6328 3460
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 15844 3519 15896 3528
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 4344 3340 4396 3392
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 13544 3408 13596 3460
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 18512 3476 18564 3528
rect 20720 3476 20772 3528
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 23572 3519 23624 3528
rect 21456 3476 21508 3485
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 15016 3408 15068 3460
rect 18144 3408 18196 3460
rect 22652 3451 22704 3460
rect 22652 3417 22661 3451
rect 22661 3417 22695 3451
rect 22695 3417 22704 3451
rect 22652 3408 22704 3417
rect 7472 3340 7524 3392
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 14556 3340 14608 3392
rect 17040 3383 17092 3392
rect 17040 3349 17049 3383
rect 17049 3349 17083 3383
rect 17083 3349 17092 3383
rect 17040 3340 17092 3349
rect 18788 3340 18840 3392
rect 19892 3383 19944 3392
rect 19892 3349 19901 3383
rect 19901 3349 19935 3383
rect 19935 3349 19944 3383
rect 19892 3340 19944 3349
rect 24768 3340 24820 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3424 3136 3476 3188
rect 6092 3136 6144 3188
rect 7196 3136 7248 3188
rect 8300 3136 8352 3188
rect 6276 3043 6328 3052
rect 6276 3009 6285 3043
rect 6285 3009 6319 3043
rect 6319 3009 6328 3043
rect 7288 3043 7340 3052
rect 6276 3000 6328 3009
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 11152 3136 11204 3188
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 13544 3179 13596 3188
rect 12440 3136 12492 3145
rect 13544 3145 13553 3179
rect 13553 3145 13587 3179
rect 13587 3145 13596 3179
rect 13544 3136 13596 3145
rect 14096 3136 14148 3188
rect 15844 3136 15896 3188
rect 17316 3136 17368 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18696 3136 18748 3188
rect 20996 3136 21048 3188
rect 21548 3136 21600 3188
rect 22560 3136 22612 3188
rect 23848 3136 23900 3188
rect 25504 3179 25556 3188
rect 25504 3145 25513 3179
rect 25513 3145 25547 3179
rect 25547 3145 25556 3179
rect 25504 3136 25556 3145
rect 11796 3068 11848 3120
rect 11980 3068 12032 3120
rect 12348 3068 12400 3120
rect 11336 3043 11388 3052
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 3884 2932 3936 2984
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 4344 2932 4396 2984
rect 5632 2932 5684 2984
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 1676 2864 1728 2916
rect 2688 2864 2740 2916
rect 11336 3009 11345 3043
rect 11345 3009 11379 3043
rect 11379 3009 11388 3043
rect 11336 3000 11388 3009
rect 12900 3043 12952 3052
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 26056 3111 26108 3120
rect 26056 3077 26065 3111
rect 26065 3077 26099 3111
rect 26099 3077 26108 3111
rect 26056 3068 26108 3077
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 8668 2932 8720 2984
rect 9680 2932 9732 2984
rect 10140 2932 10192 2984
rect 12164 2975 12216 2984
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 12532 2932 12584 2984
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 14832 2932 14884 2984
rect 15016 2975 15068 2984
rect 15016 2941 15039 2975
rect 15039 2941 15068 2975
rect 15016 2932 15068 2941
rect 15568 2932 15620 2984
rect 18144 2932 18196 2984
rect 20904 2975 20956 2984
rect 20904 2941 20938 2975
rect 20938 2941 20956 2975
rect 7472 2864 7524 2916
rect 7564 2864 7616 2916
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 9864 2796 9916 2848
rect 10692 2796 10744 2848
rect 11612 2796 11664 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 17224 2796 17276 2848
rect 20904 2932 20956 2941
rect 22100 2932 22152 2984
rect 23572 2932 23624 2984
rect 24768 2932 24820 2984
rect 23756 2864 23808 2916
rect 20812 2796 20864 2848
rect 22008 2839 22060 2848
rect 22008 2805 22017 2839
rect 22017 2805 22051 2839
rect 22051 2805 22060 2839
rect 22008 2796 22060 2805
rect 22560 2839 22612 2848
rect 22560 2805 22569 2839
rect 22569 2805 22603 2839
rect 22603 2805 22612 2839
rect 22560 2796 22612 2805
rect 24124 2796 24176 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 1952 2592 2004 2644
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3884 2635 3936 2644
rect 3884 2601 3893 2635
rect 3893 2601 3927 2635
rect 3927 2601 3936 2635
rect 3884 2592 3936 2601
rect 5632 2592 5684 2644
rect 6368 2592 6420 2644
rect 1768 2524 1820 2576
rect 4252 2524 4304 2576
rect 4620 2499 4672 2508
rect 2964 2388 3016 2440
rect 4620 2465 4654 2499
rect 4654 2465 4672 2499
rect 4620 2456 4672 2465
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 7564 2456 7616 2508
rect 9680 2592 9732 2644
rect 11612 2592 11664 2644
rect 11520 2524 11572 2576
rect 14740 2592 14792 2644
rect 16856 2635 16908 2644
rect 12716 2524 12768 2576
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 8116 2388 8168 2440
rect 10048 2456 10100 2508
rect 10232 2431 10284 2440
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 10692 2456 10744 2508
rect 11796 2456 11848 2508
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 11152 2388 11204 2440
rect 18512 2592 18564 2644
rect 20812 2592 20864 2644
rect 18696 2524 18748 2576
rect 20720 2524 20772 2576
rect 21916 2592 21968 2644
rect 22560 2635 22612 2644
rect 22560 2601 22569 2635
rect 22569 2601 22603 2635
rect 22603 2601 22612 2635
rect 22560 2592 22612 2601
rect 24216 2635 24268 2644
rect 24216 2601 24225 2635
rect 24225 2601 24259 2635
rect 24259 2601 24268 2635
rect 24216 2592 24268 2601
rect 21456 2567 21508 2576
rect 21456 2533 21490 2567
rect 21490 2533 21508 2567
rect 21456 2524 21508 2533
rect 23756 2456 23808 2508
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 24768 2431 24820 2440
rect 24768 2397 24777 2431
rect 24777 2397 24811 2431
rect 24811 2397 24820 2431
rect 24768 2388 24820 2397
rect 9128 2363 9180 2372
rect 9128 2329 9137 2363
rect 9137 2329 9171 2363
rect 9171 2329 9180 2363
rect 9128 2320 9180 2329
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 23756 2295 23808 2304
rect 23756 2261 23765 2295
rect 23765 2261 23799 2295
rect 23799 2261 23808 2295
rect 23756 2252 23808 2261
rect 24032 2252 24084 2304
rect 24768 2252 24820 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 19432 620 19484 672
rect 4344 552 4396 604
rect 5264 552 5316 604
rect 8208 552 8260 604
rect 9588 552 9640 604
rect 20168 552 20220 604
rect 20628 552 20680 604
rect 21272 552 21324 604
<< metal2 >>
rect 1858 27568 1914 27577
rect 4618 27520 4674 28000
rect 13910 27520 13966 28000
rect 23202 27520 23258 28000
rect 24766 27568 24822 27577
rect 1858 27503 1914 27512
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1596 23322 1624 24783
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1412 22438 1440 23122
rect 1400 22432 1452 22438
rect 1400 22374 1452 22380
rect 1582 22128 1638 22137
rect 1582 22063 1638 22072
rect 1490 21448 1546 21457
rect 1490 21383 1546 21392
rect 1398 20768 1454 20777
rect 1398 20703 1454 20712
rect 1412 19174 1440 20703
rect 1504 20058 1532 21383
rect 1596 20602 1624 22063
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1582 20088 1638 20097
rect 1492 20052 1544 20058
rect 1582 20023 1638 20032
rect 1492 19994 1544 20000
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1490 18728 1546 18737
rect 1490 18663 1546 18672
rect 1398 17368 1454 17377
rect 1504 17338 1532 18663
rect 1596 18426 1624 20023
rect 1766 19408 1822 19417
rect 1872 19378 1900 27503
rect 4632 27418 4660 27520
rect 13924 27418 13952 27520
rect 4172 27390 4660 27418
rect 13832 27390 13952 27418
rect 2962 26888 3018 26897
rect 2962 26823 3018 26832
rect 2226 26208 2282 26217
rect 2226 26143 2282 26152
rect 1950 25528 2006 25537
rect 1950 25463 2006 25472
rect 1766 19343 1822 19352
rect 1860 19372 1912 19378
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1688 18766 1716 19246
rect 1676 18760 1728 18766
rect 1674 18728 1676 18737
rect 1728 18728 1730 18737
rect 1674 18663 1730 18672
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1582 18048 1638 18057
rect 1582 17983 1638 17992
rect 1398 17303 1454 17312
rect 1492 17332 1544 17338
rect 1412 15706 1440 17303
rect 1492 17274 1544 17280
rect 1596 16794 1624 17983
rect 1780 17882 1808 19343
rect 1860 19314 1912 19320
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1504 15978 1532 16594
rect 1582 16008 1638 16017
rect 1492 15972 1544 15978
rect 1582 15943 1638 15952
rect 1492 15914 1544 15920
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 1412 11218 1440 13194
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 8090 1440 11154
rect 1504 10985 1532 15914
rect 1596 14618 1624 15943
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 1688 14822 1716 15506
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 1596 12986 1624 13903
rect 1688 13841 1716 14758
rect 1674 13832 1730 13841
rect 1674 13767 1730 13776
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1872 12889 1900 15846
rect 1964 14074 1992 25463
rect 2134 23488 2190 23497
rect 2134 23423 2190 23432
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 2056 20058 2084 20198
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 2044 18080 2096 18086
rect 2042 18048 2044 18057
rect 2096 18048 2098 18057
rect 2042 17983 2098 17992
rect 2044 16992 2096 16998
rect 2042 16960 2044 16969
rect 2096 16960 2098 16969
rect 2042 16895 2098 16904
rect 2042 16688 2098 16697
rect 2042 16623 2098 16632
rect 2056 15162 2084 16623
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2056 13705 2084 13806
rect 2042 13696 2098 13705
rect 2042 13631 2098 13640
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1964 12986 1992 13330
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1858 12880 1914 12889
rect 1858 12815 1914 12824
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1872 12102 1900 12718
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1412 6866 1440 7686
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 296 4140 348 4146
rect 296 4082 348 4088
rect 308 480 336 4082
rect 1412 3505 1440 6802
rect 1504 6089 1532 10911
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1596 9722 1624 10066
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1688 7585 1716 10406
rect 1872 10266 1900 12038
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1964 9897 1992 12922
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1950 9888 2006 9897
rect 1950 9823 2006 9832
rect 2056 9466 2084 11494
rect 2148 10810 2176 23423
rect 2240 14006 2268 26143
rect 2778 24168 2834 24177
rect 2778 24103 2834 24112
rect 2688 22432 2740 22438
rect 2688 22374 2740 22380
rect 2700 20602 2728 22374
rect 2688 20596 2740 20602
rect 2688 20538 2740 20544
rect 2792 20482 2820 24103
rect 2516 20454 2820 20482
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2424 19174 2452 19858
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2332 17338 2360 17682
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2332 16250 2360 17274
rect 2424 17105 2452 19110
rect 2410 17096 2466 17105
rect 2410 17031 2466 17040
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2410 14512 2466 14521
rect 2410 14447 2412 14456
rect 2464 14447 2466 14456
rect 2412 14418 2464 14424
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2240 11354 2268 13330
rect 2332 12442 2360 14350
rect 2424 14074 2452 14418
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2516 13530 2544 20454
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2608 19174 2636 19858
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2608 17785 2636 19110
rect 2594 17776 2650 17785
rect 2594 17711 2650 17720
rect 2976 16114 3004 26823
rect 3882 22808 3938 22817
rect 3882 22743 3938 22752
rect 3056 20256 3108 20262
rect 3056 20198 3108 20204
rect 3068 19961 3096 20198
rect 3054 19952 3110 19961
rect 3054 19887 3110 19896
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2700 15978 2820 15994
rect 2688 15972 2832 15978
rect 2740 15966 2780 15972
rect 2688 15914 2740 15920
rect 2780 15914 2832 15920
rect 2688 15496 2740 15502
rect 2740 15456 2820 15484
rect 2688 15438 2740 15444
rect 2688 15360 2740 15366
rect 2594 15328 2650 15337
rect 2688 15302 2740 15308
rect 2594 15263 2650 15272
rect 2608 14618 2636 15263
rect 2700 15162 2728 15302
rect 2792 15162 2820 15456
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2686 14648 2742 14657
rect 2596 14612 2648 14618
rect 2686 14583 2742 14592
rect 2596 14554 2648 14560
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2608 12442 2636 14282
rect 2700 13530 2728 14583
rect 3054 13560 3110 13569
rect 2688 13524 2740 13530
rect 3054 13495 3110 13504
rect 2688 13466 2740 13472
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2700 12322 2728 13262
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2872 12368 2924 12374
rect 2700 12306 2820 12322
rect 2872 12310 2924 12316
rect 2688 12300 2820 12306
rect 2740 12294 2820 12300
rect 2688 12242 2740 12248
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11801 2360 12038
rect 2318 11792 2374 11801
rect 2318 11727 2320 11736
rect 2372 11727 2374 11736
rect 2320 11698 2372 11704
rect 2332 11667 2360 11698
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2332 11150 2360 11494
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1872 9438 2084 9466
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1582 6760 1638 6769
rect 1582 6695 1584 6704
rect 1636 6695 1638 6704
rect 1584 6666 1636 6672
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1584 6112 1636 6118
rect 1490 6080 1546 6089
rect 1584 6054 1636 6060
rect 1490 6015 1546 6024
rect 1596 5914 1624 6054
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1596 5166 1624 5850
rect 1688 5370 1716 6598
rect 1676 5364 1728 5370
rect 1728 5324 1808 5352
rect 1676 5306 1728 5312
rect 1584 5160 1636 5166
rect 1490 5128 1546 5137
rect 1584 5102 1636 5108
rect 1490 5063 1546 5072
rect 1504 5030 1532 5063
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4826 1532 4966
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1596 2990 1624 3878
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 846 2816 902 2825
rect 846 2751 902 2760
rect 860 480 888 2751
rect 1596 2650 1624 2926
rect 1688 2922 1716 3334
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1780 2582 1808 5324
rect 1872 3233 1900 9438
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1964 7313 1992 8910
rect 2056 8401 2084 9318
rect 2136 8424 2188 8430
rect 2042 8392 2098 8401
rect 2136 8366 2188 8372
rect 2042 8327 2098 8336
rect 2148 7546 2176 8366
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1950 7304 2006 7313
rect 1950 7239 2006 7248
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2148 6458 2176 6802
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5234 2084 5510
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2134 4992 2190 5001
rect 1950 4856 2006 4865
rect 1950 4791 1952 4800
rect 2004 4791 2006 4800
rect 1952 4762 2004 4768
rect 2056 4214 2084 4966
rect 2134 4927 2190 4936
rect 2044 4208 2096 4214
rect 2044 4150 2096 4156
rect 2042 3904 2098 3913
rect 2042 3839 2098 3848
rect 2056 3738 2084 3839
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1858 3224 1914 3233
rect 1858 3159 1914 3168
rect 1964 2650 1992 3538
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 1768 2576 1820 2582
rect 2148 2530 2176 4927
rect 1768 2518 1820 2524
rect 2056 2502 2176 2530
rect 1398 1728 1454 1737
rect 1398 1663 1454 1672
rect 1412 480 1440 1663
rect 2056 480 2084 2502
rect 2240 1057 2268 11018
rect 2332 10266 2360 11086
rect 2608 11082 2636 11494
rect 2792 11354 2820 12294
rect 2884 11898 2912 12310
rect 2976 12238 3004 12582
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2424 10146 2452 10950
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2332 10118 2452 10146
rect 2504 10192 2556 10198
rect 2608 10169 2636 10202
rect 2504 10134 2556 10140
rect 2594 10160 2650 10169
rect 2332 9926 2360 10118
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2332 9722 2360 9862
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2516 9178 2544 10134
rect 2594 10095 2650 10104
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2608 8838 2636 9998
rect 2700 9160 2728 11290
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2778 10296 2834 10305
rect 2778 10231 2780 10240
rect 2832 10231 2834 10240
rect 2780 10202 2832 10208
rect 2884 10146 2912 11222
rect 2792 10118 2912 10146
rect 2792 9654 2820 10118
rect 2872 10056 2924 10062
rect 2870 10024 2872 10033
rect 2964 10056 3016 10062
rect 2924 10024 2926 10033
rect 2964 9998 3016 10004
rect 2870 9959 2926 9968
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2780 9172 2832 9178
rect 2700 9132 2780 9160
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2332 8362 2360 8774
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2332 7970 2360 8298
rect 2332 7942 2452 7970
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 7002 2360 7754
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6798 2452 7942
rect 2516 7818 2544 8570
rect 2700 8022 2728 9132
rect 2780 9114 2832 9120
rect 2976 9110 3004 9998
rect 3068 9217 3096 13495
rect 3160 12986 3188 14758
rect 3238 13968 3294 13977
rect 3238 13903 3240 13912
rect 3292 13903 3294 13912
rect 3240 13874 3292 13880
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3344 12374 3372 19314
rect 3606 14376 3662 14385
rect 3606 14311 3662 14320
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 12714 3464 14214
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12850 3556 13126
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3332 12368 3384 12374
rect 3330 12336 3332 12345
rect 3384 12336 3386 12345
rect 3330 12271 3386 12280
rect 3424 12300 3476 12306
rect 3344 12245 3372 12271
rect 3424 12242 3476 12248
rect 3436 12209 3464 12242
rect 3422 12200 3478 12209
rect 3332 12164 3384 12170
rect 3422 12135 3478 12144
rect 3332 12106 3384 12112
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 3054 9208 3110 9217
rect 3054 9143 3110 9152
rect 2964 9104 3016 9110
rect 2870 9072 2926 9081
rect 2964 9046 3016 9052
rect 2870 9007 2872 9016
rect 2924 9007 2926 9016
rect 2872 8978 2924 8984
rect 2884 8090 2912 8978
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8294 3096 8910
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3068 8022 3096 8230
rect 2688 8016 2740 8022
rect 2594 7984 2650 7993
rect 2688 7958 2740 7964
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2594 7919 2596 7928
rect 2648 7919 2650 7928
rect 2596 7890 2648 7896
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2608 7002 2636 7890
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2700 7041 2728 7822
rect 2686 7032 2742 7041
rect 2596 6996 2648 7002
rect 2686 6967 2742 6976
rect 2596 6938 2648 6944
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2700 6746 2728 6967
rect 2870 6896 2926 6905
rect 2870 6831 2926 6840
rect 2884 6798 2912 6831
rect 2872 6792 2924 6798
rect 2700 6718 2820 6746
rect 2872 6734 2924 6740
rect 2792 6458 2820 6718
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2884 6390 2912 6734
rect 3160 6458 3188 11018
rect 3252 10849 3280 12038
rect 3238 10840 3294 10849
rect 3238 10775 3294 10784
rect 3252 9518 3280 10775
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3240 9376 3292 9382
rect 3344 9330 3372 12106
rect 3436 11898 3464 12135
rect 3514 11928 3570 11937
rect 3424 11892 3476 11898
rect 3514 11863 3570 11872
rect 3424 11834 3476 11840
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 9994 3464 10474
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3436 9586 3464 9930
rect 3528 9761 3556 11863
rect 3620 11218 3648 14311
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3804 13190 3832 13738
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12850 3832 13126
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3896 10130 3924 22743
rect 4172 14346 4200 27390
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 13832 23338 13860 27390
rect 14096 26308 14148 26314
rect 14096 26250 14148 26256
rect 13740 23310 13860 23338
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 13266 22672 13322 22681
rect 13266 22607 13322 22616
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 12346 19952 12402 19961
rect 12346 19887 12402 19896
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 12360 18970 12388 19887
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12440 18760 12492 18766
rect 11518 18728 11574 18737
rect 12440 18702 12492 18708
rect 11518 18663 11574 18672
rect 12256 18692 12308 18698
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 7194 18048 7250 18057
rect 7194 17983 7250 17992
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 4802 16960 4858 16969
rect 4802 16895 4858 16904
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 14958 4292 15302
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4264 14618 4292 14894
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4172 14006 4200 14282
rect 4448 14074 4476 14418
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 4172 13394 4200 13942
rect 4160 13388 4212 13394
rect 4212 13348 4292 13376
rect 4160 13330 4212 13336
rect 4264 12986 4292 13348
rect 4252 12980 4304 12986
rect 4304 12940 4384 12968
rect 4252 12922 4304 12928
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4264 12170 4292 12650
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4356 11694 4384 12940
rect 4448 12442 4476 14010
rect 4528 13864 4580 13870
rect 4632 13852 4660 14350
rect 4580 13824 4660 13852
rect 4710 13832 4766 13841
rect 4528 13806 4580 13812
rect 4710 13767 4766 13776
rect 4618 13696 4674 13705
rect 4618 13631 4674 13640
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4540 12850 4568 13330
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4632 12782 4660 13631
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4344 11688 4396 11694
rect 4396 11648 4476 11676
rect 4344 11630 4396 11636
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3988 11082 4016 11562
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3514 9752 3570 9761
rect 3514 9687 3570 9696
rect 3620 9636 3648 9998
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3528 9608 3648 9636
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3528 9382 3556 9608
rect 3292 9324 3372 9330
rect 3240 9318 3372 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3252 9302 3372 9318
rect 3252 8566 3280 9302
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3606 8256 3662 8265
rect 3606 8191 3662 8200
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 6730 3280 7210
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 3160 6254 3188 6394
rect 3344 6322 3372 7754
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6798 3556 7142
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3528 6322 3556 6734
rect 3620 6497 3648 8191
rect 3896 7818 3924 9862
rect 4172 9654 4200 10066
rect 4356 9654 4384 11290
rect 4448 10606 4476 11648
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4632 10810 4660 11086
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 10062 4476 10542
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 9042 4200 9318
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3792 7744 3844 7750
rect 3698 7712 3754 7721
rect 3792 7686 3844 7692
rect 3698 7647 3754 7656
rect 3712 7449 3740 7647
rect 3698 7440 3754 7449
rect 3698 7375 3754 7384
rect 3606 6488 3662 6497
rect 3606 6423 3662 6432
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2686 6080 2742 6089
rect 2686 6015 2742 6024
rect 2700 5914 2728 6015
rect 3528 5914 3556 6258
rect 2688 5908 2740 5914
rect 3516 5908 3568 5914
rect 2740 5868 2820 5896
rect 2688 5850 2740 5856
rect 2700 5785 2728 5850
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 4826 2360 5510
rect 2608 5137 2636 5714
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2700 5234 2728 5578
rect 2792 5370 2820 5868
rect 3516 5850 3568 5856
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2594 5128 2650 5137
rect 2594 5063 2650 5072
rect 2608 5030 2636 5063
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2502 4856 2558 4865
rect 2320 4820 2372 4826
rect 2502 4791 2558 4800
rect 2320 4762 2372 4768
rect 2516 3738 2544 4791
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2608 4078 2636 4558
rect 2700 4486 2728 5170
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2608 3738 2636 4014
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2700 2922 2728 4422
rect 3804 4185 3832 7686
rect 3988 7478 4016 8842
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4080 8129 4108 8774
rect 4172 8344 4200 8978
rect 4356 8634 4384 8978
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4252 8356 4304 8362
rect 4172 8316 4252 8344
rect 4252 8298 4304 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3976 7472 4028 7478
rect 4172 7449 4200 7890
rect 3976 7414 4028 7420
rect 4158 7440 4214 7449
rect 4158 7375 4160 7384
rect 4212 7375 4214 7384
rect 4160 7346 4212 7352
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3988 5817 4016 6938
rect 4264 6610 4292 8298
rect 4724 8090 4752 13767
rect 4816 12714 4844 16895
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6366 15192 6422 15201
rect 6366 15127 6422 15136
rect 4986 15056 5042 15065
rect 4986 14991 5042 15000
rect 5724 15020 5776 15026
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4816 12102 4844 12650
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4816 11257 4844 12038
rect 4802 11248 4858 11257
rect 4802 11183 4858 11192
rect 4894 10840 4950 10849
rect 4894 10775 4896 10784
rect 4948 10775 4950 10784
rect 4896 10746 4948 10752
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4620 7880 4672 7886
rect 4434 7848 4490 7857
rect 4620 7822 4672 7828
rect 4434 7783 4490 7792
rect 4172 6582 4292 6610
rect 4172 6390 4200 6582
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3974 5808 4030 5817
rect 3974 5743 4030 5752
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3974 5672 4030 5681
rect 3974 5607 3976 5616
rect 4028 5607 4030 5616
rect 3976 5578 4028 5584
rect 4080 5370 4108 5714
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4172 5166 4200 6326
rect 4448 5914 4476 7783
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4172 4486 4200 5102
rect 4264 4690 4292 5510
rect 4448 5370 4476 5850
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3790 4176 3846 4185
rect 3790 4111 3846 4120
rect 3422 4040 3478 4049
rect 3422 3975 3478 3984
rect 3606 4040 3662 4049
rect 3606 3975 3662 3984
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2778 3768 2834 3777
rect 2778 3703 2834 3712
rect 2792 3097 2820 3703
rect 2884 3534 2912 3878
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2778 3088 2834 3097
rect 2778 3023 2834 3032
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 2318 2680 2374 2689
rect 2884 2650 2912 3470
rect 2976 3194 3004 3674
rect 3436 3194 3464 3975
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 2318 2615 2320 2624
rect 2372 2615 2374 2624
rect 2872 2644 2924 2650
rect 2320 2586 2372 2592
rect 2872 2586 2924 2592
rect 2976 2446 3004 3130
rect 3146 3088 3202 3097
rect 3146 3023 3202 3032
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2594 2000 2650 2009
rect 2594 1935 2650 1944
rect 2226 1048 2282 1057
rect 2226 983 2282 992
rect 2608 480 2636 1935
rect 3160 480 3188 3023
rect 3620 2417 3648 3975
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3670 4108 3878
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4068 3528 4120 3534
rect 4172 3482 4200 4422
rect 4120 3476 4200 3482
rect 4068 3470 4200 3476
rect 4080 3454 4200 3470
rect 3790 3224 3846 3233
rect 3790 3159 3846 3168
rect 3804 2961 3832 3159
rect 4080 2990 4108 3454
rect 3884 2984 3936 2990
rect 3790 2952 3846 2961
rect 3884 2926 3936 2932
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 3790 2887 3846 2896
rect 3606 2408 3662 2417
rect 3606 2343 3662 2352
rect 3804 480 3832 2887
rect 3896 2650 3924 2926
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 4264 2582 4292 4626
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4356 2990 4384 3334
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 4540 2417 4568 7482
rect 4632 6662 4660 7822
rect 4724 7546 4752 8026
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4894 7168 4950 7177
rect 4894 7103 4950 7112
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4908 6118 4936 7103
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5098 4752 5510
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4724 4554 4752 5034
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4618 2544 4674 2553
rect 4618 2479 4620 2488
rect 4672 2479 4674 2488
rect 4620 2450 4672 2456
rect 4526 2408 4582 2417
rect 4526 2343 4582 2352
rect 4066 1320 4122 1329
rect 4066 1255 4122 1264
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 2042 0 2098 480
rect 2594 0 2650 480
rect 3146 0 3202 480
rect 3790 0 3846 480
rect 4080 377 4108 1255
rect 4344 604 4396 610
rect 4344 546 4396 552
rect 4356 480 4384 546
rect 4908 480 4936 6054
rect 5000 1873 5028 14991
rect 5724 14962 5776 14968
rect 5736 14550 5764 14962
rect 5724 14544 5776 14550
rect 5552 14504 5724 14532
rect 5552 14074 5580 14504
rect 5724 14486 5776 14492
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 6012 14006 6040 14214
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5644 13530 5672 13738
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5080 12776 5132 12782
rect 5078 12744 5080 12753
rect 5132 12744 5134 12753
rect 5078 12679 5134 12688
rect 5184 12594 5212 12786
rect 5092 12566 5212 12594
rect 5092 12238 5120 12566
rect 6184 12368 6236 12374
rect 5998 12336 6054 12345
rect 6184 12310 6236 12316
rect 5998 12271 6054 12280
rect 6092 12300 6144 12306
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5092 11898 5120 12174
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 6012 11218 6040 12271
rect 6092 12242 6144 12248
rect 6104 11626 6132 12242
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5540 11076 5592 11082
rect 5460 11036 5540 11064
rect 5080 11008 5132 11014
rect 5078 10976 5080 10985
rect 5132 10976 5134 10985
rect 5078 10911 5134 10920
rect 5092 10674 5120 10911
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5354 10568 5410 10577
rect 5354 10503 5356 10512
rect 5408 10503 5410 10512
rect 5356 10474 5408 10480
rect 5172 9920 5224 9926
rect 5368 9897 5396 10474
rect 5172 9862 5224 9868
rect 5354 9888 5410 9897
rect 5184 9586 5212 9862
rect 5354 9823 5410 9832
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5460 9518 5488 11036
rect 5540 11018 5592 11024
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10674 6040 10950
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5998 9888 6054 9897
rect 5622 9820 5918 9840
rect 5998 9823 6054 9832
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9722 6040 9823
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8498 5488 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 8090 5304 8366
rect 5538 8120 5594 8129
rect 5264 8084 5316 8090
rect 5538 8055 5594 8064
rect 5814 8120 5870 8129
rect 5814 8055 5816 8064
rect 5264 8026 5316 8032
rect 5552 7342 5580 8055
rect 5868 8055 5870 8064
rect 5816 8026 5868 8032
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5540 7200 5592 7206
rect 5460 7148 5540 7154
rect 5460 7142 5592 7148
rect 5460 7126 5580 7142
rect 5460 6798 5488 7126
rect 5828 6934 5856 7346
rect 6012 7342 6040 9318
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6012 6934 6040 7278
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6322 5120 6598
rect 5460 6390 5488 6734
rect 5552 6458 5580 6802
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5630 6216 5686 6225
rect 5630 6151 5686 6160
rect 5644 5914 5672 6151
rect 5632 5908 5684 5914
rect 5368 5868 5632 5896
rect 5264 5704 5316 5710
rect 5170 5672 5226 5681
rect 5264 5646 5316 5652
rect 5170 5607 5226 5616
rect 5184 4826 5212 5607
rect 5276 5234 5304 5646
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4986 1864 5042 1873
rect 4986 1799 5042 1808
rect 5276 610 5304 5170
rect 5368 4826 5396 5868
rect 5632 5850 5684 5856
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5540 5568 5592 5574
rect 6012 5545 6040 5714
rect 5540 5510 5592 5516
rect 5998 5536 6054 5545
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5460 4622 5488 4966
rect 5552 4865 5580 5510
rect 5622 5468 5918 5488
rect 5998 5471 6054 5480
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5814 5128 5870 5137
rect 5814 5063 5870 5072
rect 5828 4865 5856 5063
rect 5538 4856 5594 4865
rect 5538 4791 5594 4800
rect 5814 4856 5870 4865
rect 5814 4791 5870 4800
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5356 4480 5408 4486
rect 5354 4448 5356 4457
rect 5408 4448 5410 4457
rect 5354 4383 5410 4392
rect 5460 4214 5488 4558
rect 6012 4486 6040 5471
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5552 4078 5580 4111
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5552 480 5580 3878
rect 6104 3584 6132 11562
rect 6196 11558 6224 12310
rect 6380 12306 6408 15127
rect 6748 14890 6776 15438
rect 6840 15026 6868 15506
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7116 15162 7144 15438
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6748 14793 6776 14826
rect 6734 14784 6790 14793
rect 6734 14719 6790 14728
rect 7024 14006 7052 14826
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7102 13968 7158 13977
rect 6826 12472 6882 12481
rect 6826 12407 6882 12416
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6184 11552 6236 11558
rect 6182 11520 6184 11529
rect 6236 11520 6238 11529
rect 6182 11455 6238 11464
rect 6288 11286 6316 12038
rect 6656 11354 6684 12038
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6196 10538 6224 11086
rect 6274 10840 6330 10849
rect 6274 10775 6330 10784
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6288 10198 6316 10775
rect 6472 10674 6500 11086
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6472 10130 6500 10610
rect 6564 10470 6592 11154
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6472 9926 6500 10066
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6196 7342 6224 7890
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6196 6322 6224 7278
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 4078 6224 6054
rect 6288 5681 6316 8774
rect 6380 7041 6408 9318
rect 6472 8498 6500 9862
rect 6564 9330 6592 10406
rect 6564 9302 6684 9330
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6564 8362 6592 8910
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6472 7478 6500 7890
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6366 7032 6422 7041
rect 6366 6967 6422 6976
rect 6274 5672 6330 5681
rect 6274 5607 6330 5616
rect 6460 5160 6512 5166
rect 6366 5128 6422 5137
rect 6460 5102 6512 5108
rect 6366 5063 6422 5072
rect 6380 4826 6408 5063
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6472 4554 6500 5102
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6196 3738 6224 4014
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6104 3556 6224 3584
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6104 3194 6132 3334
rect 6092 3188 6144 3194
rect 6012 3148 6092 3176
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2650 5672 2926
rect 6012 2689 6040 3148
rect 6092 3130 6144 3136
rect 6196 2836 6224 3556
rect 6288 3466 6316 4422
rect 6564 3942 6592 8298
rect 6656 7954 6684 9302
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6748 8498 6776 8774
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6642 6352 6698 6361
rect 6642 6287 6698 6296
rect 6656 5234 6684 6287
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6734 5128 6790 5137
rect 6734 5063 6790 5072
rect 6748 4826 6776 5063
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6642 4720 6698 4729
rect 6642 4655 6644 4664
rect 6696 4655 6698 4664
rect 6644 4626 6696 4632
rect 6748 4214 6776 4762
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6840 4060 6868 12407
rect 7024 11898 7052 13942
rect 7102 13903 7158 13912
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7024 11286 7052 11834
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7116 10810 7144 13903
rect 7208 10985 7236 17983
rect 9692 17898 9720 18294
rect 10980 18290 11008 18566
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9600 17882 9720 17898
rect 9588 17876 9720 17882
rect 9640 17870 9720 17876
rect 9588 17818 9640 17824
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7286 16688 7342 16697
rect 7286 16623 7342 16632
rect 7194 10976 7250 10985
rect 7194 10911 7250 10920
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7208 10742 7236 10911
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7194 10024 7250 10033
rect 7104 9988 7156 9994
rect 7194 9959 7250 9968
rect 7104 9930 7156 9936
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7342 6960 7754
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 6730 6960 7278
rect 7024 7002 7052 9318
rect 7116 9178 7144 9930
rect 7208 9178 7236 9959
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7116 7750 7144 8298
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7177 7144 7686
rect 7102 7168 7158 7177
rect 7102 7103 7158 7112
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6458 6960 6666
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6932 5914 6960 6394
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6932 5166 6960 5510
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4622 6960 4966
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6932 4282 6960 4558
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6748 4032 6868 4060
rect 6552 3936 6604 3942
rect 6366 3904 6422 3913
rect 6552 3878 6604 3884
rect 6366 3839 6422 3848
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6288 2961 6316 2994
rect 6274 2952 6330 2961
rect 6274 2887 6330 2896
rect 6196 2808 6316 2836
rect 5998 2680 6054 2689
rect 5632 2644 5684 2650
rect 6288 2666 6316 2808
rect 5998 2615 6054 2624
rect 6104 2638 6316 2666
rect 6380 2650 6408 3839
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6564 2854 6592 3538
rect 6552 2848 6604 2854
rect 6550 2816 6552 2825
rect 6604 2816 6606 2825
rect 6550 2751 6606 2760
rect 6748 2666 6776 4032
rect 7300 3738 7328 16623
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 11694 7420 14758
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13802 7512 14214
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7484 13462 7512 13738
rect 7576 13530 7604 15914
rect 8208 15156 8260 15162
rect 8312 15144 8340 17138
rect 9600 17134 9628 17818
rect 9678 17776 9734 17785
rect 9678 17711 9734 17720
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8260 15116 8340 15144
rect 8208 15098 8260 15104
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 8036 14618 8064 14826
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8036 14074 8064 14554
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 7484 12170 7512 13398
rect 8036 12986 8064 13398
rect 8128 13326 8156 13738
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7760 12442 7788 12922
rect 8128 12918 8156 13262
rect 8220 12986 8248 13330
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 8114 12608 8170 12617
rect 8114 12543 8170 12552
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7562 12336 7618 12345
rect 8128 12306 8156 12543
rect 7562 12271 7618 12280
rect 8116 12300 8168 12306
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 11354 7420 11630
rect 7484 11506 7512 12106
rect 7576 11801 7604 12271
rect 8116 12242 8168 12248
rect 7932 12232 7984 12238
rect 7838 12200 7894 12209
rect 7932 12174 7984 12180
rect 7838 12135 7894 12144
rect 7562 11792 7618 11801
rect 7562 11727 7618 11736
rect 7852 11694 7880 12135
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7484 11478 7604 11506
rect 7470 11384 7526 11393
rect 7380 11348 7432 11354
rect 7470 11319 7526 11328
rect 7380 11290 7432 11296
rect 7378 10296 7434 10305
rect 7378 10231 7380 10240
rect 7432 10231 7434 10240
rect 7380 10202 7432 10208
rect 7484 10146 7512 11319
rect 7576 11218 7604 11478
rect 7944 11354 7972 12174
rect 8312 11937 8340 15116
rect 8404 14618 8432 15642
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8496 14822 8524 15438
rect 8588 15201 8616 15846
rect 9232 15706 9260 16934
rect 9324 16794 9352 16934
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9324 16250 9352 16730
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9416 16153 9444 16390
rect 9402 16144 9458 16153
rect 9312 16108 9364 16114
rect 9402 16079 9458 16088
rect 9312 16050 9364 16056
rect 9324 16017 9352 16050
rect 9416 16046 9444 16079
rect 9404 16040 9456 16046
rect 9310 16008 9366 16017
rect 9404 15982 9456 15988
rect 9310 15943 9366 15952
rect 9692 15910 9720 17711
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9784 15722 9812 18022
rect 10060 17542 10088 18090
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 16130 10088 17478
rect 10336 17338 10364 17682
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10324 17332 10376 17338
rect 10152 17292 10324 17320
rect 10152 16250 10180 17292
rect 10324 17274 10376 17280
rect 10888 17134 10916 17478
rect 10876 17128 10928 17134
rect 10598 17096 10654 17105
rect 10598 17031 10600 17040
rect 10652 17031 10654 17040
rect 10796 17088 10876 17116
rect 10600 17002 10652 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10692 16720 10744 16726
rect 10796 16697 10824 17088
rect 10876 17070 10928 17076
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16726 10916 16934
rect 10876 16720 10928 16726
rect 10692 16662 10744 16668
rect 10782 16688 10838 16697
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10060 16102 10180 16130
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9692 15694 9812 15722
rect 9586 15600 9642 15609
rect 9586 15535 9642 15544
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8574 15192 8630 15201
rect 8574 15127 8630 15136
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8680 14618 8708 15370
rect 9600 15366 9628 15535
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9496 14952 9548 14958
rect 8850 14920 8906 14929
rect 9496 14894 9548 14900
rect 8850 14855 8906 14864
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8864 14521 8892 14855
rect 8850 14512 8906 14521
rect 8850 14447 8906 14456
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8588 13530 8616 14010
rect 8576 13524 8628 13530
rect 8628 13484 8708 13512
rect 8576 13466 8628 13472
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8404 12238 8432 12786
rect 8588 12782 8616 13262
rect 8680 12850 8708 13484
rect 8758 13016 8814 13025
rect 8758 12951 8814 12960
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8772 12714 8800 12951
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8298 11928 8354 11937
rect 8404 11898 8432 12174
rect 8298 11863 8354 11872
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7656 11280 7708 11286
rect 8024 11280 8076 11286
rect 7656 11222 7708 11228
rect 7838 11248 7894 11257
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7668 10674 7696 11222
rect 8024 11222 8076 11228
rect 7838 11183 7894 11192
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7562 10296 7618 10305
rect 7562 10231 7618 10240
rect 7392 10118 7512 10146
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7116 3097 7144 3538
rect 7194 3224 7250 3233
rect 7194 3159 7196 3168
rect 7248 3159 7250 3168
rect 7196 3130 7248 3136
rect 7102 3088 7158 3097
rect 7102 3023 7158 3032
rect 7208 2990 7236 3130
rect 7286 3088 7342 3097
rect 7286 3023 7288 3032
rect 7340 3023 7342 3032
rect 7288 2994 7340 3000
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7392 2802 7420 10118
rect 7470 9616 7526 9625
rect 7470 9551 7526 9560
rect 7484 8537 7512 9551
rect 7576 8634 7604 10231
rect 7668 9518 7696 10610
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7470 8528 7526 8537
rect 7470 8463 7526 8472
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 8090 7512 8230
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7484 6254 7512 8026
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 7585 7696 7686
rect 7654 7576 7710 7585
rect 7654 7511 7710 7520
rect 7760 7426 7788 7822
rect 7668 7398 7788 7426
rect 7668 6662 7696 7398
rect 7852 7290 7880 11183
rect 8036 10810 8064 11222
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8208 10600 8260 10606
rect 8312 10588 8340 11494
rect 8392 11280 8444 11286
rect 8390 11248 8392 11257
rect 8444 11248 8446 11257
rect 8390 11183 8446 11192
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8404 10985 8432 11086
rect 8390 10976 8446 10985
rect 8390 10911 8446 10920
rect 8260 10560 8340 10588
rect 8208 10542 8260 10548
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 10130 8156 10474
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 7944 9382 7972 10066
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 8673 7972 9318
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7930 8664 7986 8673
rect 7930 8599 7986 8608
rect 8036 8430 8064 9114
rect 8128 8820 8156 10066
rect 8220 10062 8248 10542
rect 8496 10266 8524 11086
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8312 9178 8340 10202
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8588 8974 8616 9386
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8838 8616 8910
rect 8300 8832 8352 8838
rect 8128 8800 8300 8820
rect 8576 8832 8628 8838
rect 8352 8800 8354 8809
rect 8128 8792 8298 8800
rect 8576 8774 8628 8780
rect 8298 8735 8354 8744
rect 8482 8528 8538 8537
rect 8482 8463 8538 8472
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8036 8276 8064 8366
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8116 8288 8168 8294
rect 8036 8248 8116 8276
rect 8312 8242 8340 8298
rect 8116 8230 8168 8236
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 8036 7478 8064 7890
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8036 7313 8064 7414
rect 7760 7262 7880 7290
rect 8022 7304 8078 7313
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7484 4146 7512 4927
rect 7576 4554 7604 6054
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7576 4146 7604 4490
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7668 3777 7696 6598
rect 7654 3768 7710 3777
rect 7654 3703 7710 3712
rect 7760 3670 7788 7262
rect 8022 7239 8078 7248
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8036 5914 8064 6802
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4185 7972 4422
rect 7930 4176 7986 4185
rect 7930 4111 7986 4120
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 7944 3777 7972 3946
rect 7930 3768 7986 3777
rect 7840 3732 7892 3738
rect 7930 3703 7986 3712
rect 7840 3674 7892 3680
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 2922 7512 3334
rect 7576 2922 7604 3606
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 6368 2644 6420 2650
rect 5632 2586 5684 2592
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 480 6132 2638
rect 6368 2586 6420 2592
rect 6656 2638 6776 2666
rect 7208 2774 7420 2802
rect 7208 2666 7236 2774
rect 7208 2638 7328 2666
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6380 2009 6408 2450
rect 6366 2000 6422 2009
rect 6366 1935 6422 1944
rect 6656 480 6684 2638
rect 7300 480 7328 2638
rect 7484 2446 7512 2858
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7392 1737 7420 2382
rect 7576 1873 7604 2450
rect 7562 1864 7618 1873
rect 7562 1799 7618 1808
rect 7378 1728 7434 1737
rect 7378 1663 7434 1672
rect 7852 480 7880 3674
rect 8128 3482 8156 8230
rect 8220 8214 8340 8242
rect 8220 6254 8248 8214
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8312 5001 8340 7142
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8404 5642 8432 6122
rect 8496 5778 8524 8463
rect 8588 8362 8616 8774
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8390 5536 8446 5545
rect 8390 5471 8446 5480
rect 8298 4992 8354 5001
rect 8298 4927 8354 4936
rect 8312 4826 8340 4927
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8220 3602 8248 4626
rect 8312 4185 8340 4762
rect 8298 4176 8354 4185
rect 8298 4111 8354 4120
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8128 3454 8248 3482
rect 8114 2816 8170 2825
rect 8114 2751 8170 2760
rect 8128 2446 8156 2751
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8220 610 8248 3454
rect 8312 3194 8340 4014
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8208 604 8260 610
rect 8208 546 8260 552
rect 8404 480 8432 5471
rect 8496 5302 8524 5714
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8496 3738 8524 4558
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8588 1465 8616 5306
rect 8680 3670 8708 7958
rect 8772 4434 8800 8026
rect 8864 5914 8892 14447
rect 9402 13968 9458 13977
rect 9402 13903 9458 13912
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9324 12481 9352 12718
rect 9310 12472 9366 12481
rect 9310 12407 9366 12416
rect 9310 10568 9366 10577
rect 9310 10503 9366 10512
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8942 10024 8998 10033
rect 8942 9959 8944 9968
rect 8996 9959 8998 9968
rect 8944 9930 8996 9936
rect 9048 9518 9076 10406
rect 9324 9654 9352 10503
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9036 9512 9088 9518
rect 9034 9480 9036 9489
rect 9088 9480 9090 9489
rect 9034 9415 9090 9424
rect 9324 9042 9352 9590
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9324 8430 9352 8978
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9312 7472 9364 7478
rect 9310 7440 9312 7449
rect 9364 7440 9366 7449
rect 9310 7375 9366 7384
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 6662 9352 7142
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 8956 6225 8984 6598
rect 8942 6216 8998 6225
rect 8942 6151 8998 6160
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8864 5370 8892 5850
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8956 4554 8984 5102
rect 9048 4826 9076 5578
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9140 4690 9168 6598
rect 9416 5658 9444 13903
rect 9508 11778 9536 14894
rect 9692 12322 9720 15694
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9784 14482 9812 15098
rect 9864 14816 9916 14822
rect 10046 14784 10102 14793
rect 9916 14764 9996 14770
rect 9864 14758 9996 14764
rect 9876 14742 9996 14758
rect 9968 14482 9996 14742
rect 10046 14719 10102 14728
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9784 14074 9812 14418
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9968 13870 9996 14418
rect 9956 13864 10008 13870
rect 9770 13832 9826 13841
rect 9956 13806 10008 13812
rect 9770 13767 9826 13776
rect 9600 12294 9720 12322
rect 9600 12073 9628 12294
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9586 12064 9642 12073
rect 9586 11999 9642 12008
rect 9692 11937 9720 12174
rect 9678 11928 9734 11937
rect 9678 11863 9680 11872
rect 9732 11863 9734 11872
rect 9680 11834 9732 11840
rect 9508 11762 9720 11778
rect 9508 11756 9732 11762
rect 9508 11750 9680 11756
rect 9680 11698 9732 11704
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9508 10266 9536 10678
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 10305 9720 10406
rect 9678 10296 9734 10305
rect 9496 10260 9548 10266
rect 9678 10231 9734 10240
rect 9496 10202 9548 10208
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9692 8072 9720 9658
rect 9600 8044 9720 8072
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9508 6458 9536 6734
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9324 5630 9444 5658
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8772 4406 8984 4434
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8680 2990 8708 3606
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8956 2428 8984 4406
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9048 2961 9076 3878
rect 9324 3738 9352 5630
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5098 9444 5510
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9600 4604 9628 8044
rect 9678 7984 9734 7993
rect 9678 7919 9734 7928
rect 9692 7546 9720 7919
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 6866 9720 7278
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 4729 9720 6598
rect 9678 4720 9734 4729
rect 9678 4655 9734 4664
rect 9600 4576 9720 4604
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9586 3632 9642 3641
rect 9586 3567 9588 3576
rect 9640 3567 9642 3576
rect 9588 3538 9640 3544
rect 9692 2990 9720 4576
rect 9680 2984 9732 2990
rect 9034 2952 9090 2961
rect 9680 2926 9732 2932
rect 9034 2887 9090 2896
rect 9048 2553 9076 2887
rect 9784 2802 9812 13767
rect 9954 13560 10010 13569
rect 9954 13495 10010 13504
rect 9968 13258 9996 13495
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9876 12170 9904 12786
rect 9956 12640 10008 12646
rect 9954 12608 9956 12617
rect 10008 12608 10010 12617
rect 9954 12543 10010 12552
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9862 11928 9918 11937
rect 9862 11863 9918 11872
rect 9876 11529 9904 11863
rect 10060 11665 10088 14719
rect 10152 11937 10180 16102
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15706 10732 16662
rect 10876 16662 10928 16668
rect 10782 16623 10838 16632
rect 10784 16040 10836 16046
rect 10980 16028 11008 18226
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11336 17876 11388 17882
rect 11336 17818 11388 17824
rect 11348 17202 11376 17818
rect 11440 17542 11468 18022
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11440 17270 11468 17478
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11256 16969 11284 17002
rect 11242 16960 11298 16969
rect 11242 16895 11298 16904
rect 11348 16794 11376 17138
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11336 16652 11388 16658
rect 11440 16640 11468 17206
rect 11388 16612 11468 16640
rect 11336 16594 11388 16600
rect 11440 16250 11468 16612
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 10980 16017 11100 16028
rect 10980 16008 11114 16017
rect 10980 16000 11058 16008
rect 10784 15982 10836 15988
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10336 15162 10364 15506
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10704 15094 10732 15642
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14006 10732 15030
rect 10796 14074 10824 15982
rect 10876 15972 10928 15978
rect 11058 15943 11114 15952
rect 10876 15914 10928 15920
rect 10888 15162 10916 15914
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10796 13530 10824 13738
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10796 13297 10824 13330
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10796 12918 10824 13223
rect 10784 12912 10836 12918
rect 10782 12880 10784 12889
rect 10836 12880 10838 12889
rect 10782 12815 10838 12824
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10704 12646 10732 12718
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12481 10732 12582
rect 10690 12472 10746 12481
rect 10690 12407 10746 12416
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10520 12186 10548 12242
rect 10520 12158 10732 12186
rect 10138 11928 10194 11937
rect 10138 11863 10194 11872
rect 10140 11688 10192 11694
rect 10046 11656 10102 11665
rect 10140 11630 10192 11636
rect 10046 11591 10102 11600
rect 9956 11552 10008 11558
rect 9862 11520 9918 11529
rect 9956 11494 10008 11500
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9862 11455 9918 11464
rect 9876 9722 9904 11455
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9876 8265 9904 9454
rect 9968 8537 9996 11494
rect 10060 11393 10088 11494
rect 10046 11384 10102 11393
rect 10046 11319 10102 11328
rect 10152 11082 10180 11630
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11218 10732 12158
rect 10782 12064 10838 12073
rect 10782 11999 10838 12008
rect 10796 11898 10824 11999
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10968 11212 11020 11218
rect 11072 11200 11100 15943
rect 11440 15706 11468 16186
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11440 14822 11468 15506
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11348 12918 11376 14758
rect 11440 14278 11468 14758
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11440 13326 11468 14214
rect 11532 13530 11560 18663
rect 12256 18634 12308 18640
rect 12268 18358 12296 18634
rect 12452 18426 12480 18702
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11900 16794 11928 17682
rect 12452 17338 12480 18362
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17814 12756 18090
rect 12912 17882 12940 18770
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11992 16674 12020 16934
rect 12544 16794 12572 17138
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12912 16726 12940 16934
rect 13096 16726 13124 17070
rect 11900 16646 12020 16674
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 11704 15360 11756 15366
rect 11624 15320 11704 15348
rect 11624 15026 11652 15320
rect 11704 15302 11756 15308
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 14618 11652 14962
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 14074 11744 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11716 13870 11744 14010
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11532 12986 11560 13466
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11808 12986 11836 13262
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11020 11172 11100 11200
rect 10968 11154 11020 11160
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10046 10976 10102 10985
rect 10046 10911 10102 10920
rect 10060 9110 10088 10911
rect 10152 10849 10180 11018
rect 10138 10840 10194 10849
rect 10704 10810 10732 11154
rect 10138 10775 10194 10784
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 10406
rect 10874 10296 10930 10305
rect 10692 10260 10744 10266
rect 10980 10266 11008 11154
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 10874 10231 10930 10240
rect 10968 10260 11020 10266
rect 10692 10202 10744 10208
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10152 8838 10180 10066
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 9602 10640 9862
rect 10704 9722 10732 10202
rect 10888 9761 10916 10231
rect 10968 10202 11020 10208
rect 11164 10169 11192 10474
rect 11150 10160 11206 10169
rect 11060 10124 11112 10130
rect 11150 10095 11206 10104
rect 11060 10066 11112 10072
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10874 9752 10930 9761
rect 10692 9716 10744 9722
rect 10874 9687 10930 9696
rect 10692 9658 10744 9664
rect 10612 9586 10732 9602
rect 10612 9580 10744 9586
rect 10612 9574 10692 9580
rect 10692 9522 10744 9528
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10704 9160 10732 9522
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10784 9376 10836 9382
rect 10782 9344 10784 9353
rect 10836 9344 10838 9353
rect 10782 9279 10838 9288
rect 10612 9132 10732 9160
rect 10612 9042 10640 9132
rect 10888 9110 10916 9454
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 9954 8528 10010 8537
rect 10336 8498 10364 8910
rect 10612 8634 10640 8978
rect 10692 8832 10744 8838
rect 10744 8792 10824 8820
rect 10692 8774 10744 8780
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 9954 8463 10010 8472
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10046 8392 10102 8401
rect 10046 8327 10102 8336
rect 9862 8256 9918 8265
rect 9862 8191 9918 8200
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 6934 9904 7686
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9876 5914 9904 6870
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9876 3777 9904 5714
rect 9968 4826 9996 5714
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9968 3942 9996 4082
rect 9956 3936 10008 3942
rect 9954 3904 9956 3913
rect 10008 3904 10010 3913
rect 9954 3839 10010 3848
rect 9862 3768 9918 3777
rect 10060 3738 10088 8327
rect 10690 8256 10746 8265
rect 10289 8188 10585 8208
rect 10690 8191 10746 8200
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8191
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10140 8016 10192 8022
rect 10138 7984 10140 7993
rect 10192 7984 10194 7993
rect 10138 7919 10194 7928
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7410 10180 7754
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10152 6322 10180 7346
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10690 6896 10746 6905
rect 10690 6831 10746 6840
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10508 6384 10560 6390
rect 10506 6352 10508 6361
rect 10560 6352 10562 6361
rect 10140 6316 10192 6322
rect 10612 6338 10640 6598
rect 10704 6458 10732 6831
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10612 6310 10732 6338
rect 10506 6287 10562 6296
rect 10140 6258 10192 6264
rect 10152 6118 10180 6258
rect 10704 6254 10732 6310
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5846 10180 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10152 5545 10180 5646
rect 10138 5536 10194 5545
rect 10138 5471 10194 5480
rect 10336 5273 10364 5646
rect 10322 5264 10378 5273
rect 10322 5199 10378 5208
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4049 10732 6190
rect 10796 5409 10824 8792
rect 10980 7002 11008 9930
rect 11072 9722 11100 10066
rect 11150 10024 11206 10033
rect 11150 9959 11152 9968
rect 11204 9959 11206 9968
rect 11152 9930 11204 9936
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 11072 8090 11100 9658
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11164 7886 11192 8434
rect 11256 8401 11284 12582
rect 11532 12374 11560 12922
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11518 12200 11574 12209
rect 11518 12135 11520 12144
rect 11572 12135 11574 12144
rect 11520 12106 11572 12112
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11348 9654 11376 10950
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11440 9586 11468 10610
rect 11532 10146 11560 11562
rect 11624 11286 11652 12650
rect 11702 11384 11758 11393
rect 11702 11319 11758 11328
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11624 10266 11652 10678
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11532 10118 11652 10146
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11348 8498 11376 9386
rect 11440 9178 11468 9522
rect 11532 9382 11560 9930
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11242 8392 11298 8401
rect 11242 8327 11298 8336
rect 11242 8120 11298 8129
rect 11242 8055 11298 8064
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7546 11192 7822
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11058 6896 11114 6905
rect 11058 6831 11060 6840
rect 11112 6831 11114 6840
rect 11060 6802 11112 6808
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10782 5400 10838 5409
rect 10782 5335 10838 5344
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10796 4865 10824 5102
rect 10782 4856 10838 4865
rect 10782 4791 10838 4800
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10796 4078 10824 4422
rect 10784 4072 10836 4078
rect 10690 4040 10746 4049
rect 10784 4014 10836 4020
rect 10690 3975 10746 3984
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10692 3936 10744 3942
rect 10796 3913 10824 4014
rect 10692 3878 10744 3884
rect 10782 3904 10838 3913
rect 9862 3703 9918 3712
rect 10048 3732 10100 3738
rect 9876 2854 9904 3703
rect 10048 3674 10100 3680
rect 10152 3505 10180 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3777 10732 3878
rect 10782 3839 10838 3848
rect 10690 3768 10746 3777
rect 10690 3703 10746 3712
rect 10784 3732 10836 3738
rect 10888 3720 10916 6054
rect 11072 5914 11100 6802
rect 11164 6662 11192 7482
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6186 11192 6598
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11164 5778 11192 6122
rect 11256 5914 11284 8055
rect 11440 8022 11468 9114
rect 11532 8498 11560 9318
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11440 7546 11468 7958
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11624 7154 11652 10118
rect 11716 9081 11744 11319
rect 11794 9888 11850 9897
rect 11794 9823 11850 9832
rect 11702 9072 11758 9081
rect 11702 9007 11758 9016
rect 11808 7698 11836 9823
rect 11440 7126 11652 7154
rect 11716 7670 11836 7698
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11348 6225 11376 6326
rect 11334 6216 11390 6225
rect 11334 6151 11390 6160
rect 11348 6118 11376 6151
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11164 4690 11192 5714
rect 11256 4758 11284 5850
rect 11334 5536 11390 5545
rect 11334 5471 11390 5480
rect 11348 5370 11376 5471
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10836 3692 10916 3720
rect 10784 3674 10836 3680
rect 10138 3496 10194 3505
rect 10138 3431 10194 3440
rect 9956 3392 10008 3398
rect 10888 3369 10916 3692
rect 10980 3505 11008 4490
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4049 11100 4422
rect 11164 4282 11192 4626
rect 11348 4593 11376 5306
rect 11334 4584 11390 4593
rect 11334 4519 11390 4528
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 9956 3334 10008 3340
rect 10874 3360 10930 3369
rect 9968 3233 9996 3334
rect 10874 3295 10930 3304
rect 9954 3224 10010 3233
rect 9954 3159 10010 3168
rect 11072 3097 11100 3878
rect 11164 3738 11192 4218
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11164 3194 11192 3674
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11058 3088 11114 3097
rect 11058 3023 11114 3032
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9692 2774 9812 2802
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9692 2650 9720 2774
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9034 2544 9090 2553
rect 9034 2479 9090 2488
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 8956 2400 9076 2428
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 2009 8800 2246
rect 8758 2000 8814 2009
rect 8758 1935 8814 1944
rect 8574 1456 8630 1465
rect 8574 1391 8630 1400
rect 9048 480 9076 2400
rect 9126 2408 9182 2417
rect 9126 2343 9128 2352
rect 9180 2343 9182 2352
rect 9128 2314 9180 2320
rect 10060 2281 10088 2450
rect 10046 2272 10102 2281
rect 10046 2207 10102 2216
rect 9588 604 9640 610
rect 9588 546 9640 552
rect 9600 480 9628 546
rect 10152 480 10180 2926
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10230 2544 10286 2553
rect 10704 2514 10732 2790
rect 10782 2680 10838 2689
rect 10782 2615 10838 2624
rect 10230 2479 10286 2488
rect 10692 2508 10744 2514
rect 10244 2446 10272 2479
rect 10692 2450 10744 2456
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10796 480 10824 2615
rect 11164 2446 11192 3130
rect 11334 3088 11390 3097
rect 11334 3023 11336 3032
rect 11388 3023 11390 3032
rect 11336 2994 11388 3000
rect 11440 2938 11468 7126
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11624 6390 11652 6938
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11716 5794 11744 7670
rect 11794 7576 11850 7585
rect 11794 7511 11850 7520
rect 11624 5766 11744 5794
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 5137 11560 5510
rect 11518 5128 11574 5137
rect 11518 5063 11574 5072
rect 11624 4842 11652 5766
rect 11704 5704 11756 5710
rect 11702 5672 11704 5681
rect 11756 5672 11758 5681
rect 11702 5607 11758 5616
rect 11808 5370 11836 7511
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11532 4814 11652 4842
rect 11532 3602 11560 4814
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11624 4282 11652 4694
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11348 2910 11468 2938
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11348 480 11376 2910
rect 11532 2582 11560 3538
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11624 2650 11652 2790
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11808 2514 11836 3062
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1601 11652 2246
rect 11610 1592 11666 1601
rect 11610 1527 11666 1536
rect 11900 480 11928 16646
rect 13174 16144 13230 16153
rect 13174 16079 13230 16088
rect 12898 16008 12954 16017
rect 12898 15943 12954 15952
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12360 14822 12388 14894
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11992 13870 12020 14418
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11992 11626 12020 13806
rect 12452 13734 12480 14350
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12162 13424 12218 13433
rect 12162 13359 12218 13368
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 12084 11354 12112 12242
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12176 10441 12204 13359
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12256 12640 12308 12646
rect 12254 12608 12256 12617
rect 12308 12608 12310 12617
rect 12254 12543 12310 12552
rect 12360 11898 12388 12786
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12452 11558 12480 13670
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12714 12664 13330
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12714 12336 12770 12345
rect 12714 12271 12770 12280
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10577 12296 10610
rect 12254 10568 12310 10577
rect 12254 10503 12310 10512
rect 12162 10432 12218 10441
rect 12162 10367 12218 10376
rect 12176 9518 12204 10367
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12268 9654 12296 10134
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11978 8528 12034 8537
rect 11978 8463 12034 8472
rect 11992 3126 12020 8463
rect 12176 8362 12204 8910
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12176 7857 12204 8298
rect 12162 7848 12218 7857
rect 12162 7783 12218 7792
rect 12070 7440 12126 7449
rect 12070 7375 12126 7384
rect 12084 4146 12112 7375
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 4758 12204 6938
rect 12268 6866 12296 8978
rect 12452 8945 12480 11222
rect 12544 10810 12572 11630
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12544 10470 12572 10542
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12530 9616 12586 9625
rect 12530 9551 12586 9560
rect 12544 9353 12572 9551
rect 12530 9344 12586 9353
rect 12530 9279 12586 9288
rect 12438 8936 12494 8945
rect 12438 8871 12494 8880
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8430 12388 8774
rect 12438 8528 12494 8537
rect 12438 8463 12494 8472
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12162 4312 12218 4321
rect 12162 4247 12218 4256
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12176 3369 12204 4247
rect 12268 3890 12296 6802
rect 12452 6066 12480 8463
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12544 8090 12572 8366
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12636 7954 12664 11494
rect 12728 11098 12756 12271
rect 12820 11937 12848 13126
rect 12806 11928 12862 11937
rect 12806 11863 12862 11872
rect 12806 11520 12862 11529
rect 12806 11455 12862 11464
rect 12820 11257 12848 11455
rect 12806 11248 12862 11257
rect 12806 11183 12862 11192
rect 12728 11070 12848 11098
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10606 12756 10950
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10266 12756 10542
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12820 10010 12848 11070
rect 12912 10742 12940 15943
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13004 15162 13032 15506
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 13004 14414 13032 14894
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14074 13032 14350
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12782 13124 13126
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12992 12640 13044 12646
rect 13188 12628 13216 16079
rect 12992 12582 13044 12588
rect 13096 12600 13216 12628
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12728 9982 12848 10010
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12452 6038 12572 6066
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12360 4978 12388 5306
rect 12452 5166 12480 5850
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12544 5098 12572 6038
rect 12622 5128 12678 5137
rect 12532 5092 12584 5098
rect 12622 5063 12678 5072
rect 12532 5034 12584 5040
rect 12636 5030 12664 5063
rect 12624 5024 12676 5030
rect 12360 4950 12572 4978
rect 12624 4966 12676 4972
rect 12438 3904 12494 3913
rect 12268 3862 12388 3890
rect 12360 3738 12388 3862
rect 12438 3839 12494 3848
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12268 3641 12296 3674
rect 12254 3632 12310 3641
rect 12254 3567 12310 3576
rect 12162 3360 12218 3369
rect 12162 3295 12218 3304
rect 12452 3194 12480 3839
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12164 2984 12216 2990
rect 12162 2952 12164 2961
rect 12360 2972 12388 3062
rect 12544 2990 12572 4950
rect 12728 4826 12756 9982
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9450 12848 9862
rect 12898 9616 12954 9625
rect 12898 9551 12954 9560
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 7041 12848 7142
rect 12806 7032 12862 7041
rect 12806 6967 12862 6976
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12820 5778 12848 6190
rect 12912 5817 12940 9551
rect 13004 8129 13032 12582
rect 13096 12238 13124 12600
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11354 13124 12174
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11801 13216 12038
rect 13174 11792 13230 11801
rect 13174 11727 13230 11736
rect 13174 11520 13230 11529
rect 13174 11455 13230 11464
rect 13188 11354 13216 11455
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13188 10810 13216 11154
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13174 10296 13230 10305
rect 13174 10231 13176 10240
rect 13228 10231 13230 10240
rect 13176 10202 13228 10208
rect 13188 9654 13216 10202
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8634 13124 8842
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12990 8120 13046 8129
rect 12990 8055 13046 8064
rect 13096 7970 13124 8570
rect 13188 8090 13216 8978
rect 13280 8090 13308 22607
rect 13740 20398 13768 23310
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13464 19718 13492 20334
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13464 19174 13492 19654
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13372 17202 13400 17478
rect 13464 17270 13492 19110
rect 13832 18630 13860 19178
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13832 18086 13860 18566
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 16250 13400 16526
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13372 16153 13400 16186
rect 13358 16144 13414 16153
rect 13358 16079 13414 16088
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15609 13400 15846
rect 13358 15600 13414 15609
rect 13358 15535 13414 15544
rect 13464 14822 13492 17206
rect 13556 16794 13584 17682
rect 13832 17610 13860 18022
rect 13924 17746 13952 18702
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 14016 17134 14044 17614
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 16114 13676 16390
rect 13832 16266 13860 16934
rect 14108 16794 14136 26250
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 17882 14688 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 23216 19281 23244 27520
rect 24766 27503 24822 27512
rect 24030 26888 24086 26897
rect 24030 26823 24086 26832
rect 23662 22672 23718 22681
rect 23662 22607 23718 22616
rect 23676 22574 23704 22607
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23478 20088 23534 20097
rect 23478 20023 23534 20032
rect 14830 19272 14886 19281
rect 14830 19207 14886 19216
rect 23202 19272 23258 19281
rect 23202 19207 23258 19216
rect 14844 19174 14872 19207
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14844 18834 14872 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 22834 18864 22890 18873
rect 14832 18828 14884 18834
rect 22834 18799 22890 18808
rect 14832 18770 14884 18776
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 22650 18048 22706 18057
rect 19622 17980 19918 18000
rect 22650 17983 22706 17992
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14660 17202 14688 17818
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15658 17232 15714 17241
rect 14648 17196 14700 17202
rect 15658 17167 15714 17176
rect 14648 17138 14700 17144
rect 14660 16794 14688 17138
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13740 16238 13860 16266
rect 14016 16250 14044 16662
rect 14660 16590 14688 16730
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14004 16244 14056 16250
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 15706 13676 16050
rect 13740 16046 13768 16238
rect 14004 16186 14056 16192
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 14660 15978 14688 16526
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13634 15464 13690 15473
rect 13634 15399 13636 15408
rect 13688 15399 13690 15408
rect 13636 15370 13688 15376
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 13734 13492 14758
rect 13740 14618 13768 15642
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13832 15162 13860 15574
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 14568 14958 14596 15846
rect 14660 15502 14688 15914
rect 14844 15638 14872 17002
rect 15476 16992 15528 16998
rect 15528 16952 15608 16980
rect 15476 16934 15528 16940
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 15978 15332 16526
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16046 15516 16390
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 15488 15570 15516 15982
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13634 14512 13690 14521
rect 13634 14447 13690 14456
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13372 10146 13400 12650
rect 13464 11694 13492 13670
rect 13648 13530 13676 14447
rect 13832 13870 13860 14758
rect 13924 14618 13952 14826
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 13820 13864 13872 13870
rect 14384 13841 14412 14214
rect 13820 13806 13872 13812
rect 14370 13832 14426 13841
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13832 13462 13860 13806
rect 14370 13767 14426 13776
rect 14660 13462 14688 14418
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13870 14780 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14832 13728 14884 13734
rect 14738 13696 14794 13705
rect 14832 13670 14884 13676
rect 14738 13631 14794 13640
rect 13820 13456 13872 13462
rect 14648 13456 14700 13462
rect 13820 13398 13872 13404
rect 14646 13424 14648 13433
rect 14700 13424 14702 13433
rect 13832 13138 13860 13398
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14556 13388 14608 13394
rect 14646 13359 14702 13368
rect 14556 13330 14608 13336
rect 13832 13110 13952 13138
rect 13726 13016 13782 13025
rect 13726 12951 13782 12960
rect 13820 12980 13872 12986
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13542 12472 13598 12481
rect 13542 12407 13598 12416
rect 13556 12306 13584 12407
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13556 11898 13584 12242
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13544 10192 13596 10198
rect 13372 10118 13492 10146
rect 13544 10134 13596 10140
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13372 9722 13400 9998
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13372 9489 13400 9658
rect 13358 9480 13414 9489
rect 13358 9415 13414 9424
rect 13464 8922 13492 10118
rect 13372 8894 13492 8922
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13004 7942 13124 7970
rect 13004 7750 13032 7942
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 6905 13032 7686
rect 13188 7410 13216 8026
rect 13372 7698 13400 8894
rect 13450 8800 13506 8809
rect 13450 8735 13506 8744
rect 13280 7670 13400 7698
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12990 6896 13046 6905
rect 12990 6831 13046 6840
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12898 5808 12954 5817
rect 12808 5772 12860 5778
rect 12898 5743 12954 5752
rect 12808 5714 12860 5720
rect 12820 5370 12848 5714
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12216 2952 12388 2972
rect 12218 2944 12388 2952
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12162 2887 12218 2896
rect 12636 2802 12664 4694
rect 12452 2774 12664 2802
rect 12452 2666 12480 2774
rect 12452 2638 12572 2666
rect 12544 480 12572 2638
rect 12728 2582 12756 4762
rect 12912 4457 12940 5034
rect 12898 4448 12954 4457
rect 12898 4383 12954 4392
rect 12912 4078 12940 4383
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 13004 3754 13032 6394
rect 13096 4622 13124 7210
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13188 5302 13216 5782
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13096 3942 13124 4558
rect 13188 4486 13216 5238
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4214 13216 4422
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13176 3936 13228 3942
rect 13280 3913 13308 7670
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13372 7002 13400 7482
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6497 13400 6734
rect 13358 6488 13414 6497
rect 13358 6423 13360 6432
rect 13412 6423 13414 6432
rect 13360 6394 13412 6400
rect 13464 4434 13492 8735
rect 13556 5914 13584 10134
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 5545 13676 12718
rect 13740 11218 13768 12951
rect 13820 12922 13872 12928
rect 13832 12374 13860 12922
rect 13924 12850 13952 13110
rect 14016 12986 14044 13330
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13924 12442 13952 12786
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13924 11694 13952 12174
rect 14002 11928 14058 11937
rect 14002 11863 14058 11872
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 10470 13768 11154
rect 13924 11150 13952 11630
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10810 13952 11086
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9586 13768 9862
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13740 8945 13768 8978
rect 13726 8936 13782 8945
rect 13726 8871 13782 8880
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13740 8265 13768 8774
rect 13726 8256 13782 8265
rect 13726 8191 13782 8200
rect 13740 8090 13768 8191
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13832 6882 13860 8774
rect 13910 8392 13966 8401
rect 13910 8327 13966 8336
rect 13740 6854 13860 6882
rect 13740 6662 13768 6854
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13728 6112 13780 6118
rect 13726 6080 13728 6089
rect 13780 6080 13782 6089
rect 13726 6015 13782 6024
rect 13634 5536 13690 5545
rect 13634 5471 13690 5480
rect 13542 5400 13598 5409
rect 13542 5335 13544 5344
rect 13596 5335 13598 5344
rect 13544 5306 13596 5312
rect 13832 5166 13860 6854
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13648 4554 13676 5034
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13832 4554 13860 4694
rect 13924 4690 13952 8327
rect 14016 6866 14044 11863
rect 14108 11558 14136 12718
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 7954 14136 9862
rect 14200 8344 14228 12242
rect 14568 12238 14596 13330
rect 14646 13152 14702 13161
rect 14646 13087 14702 13096
rect 14660 12753 14688 13087
rect 14646 12744 14702 12753
rect 14646 12679 14702 12688
rect 14752 12345 14780 13631
rect 14844 13326 14872 13670
rect 15120 13530 15148 13874
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14844 12850 14872 13262
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15474 12880 15530 12889
rect 14832 12844 14884 12850
rect 15474 12815 15530 12824
rect 14832 12786 14884 12792
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15304 12442 15332 12650
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 14738 12336 14794 12345
rect 14738 12271 14794 12280
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14568 12073 14596 12174
rect 14554 12064 14610 12073
rect 14554 11999 14610 12008
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14292 11150 14320 11562
rect 14660 11354 14688 11630
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 9217 14320 9318
rect 14278 9208 14334 9217
rect 14278 9143 14334 9152
rect 14200 8316 14320 8344
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14200 7546 14228 7822
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14292 6984 14320 8316
rect 14200 6956 14320 6984
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6254 14044 6666
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14016 5914 14044 6190
rect 14108 6186 14136 6598
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 14016 4826 14044 5850
rect 14108 5370 14136 6122
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13464 4406 13676 4434
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13176 3878 13228 3884
rect 13266 3904 13322 3913
rect 13004 3726 13124 3754
rect 13188 3738 13216 3878
rect 13266 3839 13322 3848
rect 13358 3768 13414 3777
rect 12898 3224 12954 3233
rect 12898 3159 12954 3168
rect 12912 3058 12940 3159
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 13096 480 13124 3726
rect 13176 3732 13228 3738
rect 13464 3738 13492 4082
rect 13358 3703 13360 3712
rect 13176 3674 13228 3680
rect 13412 3703 13414 3712
rect 13452 3732 13504 3738
rect 13360 3674 13412 3680
rect 13452 3674 13504 3680
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13556 3194 13584 3402
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13648 480 13676 4406
rect 13924 4282 13952 4626
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13832 2854 13860 3470
rect 14108 3194 14136 5306
rect 14200 4282 14228 6956
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14292 3641 14320 6802
rect 14278 3632 14334 3641
rect 14278 3567 14334 3576
rect 14278 3360 14334 3369
rect 14278 3295 14334 3304
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14292 480 14320 3295
rect 14384 1034 14412 10406
rect 14476 3777 14504 10406
rect 14556 9920 14608 9926
rect 14752 9897 14780 11766
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 11218 15056 11494
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10810 15332 11086
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14556 9862 14608 9868
rect 14738 9888 14794 9897
rect 14568 9586 14596 9862
rect 14738 9823 14794 9832
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14844 9518 14872 9998
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14844 9178 14872 9454
rect 15028 9178 15056 9522
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 14830 9072 14886 9081
rect 14830 9007 14886 9016
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14752 8430 14780 8910
rect 14740 8424 14792 8430
rect 14844 8401 14872 9007
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14740 8366 14792 8372
rect 14830 8392 14886 8401
rect 14752 8090 14780 8366
rect 15304 8362 15332 9114
rect 14830 8327 14886 8336
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14568 4826 14596 7890
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14660 7342 14688 7686
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14660 6458 14688 7278
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14660 5234 14688 6394
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14752 5166 14780 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15120 6769 15148 6870
rect 14830 6760 14886 6769
rect 14830 6695 14886 6704
rect 15106 6760 15162 6769
rect 15106 6695 15162 6704
rect 14844 5914 14872 6695
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15290 6216 15346 6225
rect 15290 6151 15346 6160
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14752 4146 14780 4422
rect 14844 4196 14872 4626
rect 15014 4584 15070 4593
rect 15014 4519 15016 4528
rect 15068 4519 15070 4528
rect 15016 4490 15068 4496
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14844 4168 14964 4196
rect 14740 4140 14792 4146
rect 14792 4100 14872 4128
rect 14740 4082 14792 4088
rect 14646 4040 14702 4049
rect 14646 3975 14702 3984
rect 14660 3942 14688 3975
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14462 3768 14518 3777
rect 14462 3703 14518 3712
rect 14660 3670 14688 3878
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 1329 14596 3334
rect 14844 2990 14872 4100
rect 14936 3738 14964 4168
rect 15304 4078 15332 6151
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15290 3904 15346 3913
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15028 3466 15056 3878
rect 15290 3839 15346 3848
rect 15304 3738 15332 3839
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 14752 2650 14780 2926
rect 15028 2689 15056 2926
rect 15014 2680 15070 2689
rect 14740 2644 14792 2650
rect 15014 2615 15070 2624
rect 14740 2586 14792 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14554 1320 14610 1329
rect 14554 1255 14610 1264
rect 14384 1006 14872 1034
rect 14844 480 14872 1006
rect 15396 480 15424 12582
rect 15488 11558 15516 12815
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15488 8294 15516 9046
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 7478 15516 8230
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15580 7256 15608 16952
rect 15672 15706 15700 17167
rect 17682 16960 17738 16969
rect 17682 16895 17738 16904
rect 16210 16280 16266 16289
rect 16210 16215 16266 16224
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15844 15632 15896 15638
rect 15750 15600 15806 15609
rect 15844 15574 15896 15580
rect 15750 15535 15806 15544
rect 15658 15464 15714 15473
rect 15658 15399 15714 15408
rect 15672 14550 15700 15399
rect 15764 14550 15792 15535
rect 15856 15065 15884 15574
rect 15842 15056 15898 15065
rect 15842 14991 15898 15000
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15672 13938 15700 14486
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15764 13530 15792 14486
rect 15856 14346 15884 14991
rect 15948 14890 15976 15846
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 16040 15162 16068 15642
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15948 14414 15976 14826
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15948 14074 15976 14350
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16040 13954 16068 15098
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16132 14006 16160 14418
rect 16120 14000 16172 14006
rect 15948 13926 16068 13954
rect 16118 13968 16120 13977
rect 16172 13968 16174 13977
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 12986 15792 13194
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15856 12646 15884 13262
rect 15844 12640 15896 12646
rect 15658 12608 15714 12617
rect 15844 12582 15896 12588
rect 15658 12543 15714 12552
rect 15672 9654 15700 12543
rect 15856 12238 15884 12582
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15764 10266 15792 10542
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15948 9353 15976 13926
rect 16118 13903 16174 13912
rect 16224 13852 16252 16215
rect 17130 16008 17186 16017
rect 17130 15943 17186 15952
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16500 15178 16528 15302
rect 16500 15150 16712 15178
rect 16684 15026 16712 15150
rect 16672 15020 16724 15026
rect 16316 14958 16344 14989
rect 16672 14962 16724 14968
rect 16304 14952 16356 14958
rect 16302 14920 16304 14929
rect 16356 14920 16358 14929
rect 16302 14855 16358 14864
rect 16486 14920 16542 14929
rect 16486 14855 16542 14864
rect 16316 14550 16344 14855
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 16304 14000 16356 14006
rect 16302 13968 16304 13977
rect 16356 13968 16358 13977
rect 16302 13903 16358 13912
rect 16040 13824 16252 13852
rect 16040 12753 16068 13824
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16316 12986 16344 13738
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16026 12744 16082 12753
rect 16026 12679 16082 12688
rect 16040 12442 16068 12679
rect 16118 12608 16174 12617
rect 16118 12543 16174 12552
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 16040 11762 16068 12378
rect 16132 11898 16160 12543
rect 16408 12345 16436 14758
rect 16500 12782 16528 14855
rect 16684 14278 16712 14962
rect 16776 14521 16804 15302
rect 16762 14512 16818 14521
rect 16762 14447 16818 14456
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 13841 16712 14214
rect 16776 13938 16804 14447
rect 16854 14376 16910 14385
rect 16854 14311 16856 14320
rect 16908 14311 16910 14320
rect 16856 14282 16908 14288
rect 17052 14113 17080 15302
rect 17038 14104 17094 14113
rect 17038 14039 17094 14048
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16670 13832 16726 13841
rect 16670 13767 16726 13776
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16762 13152 16818 13161
rect 16762 13087 16818 13096
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16592 12442 16620 12718
rect 16776 12646 16804 13087
rect 16960 12850 16988 13330
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16854 12744 16910 12753
rect 16854 12679 16910 12688
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16394 12336 16450 12345
rect 16394 12271 16450 12280
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16776 11558 16804 12174
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16132 10266 16160 11154
rect 16408 10713 16436 11494
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16394 10704 16450 10713
rect 16394 10639 16450 10648
rect 16500 10606 16528 11290
rect 16776 10810 16804 11494
rect 16868 11354 16896 12679
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16868 11014 16896 11045
rect 16856 11008 16908 11014
rect 16854 10976 16856 10985
rect 16908 10976 16910 10985
rect 16854 10911 16910 10920
rect 16868 10810 16896 10911
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16132 9382 16160 9522
rect 16488 9512 16540 9518
rect 16592 9500 16620 9862
rect 16670 9752 16726 9761
rect 16670 9687 16726 9696
rect 16540 9472 16620 9500
rect 16488 9454 16540 9460
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16120 9376 16172 9382
rect 15934 9344 15990 9353
rect 16120 9318 16172 9324
rect 15934 9279 15990 9288
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15856 7342 15884 8978
rect 15948 8673 15976 9279
rect 15934 8664 15990 8673
rect 15934 8599 15990 8608
rect 16132 8566 16160 9318
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 16040 7274 16068 7890
rect 16028 7268 16080 7274
rect 15580 7228 15792 7256
rect 15566 7168 15622 7177
rect 15566 7103 15622 7112
rect 15580 6866 15608 7103
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 4049 15516 5510
rect 15474 4040 15530 4049
rect 15474 3975 15530 3984
rect 15566 3768 15622 3777
rect 15566 3703 15568 3712
rect 15620 3703 15622 3712
rect 15568 3674 15620 3680
rect 15580 2990 15608 3674
rect 15764 3074 15792 7228
rect 16028 7210 16080 7216
rect 15934 6896 15990 6905
rect 15934 6831 15990 6840
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 6186 15884 6734
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15856 5778 15884 6122
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15856 3534 15884 5034
rect 15948 4622 15976 6831
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16040 3913 16068 7210
rect 16132 6866 16160 8502
rect 16316 7546 16344 9386
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 8090 16620 8298
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16684 7954 16712 9687
rect 16960 9382 16988 10066
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16684 7546 16712 7890
rect 16854 7848 16910 7857
rect 16854 7783 16910 7792
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16670 7440 16726 7449
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16132 5914 16160 6802
rect 16224 6662 16252 7210
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16224 4282 16252 6598
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16026 3904 16082 3913
rect 16026 3839 16082 3848
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 3194 15884 3470
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15764 3046 16068 3074
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 16040 480 16068 3046
rect 16224 2417 16252 4014
rect 16210 2408 16266 2417
rect 16210 2343 16266 2352
rect 16316 1737 16344 6122
rect 16408 4146 16436 7414
rect 16670 7375 16726 7384
rect 16684 7342 16712 7375
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16670 6488 16726 6497
rect 16670 6423 16726 6432
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16500 5386 16528 6054
rect 16592 5914 16620 6190
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16500 5358 16620 5386
rect 16488 5296 16540 5302
rect 16486 5264 16488 5273
rect 16540 5264 16542 5273
rect 16486 5199 16542 5208
rect 16592 4758 16620 5358
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16408 3738 16436 4082
rect 16684 4010 16712 6423
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16776 5370 16804 5714
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16868 4078 16896 7783
rect 16960 4214 16988 9318
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17052 8090 17080 9114
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17052 7410 17080 8026
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17052 5846 17080 6258
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 17052 4690 17080 5782
rect 17144 4826 17172 15943
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17236 9489 17264 14826
rect 17328 14822 17356 15506
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17328 14618 17356 14758
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17316 14408 17368 14414
rect 17314 14376 17316 14385
rect 17368 14376 17370 14385
rect 17314 14311 17370 14320
rect 17328 14074 17356 14311
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17314 13016 17370 13025
rect 17314 12951 17370 12960
rect 17328 10266 17356 12951
rect 17420 12782 17448 14758
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17512 13190 17540 13874
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17512 12306 17540 13126
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17512 11898 17540 12242
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17604 10792 17632 13806
rect 17512 10764 17632 10792
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17328 9722 17356 10202
rect 17420 10062 17448 10406
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17222 9480 17278 9489
rect 17222 9415 17278 9424
rect 17236 8537 17264 9415
rect 17420 9178 17448 9998
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17222 8528 17278 8537
rect 17222 8463 17278 8472
rect 17314 7984 17370 7993
rect 17314 7919 17370 7928
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 17130 4040 17186 4049
rect 16672 4004 16724 4010
rect 17130 3975 17186 3984
rect 16672 3946 16724 3952
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16854 3632 16910 3641
rect 16854 3567 16856 3576
rect 16908 3567 16910 3576
rect 16856 3538 16908 3544
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17052 3233 17080 3334
rect 17038 3224 17094 3233
rect 17038 3159 17094 3168
rect 16854 2680 16910 2689
rect 16854 2615 16856 2624
rect 16908 2615 16910 2624
rect 16856 2586 16908 2592
rect 16302 1728 16358 1737
rect 16302 1663 16358 1672
rect 16578 1592 16634 1601
rect 16578 1527 16634 1536
rect 16592 480 16620 1527
rect 17144 480 17172 3975
rect 17236 3738 17264 4762
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17328 3670 17356 7919
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6458 17448 6598
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17512 6361 17540 10764
rect 17590 10704 17646 10713
rect 17590 10639 17646 10648
rect 17604 7546 17632 10639
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17696 6905 17724 16895
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 18052 16040 18104 16046
rect 18050 16008 18052 16017
rect 18104 16008 18106 16017
rect 18050 15943 18106 15952
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 10198 17816 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20810 15600 20866 15609
rect 18236 15564 18288 15570
rect 18236 15506 18288 15512
rect 19340 15564 19392 15570
rect 20810 15535 20866 15544
rect 19340 15506 19392 15512
rect 18248 14822 18276 15506
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 14006 17908 14214
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17880 13530 17908 13942
rect 18052 13728 18104 13734
rect 18248 13682 18276 14758
rect 18052 13670 18104 13676
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 18064 12442 18092 13670
rect 18156 13654 18276 13682
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17972 11762 18000 12038
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 11688 17920 11694
rect 18156 11642 18184 13654
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 17868 11630 17920 11636
rect 17880 11558 17908 11630
rect 17972 11614 18184 11642
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 10470 17908 11494
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17972 9704 18000 11614
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17788 9676 18000 9704
rect 17788 8090 17816 9676
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8634 17908 8910
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17972 8430 18000 9454
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17776 8084 17828 8090
rect 17880 8072 17908 8298
rect 17960 8084 18012 8090
rect 17880 8044 17960 8072
rect 17776 8026 17828 8032
rect 17960 8026 18012 8032
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7206 18000 7890
rect 18064 7342 18092 11494
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18156 10470 18184 10542
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 10146 18184 10406
rect 18248 10266 18276 13466
rect 18340 12356 18368 15302
rect 19352 14958 19380 15506
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 18512 14952 18564 14958
rect 19340 14952 19392 14958
rect 18512 14894 18564 14900
rect 19168 14900 19340 14906
rect 19168 14894 19392 14900
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13734 18460 14214
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18432 12458 18460 13670
rect 18524 13530 18552 14894
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 19168 14878 19380 14894
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18616 14521 18644 14554
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12889 18552 13126
rect 18510 12880 18566 12889
rect 18510 12815 18512 12824
rect 18564 12815 18566 12824
rect 18512 12786 18564 12792
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18524 12617 18552 12650
rect 18510 12608 18566 12617
rect 18510 12543 18566 12552
rect 18432 12430 18552 12458
rect 18340 12328 18460 12356
rect 18326 11112 18382 11121
rect 18326 11047 18382 11056
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18156 10118 18276 10146
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9518 18184 9862
rect 18248 9722 18276 10118
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18156 8650 18184 9454
rect 18340 8974 18368 11047
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18156 8634 18276 8650
rect 18156 8628 18288 8634
rect 18156 8622 18236 8628
rect 18156 7886 18184 8622
rect 18236 8570 18288 8576
rect 18340 8362 18368 8774
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18340 7818 18368 8298
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18432 7585 18460 12328
rect 18524 11286 18552 12430
rect 18616 12102 18644 13262
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18616 11801 18644 12038
rect 18602 11792 18658 11801
rect 18602 11727 18658 11736
rect 18708 11354 18736 12378
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18524 9110 18552 11086
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18616 10266 18644 10950
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18616 9178 18644 10202
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18524 8090 18552 9046
rect 18800 8090 18828 14826
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19076 14074 19104 14418
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18418 7576 18474 7585
rect 18418 7511 18474 7520
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17960 7200 18012 7206
rect 17958 7168 17960 7177
rect 18012 7168 18014 7177
rect 17958 7103 18014 7112
rect 18064 7002 18092 7278
rect 18892 7154 18920 12310
rect 18984 11529 19012 13330
rect 19062 12336 19118 12345
rect 19062 12271 19064 12280
rect 19116 12271 19118 12280
rect 19064 12242 19116 12248
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11830 19104 12038
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 18970 11520 19026 11529
rect 18970 11455 19026 11464
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18984 7274 19012 11222
rect 19062 8936 19118 8945
rect 19062 8871 19118 8880
rect 19076 8537 19104 8871
rect 19062 8528 19118 8537
rect 19062 8463 19118 8472
rect 18972 7268 19024 7274
rect 18972 7210 19024 7216
rect 18800 7126 18920 7154
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17682 6896 17738 6905
rect 17682 6831 17738 6840
rect 18144 6860 18196 6866
rect 17498 6352 17554 6361
rect 17498 6287 17554 6296
rect 17512 6186 17540 6287
rect 17696 6254 17724 6831
rect 18144 6802 18196 6808
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5370 17816 6122
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17420 3738 17448 4694
rect 17512 4622 17540 5034
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17512 4282 17540 4558
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17316 3664 17368 3670
rect 17222 3632 17278 3641
rect 17316 3606 17368 3612
rect 17222 3567 17278 3576
rect 17236 2854 17264 3567
rect 17328 3194 17356 3606
rect 17788 3194 17816 5306
rect 17868 4820 17920 4826
rect 17972 4808 18000 6598
rect 18156 6254 18184 6802
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5166 18184 5510
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 17920 4780 18000 4808
rect 17868 4762 17920 4768
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 17972 4282 18000 4422
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17972 3738 18000 4218
rect 18708 4146 18736 4422
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18708 3738 18736 4082
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18512 3528 18564 3534
rect 18142 3496 18198 3505
rect 18512 3470 18564 3476
rect 18142 3431 18144 3440
rect 18196 3431 18198 3440
rect 18144 3402 18196 3408
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 18064 2650 18092 2994
rect 18156 2990 18184 3402
rect 18326 3360 18382 3369
rect 18326 3295 18382 3304
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17774 2000 17830 2009
rect 17774 1935 17830 1944
rect 17788 480 17816 1935
rect 18340 480 18368 3295
rect 18524 2650 18552 3470
rect 18708 3194 18736 3674
rect 18800 3398 18828 7126
rect 18878 7032 18934 7041
rect 18878 6967 18880 6976
rect 18932 6967 18934 6976
rect 18880 6938 18932 6944
rect 18892 5914 18920 6938
rect 19076 6882 19104 8463
rect 18984 6854 19104 6882
rect 18984 6798 19012 6854
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18984 6390 19012 6734
rect 19076 6458 19104 6734
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18972 6384 19024 6390
rect 18972 6326 19024 6332
rect 18970 6080 19026 6089
rect 18970 6015 19026 6024
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18984 4672 19012 6015
rect 19062 5672 19118 5681
rect 19062 5607 19118 5616
rect 19076 4826 19104 5607
rect 19168 4826 19196 14878
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19260 12374 19288 13874
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11393 19288 12038
rect 19246 11384 19302 11393
rect 19246 11319 19302 11328
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19260 10146 19288 10746
rect 19352 10266 19380 14758
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19260 10118 19380 10146
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19260 8974 19288 9318
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19246 8392 19302 8401
rect 19246 8327 19248 8336
rect 19300 8327 19302 8336
rect 19248 8298 19300 8304
rect 19260 7954 19288 8298
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19260 7410 19288 7890
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19352 6934 19380 10118
rect 19444 9042 19472 15302
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 13938 19564 14418
rect 19614 13968 19670 13977
rect 19524 13932 19576 13938
rect 19614 13903 19670 13912
rect 19524 13874 19576 13880
rect 19628 13870 19656 13903
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20088 12850 20116 13466
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19522 12744 19578 12753
rect 19522 12679 19524 12688
rect 19576 12679 19578 12688
rect 19524 12650 19576 12656
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19982 11792 20038 11801
rect 19982 11727 20038 11736
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19536 11014 19564 11562
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19706 11248 19762 11257
rect 19616 11212 19668 11218
rect 19996 11218 20024 11727
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19706 11183 19708 11192
rect 19616 11154 19668 11160
rect 19760 11183 19762 11192
rect 19984 11212 20036 11218
rect 19708 11154 19760 11160
rect 19984 11154 20036 11160
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19536 10470 19564 10950
rect 19628 10810 19656 11154
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 10062 19564 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19996 10198 20024 11154
rect 20088 11150 20116 11494
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19524 10056 19576 10062
rect 19812 10033 19840 10066
rect 19524 9998 19576 10004
rect 19798 10024 19854 10033
rect 19536 9722 19564 9998
rect 19798 9959 19854 9968
rect 19982 10024 20038 10033
rect 19982 9959 19984 9968
rect 20036 9959 20038 9968
rect 19984 9930 20036 9936
rect 20088 9926 20116 11086
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20180 9194 20208 14758
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20442 13288 20498 13297
rect 20442 13223 20498 13232
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 12442 20300 12718
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20364 11121 20392 11562
rect 20456 11286 20484 13223
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20548 11121 20576 14214
rect 20824 13569 20852 15535
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 21822 15328 21878 15337
rect 21822 15263 21878 15272
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20810 13560 20866 13569
rect 20810 13495 20866 13504
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20732 11694 20760 12242
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20732 11150 20760 11630
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20720 11144 20772 11150
rect 20350 11112 20406 11121
rect 20350 11047 20406 11056
rect 20534 11112 20590 11121
rect 20534 11047 20590 11056
rect 20640 11104 20720 11132
rect 20640 10538 20668 11104
rect 20720 11086 20772 11092
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10606 20760 10950
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20732 10266 20760 10542
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20352 9920 20404 9926
rect 20352 9862 20404 9868
rect 20364 9722 20392 9862
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20548 9518 20576 10202
rect 20824 9625 20852 11494
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20536 9512 20588 9518
rect 20720 9512 20772 9518
rect 20536 9454 20588 9460
rect 20718 9480 20720 9489
rect 20772 9480 20774 9489
rect 20718 9415 20774 9424
rect 20088 9166 20208 9194
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19536 8090 19564 8842
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19614 7576 19670 7585
rect 19720 7546 19748 7822
rect 19614 7511 19670 7520
rect 19708 7540 19760 7546
rect 19628 7342 19656 7511
rect 19708 7482 19760 7488
rect 19812 7478 19840 7822
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19616 6928 19668 6934
rect 19616 6870 19668 6876
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19338 6352 19394 6361
rect 19394 6310 19472 6338
rect 19338 6287 19394 6296
rect 19340 6248 19392 6254
rect 19338 6216 19340 6225
rect 19392 6216 19394 6225
rect 19338 6151 19394 6160
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 18892 4644 19012 4672
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18708 2582 18736 3130
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18892 480 18920 4644
rect 18972 4548 19024 4554
rect 18972 4490 19024 4496
rect 18984 3942 19012 4490
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 4066 368 4122 377
rect 4066 303 4122 312
rect 4342 0 4398 480
rect 4894 0 4950 480
rect 5538 0 5594 480
rect 6090 0 6146 480
rect 6642 0 6698 480
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 9034 0 9090 480
rect 9586 0 9642 480
rect 10138 0 10194 480
rect 10782 0 10838 480
rect 11334 0 11390 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17774 0 17830 480
rect 18326 0 18382 480
rect 18878 0 18934 480
rect 18984 377 19012 3878
rect 19260 2961 19288 6054
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 4826 19380 5510
rect 19444 5284 19472 6310
rect 19536 6186 19564 6598
rect 19628 6186 19656 6870
rect 19996 6202 20024 8774
rect 20088 6866 20116 9166
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 20180 8634 20208 9046
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20442 8664 20498 8673
rect 20168 8628 20220 8634
rect 20442 8599 20498 8608
rect 20168 8570 20220 8576
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20168 7336 20220 7342
rect 20166 7304 20168 7313
rect 20220 7304 20222 7313
rect 20166 7239 20222 7248
rect 20272 7002 20300 7482
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19616 6180 19668 6186
rect 19996 6174 20208 6202
rect 19616 6122 19668 6128
rect 19536 5642 19564 6122
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 19628 5681 19656 5714
rect 19614 5672 19670 5681
rect 19524 5636 19576 5642
rect 19614 5607 19670 5616
rect 19524 5578 19576 5584
rect 19524 5296 19576 5302
rect 19444 5256 19524 5284
rect 19524 5238 19576 5244
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19430 4856 19486 4865
rect 19340 4820 19392 4826
rect 19622 4848 19918 4868
rect 19430 4791 19486 4800
rect 19340 4762 19392 4768
rect 19352 3738 19380 4762
rect 19444 4690 19472 4791
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19432 3936 19484 3942
rect 19430 3904 19432 3913
rect 19484 3904 19486 3913
rect 19430 3839 19486 3848
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19536 3670 19564 4694
rect 19800 4616 19852 4622
rect 19996 4604 20024 6054
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20088 5370 20116 5850
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20074 5128 20130 5137
rect 20074 5063 20130 5072
rect 19852 4576 20024 4604
rect 19800 4558 19852 4564
rect 19812 4282 19840 4558
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19522 3088 19578 3097
rect 19522 3023 19578 3032
rect 19246 2952 19302 2961
rect 19246 2887 19302 2896
rect 19430 2952 19486 2961
rect 19430 2887 19486 2896
rect 19444 678 19472 2887
rect 19432 672 19484 678
rect 19432 614 19484 620
rect 19536 480 19564 3023
rect 19904 2961 19932 3334
rect 19890 2952 19946 2961
rect 19890 2887 19946 2896
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20088 480 20116 5063
rect 20180 610 20208 6174
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20272 4185 20300 4966
rect 20258 4176 20314 4185
rect 20258 4111 20314 4120
rect 20364 3777 20392 7142
rect 20456 5914 20484 8599
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20640 8090 20668 8366
rect 20732 8362 20760 8774
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20732 7886 20760 8298
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20824 7886 20852 8026
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20824 7546 20852 7822
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 6118 20668 6802
rect 20824 6798 20852 7482
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20824 6458 20852 6734
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 5914 20668 6054
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20640 5234 20668 5510
rect 20810 5264 20866 5273
rect 20628 5228 20680 5234
rect 20810 5199 20866 5208
rect 20628 5170 20680 5176
rect 20824 5098 20852 5199
rect 20812 5092 20864 5098
rect 20812 5034 20864 5040
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4826 20576 4966
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20824 4690 20852 5034
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20350 3768 20406 3777
rect 20350 3703 20406 3712
rect 20640 3346 20668 4082
rect 20810 4040 20866 4049
rect 20810 3975 20866 3984
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 3534 20760 3878
rect 20824 3670 20852 3975
rect 20916 3738 20944 13806
rect 21468 13734 21496 14418
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11830 21036 12038
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 21008 10985 21036 11766
rect 21088 11552 21140 11558
rect 21086 11520 21088 11529
rect 21140 11520 21142 11529
rect 21086 11455 21142 11464
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20994 10976 21050 10985
rect 20994 10911 21050 10920
rect 21100 10674 21128 11290
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21086 10160 21142 10169
rect 21086 10095 21142 10104
rect 21100 10062 21128 10095
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 21100 9722 21128 9998
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21008 4185 21036 9318
rect 21192 9058 21220 13262
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 10266 21312 12174
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21284 9722 21312 10202
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21376 9602 21404 12582
rect 21468 10810 21496 13670
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21284 9574 21404 9602
rect 21284 9110 21312 9574
rect 21362 9208 21418 9217
rect 21362 9143 21364 9152
rect 21416 9143 21418 9152
rect 21364 9114 21416 9120
rect 21100 9030 21220 9058
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 20994 4176 21050 4185
rect 20994 4111 21050 4120
rect 21100 3738 21128 9030
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21192 7954 21220 8910
rect 21376 8634 21404 9114
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21192 7410 21220 7890
rect 21270 7576 21326 7585
rect 21270 7511 21326 7520
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21284 7342 21312 7511
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21180 3936 21232 3942
rect 21178 3904 21180 3913
rect 21232 3904 21234 3913
rect 21178 3839 21234 3848
rect 20904 3732 20956 3738
rect 21088 3732 21140 3738
rect 20904 3674 20956 3680
rect 21008 3692 21088 3720
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20640 3318 20760 3346
rect 20732 2689 20760 3318
rect 20824 3074 20852 3606
rect 21008 3194 21036 3692
rect 21088 3674 21140 3680
rect 21180 3664 21232 3670
rect 21100 3612 21180 3618
rect 21100 3606 21232 3612
rect 21100 3590 21220 3606
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20824 3046 20944 3074
rect 20916 2990 20944 3046
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20718 2680 20774 2689
rect 20824 2650 20852 2790
rect 20718 2615 20774 2624
rect 20812 2644 20864 2650
rect 20732 2582 20760 2615
rect 20812 2586 20864 2592
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 21100 1873 21128 3590
rect 21284 3369 21312 5510
rect 21376 3670 21404 7142
rect 21560 4554 21588 14418
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21638 13424 21694 13433
rect 21638 13359 21694 13368
rect 21652 4758 21680 13359
rect 21744 11898 21772 14214
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21836 11778 21864 15263
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22008 12300 22060 12306
rect 21928 12260 22008 12288
rect 21928 12102 21956 12260
rect 22008 12242 22060 12248
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21744 11750 21864 11778
rect 21744 5778 21772 11750
rect 21822 11656 21878 11665
rect 21822 11591 21878 11600
rect 21836 11558 21864 11591
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21928 11082 21956 12038
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21928 10742 21956 11018
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 22020 10554 22048 11834
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21928 10526 22048 10554
rect 21836 10130 21864 10474
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21744 5370 21772 5714
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21836 5166 21864 6054
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21652 4282 21680 4694
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21822 3768 21878 3777
rect 21928 3738 21956 10526
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 22020 10062 22048 10406
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 22020 8401 22048 8502
rect 22006 8392 22062 8401
rect 22006 8327 22062 8336
rect 22112 7426 22140 13942
rect 22296 13433 22324 15438
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22282 13424 22338 13433
rect 22282 13359 22338 13368
rect 22284 12368 22336 12374
rect 22284 12310 22336 12316
rect 22296 11898 22324 12310
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22284 11552 22336 11558
rect 22282 11520 22284 11529
rect 22336 11520 22338 11529
rect 22282 11455 22338 11464
rect 22388 11132 22416 14214
rect 22572 14074 22600 14418
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22296 11104 22416 11132
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22204 9081 22232 10542
rect 22296 10418 22324 11104
rect 22480 10470 22508 13670
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22572 11354 22600 13262
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22468 10464 22520 10470
rect 22296 10390 22416 10418
rect 22468 10406 22520 10412
rect 22388 10282 22416 10390
rect 22284 10260 22336 10266
rect 22388 10254 22508 10282
rect 22284 10202 22336 10208
rect 22296 9586 22324 10202
rect 22374 9888 22430 9897
rect 22374 9823 22430 9832
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22388 9178 22416 9823
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22190 9072 22246 9081
rect 22190 9007 22246 9016
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22296 8090 22324 8230
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22112 7398 22232 7426
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22112 7002 22140 7278
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22020 4826 22048 6054
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22112 4010 22140 4558
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 22204 3738 22232 7398
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22296 6254 22324 6394
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22296 5778 22324 6190
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22296 5030 22324 5714
rect 22480 5166 22508 10254
rect 22572 6202 22600 11154
rect 22664 10810 22692 17983
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 22756 11286 22784 14554
rect 22744 11280 22796 11286
rect 22744 11222 22796 11228
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22664 9194 22692 10406
rect 22756 10198 22784 11086
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22664 9166 22784 9194
rect 22848 9178 22876 18799
rect 23492 18057 23520 20023
rect 23478 18048 23534 18057
rect 23478 17983 23534 17992
rect 24044 17354 24072 26823
rect 24780 26314 24808 27503
rect 24768 26308 24820 26314
rect 24768 26250 24820 26256
rect 24122 26208 24178 26217
rect 24122 26143 24178 26152
rect 23768 17326 24072 17354
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22664 8362 22692 8978
rect 22652 8356 22704 8362
rect 22652 8298 22704 8304
rect 22664 7449 22692 8298
rect 22756 7993 22784 9166
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22742 7984 22798 7993
rect 22742 7919 22798 7928
rect 22836 7744 22888 7750
rect 22834 7712 22836 7721
rect 22888 7712 22890 7721
rect 22834 7647 22890 7656
rect 22650 7440 22706 7449
rect 22650 7375 22706 7384
rect 22940 7342 22968 15030
rect 23032 10441 23060 15846
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23018 10432 23074 10441
rect 23018 10367 23074 10376
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23032 9722 23060 10066
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23032 9042 23060 9658
rect 23124 9586 23152 9998
rect 23216 9654 23244 14758
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23308 9738 23336 13806
rect 23400 11540 23428 17070
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23584 14822 23612 15506
rect 23768 15450 23796 17326
rect 24136 17218 24164 26143
rect 25134 25528 25190 25537
rect 25134 25463 25190 25472
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24766 24848 24822 24857
rect 24766 24783 24822 24792
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24214 23488 24270 23497
rect 24214 23423 24270 23432
rect 24228 22114 24256 23423
rect 24780 23322 24808 24783
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23122
rect 24766 22808 24822 22817
rect 24676 22772 24728 22778
rect 24766 22743 24822 22752
rect 24676 22714 24728 22720
rect 24780 22250 24808 22743
rect 24780 22222 24900 22250
rect 24228 22086 24808 22114
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21570 24716 21966
rect 24780 21962 24808 22086
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24872 21842 24900 22222
rect 24596 21542 24716 21570
rect 24780 21814 24900 21842
rect 24596 21350 24624 21542
rect 24584 21344 24636 21350
rect 24582 21312 24584 21321
rect 24636 21312 24638 21321
rect 24582 21247 24638 21256
rect 24780 21146 24808 21814
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24216 21004 24268 21010
rect 24216 20946 24268 20952
rect 24228 20262 24256 20946
rect 24674 20768 24730 20777
rect 24289 20700 24585 20720
rect 24674 20703 24730 20712
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24216 20256 24268 20262
rect 24216 20198 24268 20204
rect 24228 17241 24256 20198
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 18873 24716 20703
rect 24766 19408 24822 19417
rect 24766 19343 24822 19352
rect 24674 18864 24730 18873
rect 24674 18799 24730 18808
rect 24674 18728 24730 18737
rect 24674 18663 24730 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 17898 24716 18663
rect 24596 17870 24716 17898
rect 24780 17882 24808 19343
rect 24858 18048 24914 18057
rect 24858 17983 24914 17992
rect 24768 17876 24820 17882
rect 24596 17610 24624 17870
rect 24768 17818 24820 17824
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24044 17190 24164 17218
rect 24214 17232 24270 17241
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23860 16182 23888 16594
rect 23848 16176 23900 16182
rect 23846 16144 23848 16153
rect 23900 16144 23902 16153
rect 23846 16079 23902 16088
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23768 15422 23888 15450
rect 23756 15360 23808 15366
rect 23754 15328 23756 15337
rect 23808 15328 23810 15337
rect 23754 15263 23810 15272
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23478 13560 23534 13569
rect 23478 13495 23534 13504
rect 23492 13394 23520 13495
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23480 11552 23532 11558
rect 23400 11512 23480 11540
rect 23480 11494 23532 11500
rect 23584 11370 23612 14758
rect 23860 14226 23888 15422
rect 23952 14929 23980 15506
rect 23938 14920 23994 14929
rect 23938 14855 23994 14864
rect 23860 14198 23980 14226
rect 23846 14104 23902 14113
rect 23846 14039 23902 14048
rect 23860 13938 23888 14039
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23846 13288 23902 13297
rect 23846 13223 23902 13232
rect 23662 13016 23718 13025
rect 23662 12951 23718 12960
rect 23676 11529 23704 12951
rect 23662 11520 23718 11529
rect 23662 11455 23718 11464
rect 23584 11342 23796 11370
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23400 10266 23428 10950
rect 23492 10606 23520 11222
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23584 10198 23612 11154
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23676 10577 23704 10678
rect 23662 10568 23718 10577
rect 23768 10554 23796 11342
rect 23860 11218 23888 13223
rect 23952 12986 23980 14198
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 24044 12442 24072 17190
rect 24688 17218 24716 17682
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24780 17338 24808 17546
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24872 17218 24900 17983
rect 24214 17167 24270 17176
rect 24412 17190 24716 17218
rect 24780 17190 24900 17218
rect 24412 16998 24440 17190
rect 24674 17096 24730 17105
rect 24674 17031 24730 17040
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16794 24440 16934
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24214 16688 24270 16697
rect 24124 16652 24176 16658
rect 24214 16623 24270 16632
rect 24124 16594 24176 16600
rect 24136 16289 24164 16594
rect 24122 16280 24178 16289
rect 24122 16215 24124 16224
rect 24176 16215 24178 16224
rect 24124 16186 24176 16192
rect 24228 15994 24256 16623
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24136 15966 24256 15994
rect 24136 14618 24164 15966
rect 24688 15706 24716 17031
rect 24780 16794 24808 17190
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24674 15328 24730 15337
rect 24289 15260 24585 15280
rect 24674 15263 24730 15272
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24400 14952 24452 14958
rect 24398 14920 24400 14929
rect 24584 14952 24636 14958
rect 24452 14920 24454 14929
rect 24584 14894 24636 14900
rect 24398 14855 24454 14864
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 24136 13870 24164 14418
rect 24596 14385 24624 14894
rect 24688 14634 24716 15263
rect 24780 15162 24808 15943
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24688 14606 24808 14634
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24582 14376 24638 14385
rect 24582 14311 24638 14320
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23952 11626 23980 12038
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 24044 11626 24072 11834
rect 23940 11620 23992 11626
rect 23940 11562 23992 11568
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 23848 11212 23900 11218
rect 23848 11154 23900 11160
rect 23952 11150 23980 11562
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 23768 10526 23888 10554
rect 23662 10503 23718 10512
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23754 10432 23810 10441
rect 23572 10192 23624 10198
rect 23572 10134 23624 10140
rect 23308 9710 23612 9738
rect 23204 9648 23256 9654
rect 23204 9590 23256 9596
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23124 9178 23152 9522
rect 23112 9172 23164 9178
rect 23112 9114 23164 9120
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23492 7857 23520 8298
rect 23478 7848 23534 7857
rect 23478 7783 23534 7792
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23492 7426 23520 7686
rect 23584 7546 23612 9710
rect 23676 9518 23704 10406
rect 23754 10367 23810 10376
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23676 9178 23704 9454
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23662 8392 23718 8401
rect 23662 8327 23718 8336
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23492 7398 23612 7426
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 22940 7002 22968 7278
rect 22928 6996 22980 7002
rect 22928 6938 22980 6944
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22940 6322 22968 6598
rect 23124 6458 23152 7278
rect 23584 7206 23612 7398
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 22572 6174 22692 6202
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5846 22600 6054
rect 22560 5840 22612 5846
rect 22560 5782 22612 5788
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22296 4622 22324 4966
rect 22480 4826 22508 5102
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22374 4176 22430 4185
rect 22374 4111 22430 4120
rect 21822 3703 21878 3712
rect 21916 3732 21968 3738
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21364 3528 21416 3534
rect 21456 3528 21508 3534
rect 21364 3470 21416 3476
rect 21454 3496 21456 3505
rect 21508 3496 21510 3505
rect 21270 3360 21326 3369
rect 21270 3295 21326 3304
rect 21376 3097 21404 3470
rect 21510 3454 21588 3482
rect 21454 3431 21510 3440
rect 21560 3194 21588 3454
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21362 3088 21418 3097
rect 21362 3023 21418 3032
rect 21454 2680 21510 2689
rect 21454 2615 21510 2624
rect 21468 2582 21496 2615
rect 21456 2576 21508 2582
rect 21456 2518 21508 2524
rect 21086 1864 21142 1873
rect 21086 1799 21142 1808
rect 20168 604 20220 610
rect 20168 546 20220 552
rect 20628 604 20680 610
rect 20628 546 20680 552
rect 21272 604 21324 610
rect 21272 546 21324 552
rect 20640 480 20668 546
rect 21284 480 21312 546
rect 21836 480 21864 3703
rect 21916 3674 21968 3680
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22100 2984 22152 2990
rect 21928 2932 22100 2938
rect 21928 2926 22152 2932
rect 21928 2910 22140 2926
rect 21928 2650 21956 2910
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 22020 2689 22048 2790
rect 22006 2680 22062 2689
rect 21916 2644 21968 2650
rect 22006 2615 22062 2624
rect 21916 2586 21968 2592
rect 22388 480 22416 4111
rect 22664 4078 22692 6174
rect 22744 5772 22796 5778
rect 22744 5714 22796 5720
rect 22756 5098 22784 5714
rect 22744 5092 22796 5098
rect 22744 5034 22796 5040
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22652 4072 22704 4078
rect 22704 4020 22784 4026
rect 22652 4014 22784 4020
rect 22664 3998 22784 4014
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22664 3777 22692 3878
rect 22650 3768 22706 3777
rect 22756 3738 22784 3998
rect 22848 3942 22876 4422
rect 23216 4185 23244 4966
rect 23202 4176 23258 4185
rect 23202 4111 23258 4120
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22650 3703 22706 3712
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22650 3496 22706 3505
rect 22650 3431 22652 3440
rect 22704 3431 22706 3440
rect 22652 3402 22704 3408
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22572 2854 22600 3130
rect 23018 2952 23074 2961
rect 23018 2887 23074 2896
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22572 2650 22600 2790
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 23032 480 23060 2887
rect 23308 2836 23336 7142
rect 23584 6798 23612 7142
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23400 5574 23428 6258
rect 23584 6254 23612 6734
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23388 5568 23440 5574
rect 23388 5510 23440 5516
rect 23400 4690 23428 5510
rect 23492 5137 23520 5782
rect 23676 5273 23704 8327
rect 23768 7478 23796 10367
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 23768 7274 23796 7414
rect 23756 7268 23808 7274
rect 23756 7210 23808 7216
rect 23754 7032 23810 7041
rect 23754 6967 23810 6976
rect 23662 5264 23718 5273
rect 23662 5199 23718 5208
rect 23478 5128 23534 5137
rect 23478 5063 23534 5072
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23400 4282 23428 4626
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23662 3904 23718 3913
rect 23584 3534 23612 3878
rect 23662 3839 23718 3848
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23584 2990 23612 3470
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23308 2808 23612 2836
rect 23584 480 23612 2808
rect 23676 1057 23704 3839
rect 23768 2922 23796 6967
rect 23860 5642 23888 10526
rect 24030 9208 24086 9217
rect 24030 9143 24086 9152
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 23952 8090 23980 8230
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23952 7410 23980 8026
rect 24044 7585 24072 9143
rect 24030 7576 24086 7585
rect 24030 7511 24086 7520
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23860 4010 23888 4422
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23860 3670 23888 3946
rect 24136 3942 24164 13806
rect 24688 13734 24716 14418
rect 24780 14090 24808 14606
rect 24780 14062 24900 14090
rect 24768 14000 24820 14006
rect 24766 13968 24768 13977
rect 24820 13968 24822 13977
rect 24766 13903 24822 13912
rect 24872 13818 24900 14062
rect 24780 13790 24900 13818
rect 24400 13728 24452 13734
rect 24400 13670 24452 13676
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24412 13530 24440 13670
rect 24780 13530 24808 13790
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12918 24716 13330
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24676 12776 24728 12782
rect 24964 12764 24992 15846
rect 24676 12718 24728 12724
rect 24780 12736 24992 12764
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24228 11082 24256 12242
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11218 24624 11494
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24228 10305 24256 11018
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10606 24716 12718
rect 24676 10600 24728 10606
rect 24306 10568 24362 10577
rect 24676 10542 24728 10548
rect 24306 10503 24362 10512
rect 24214 10296 24270 10305
rect 24214 10231 24270 10240
rect 24320 10010 24348 10503
rect 24228 9982 24348 10010
rect 24228 8498 24256 9982
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9586 24716 9862
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24596 8022 24624 8434
rect 24584 8016 24636 8022
rect 24584 7958 24636 7964
rect 24674 7848 24730 7857
rect 24674 7783 24730 7792
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24320 6934 24348 7346
rect 24308 6928 24360 6934
rect 24308 6870 24360 6876
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 5914 24716 7783
rect 24780 6882 24808 12736
rect 24858 12608 24914 12617
rect 24858 12543 24914 12552
rect 24872 11354 24900 12543
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 24858 11112 24914 11121
rect 24858 11047 24914 11056
rect 24872 7018 24900 11047
rect 24964 10810 24992 11154
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 25056 10674 25084 11494
rect 25148 11354 25176 25463
rect 25502 24168 25558 24177
rect 25502 24103 25558 24112
rect 25410 22128 25466 22137
rect 25410 22063 25466 22072
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25226 10704 25282 10713
rect 25044 10668 25096 10674
rect 25226 10639 25282 10648
rect 25044 10610 25096 10616
rect 25056 10266 25084 10610
rect 25240 10606 25268 10639
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 25226 10160 25282 10169
rect 25226 10095 25282 10104
rect 25240 9518 25268 10095
rect 25424 9654 25452 22063
rect 25516 10810 25544 24103
rect 25686 21448 25742 21457
rect 25686 21383 25742 21392
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 9110 24992 9318
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 24964 8634 24992 9046
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25148 8634 25176 8774
rect 25700 8634 25728 21383
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25148 7546 25176 8570
rect 25502 8528 25558 8537
rect 25502 8463 25558 8472
rect 25516 8430 25544 8463
rect 25504 8424 25556 8430
rect 25504 8366 25556 8372
rect 25226 7984 25282 7993
rect 25226 7919 25282 7928
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25240 7342 25268 7919
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 7410 25360 7686
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25228 7336 25280 7342
rect 25228 7278 25280 7284
rect 25412 7200 25464 7206
rect 25412 7142 25464 7148
rect 25424 7041 25452 7142
rect 25410 7032 25466 7041
rect 24872 6990 25084 7018
rect 24780 6854 24992 6882
rect 24858 6760 24914 6769
rect 24858 6695 24914 6704
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24214 5808 24270 5817
rect 24214 5743 24270 5752
rect 24228 4264 24256 5743
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5030 24716 5850
rect 24780 5234 24808 6190
rect 24872 5817 24900 6695
rect 24964 5914 24992 6854
rect 24952 5908 25004 5914
rect 24952 5850 25004 5856
rect 24858 5808 24914 5817
rect 24858 5743 24914 5752
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24872 5114 24900 5578
rect 24964 5302 24992 5850
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 24780 5098 24900 5114
rect 24780 5092 24912 5098
rect 24780 5086 24860 5092
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24780 4826 24808 5086
rect 24860 5034 24912 5040
rect 24872 5003 24900 5034
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 25056 4690 25084 6990
rect 25410 6967 25466 6976
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6254 25176 6598
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25504 6112 25556 6118
rect 25504 6054 25556 6060
rect 25516 5710 25544 6054
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 25504 5704 25556 5710
rect 25504 5646 25556 5652
rect 25148 5370 25176 5646
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24766 4448 24822 4457
rect 24289 4380 24585 4400
rect 24766 4383 24822 4392
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24228 4236 24348 4264
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 23940 3936 23992 3942
rect 23938 3904 23940 3913
rect 24124 3936 24176 3942
rect 23992 3904 23994 3913
rect 24124 3878 24176 3884
rect 23938 3839 23994 3848
rect 23848 3664 23900 3670
rect 23848 3606 23900 3612
rect 23860 3194 23888 3606
rect 24030 3360 24086 3369
rect 24030 3295 24086 3304
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23768 2310 23796 2450
rect 24044 2310 24072 3295
rect 24122 3224 24178 3233
rect 24122 3159 24178 3168
rect 24136 2961 24164 3159
rect 24122 2952 24178 2961
rect 24122 2887 24178 2896
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 23768 1873 23796 2246
rect 23754 1864 23810 1873
rect 23754 1799 23810 1808
rect 23662 1048 23718 1057
rect 23662 983 23718 992
rect 24136 480 24164 2790
rect 24228 2650 24256 3946
rect 24320 3913 24348 4236
rect 24584 4208 24636 4214
rect 24584 4150 24636 4156
rect 24596 4049 24624 4150
rect 24582 4040 24638 4049
rect 24582 3975 24638 3984
rect 24306 3904 24362 3913
rect 24306 3839 24362 3848
rect 24780 3641 24808 4383
rect 25056 4282 25084 4626
rect 27068 4480 27120 4486
rect 27068 4422 27120 4428
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 25318 4176 25374 4185
rect 25318 4111 25374 4120
rect 25504 4140 25556 4146
rect 24766 3632 24822 3641
rect 24766 3567 24822 3576
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24674 3224 24730 3233
rect 24674 3159 24730 3168
rect 24688 2825 24716 3159
rect 24780 2990 24808 3334
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 24674 2816 24730 2825
rect 24674 2751 24730 2760
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24780 2446 24808 2926
rect 24676 2440 24728 2446
rect 24674 2408 24676 2417
rect 24768 2440 24820 2446
rect 24728 2408 24730 2417
rect 24768 2382 24820 2388
rect 24674 2343 24730 2352
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24780 480 24808 2246
rect 25332 480 25360 4111
rect 25504 4082 25556 4088
rect 25516 3194 25544 4082
rect 25870 3768 25926 3777
rect 25870 3703 25926 3712
rect 25504 3188 25556 3194
rect 25504 3130 25556 3136
rect 25884 480 25912 3703
rect 26514 3496 26570 3505
rect 26514 3431 26570 3440
rect 26056 3120 26108 3126
rect 26054 3088 26056 3097
rect 26108 3088 26110 3097
rect 26054 3023 26110 3032
rect 26528 480 26556 3431
rect 27080 480 27108 4422
rect 27618 2816 27674 2825
rect 27618 2751 27674 2760
rect 27632 480 27660 2751
rect 18970 368 19026 377
rect 18970 303 19026 312
rect 19522 0 19578 480
rect 20074 0 20130 480
rect 20626 0 20682 480
rect 21270 0 21326 480
rect 21822 0 21878 480
rect 22374 0 22430 480
rect 23018 0 23074 480
rect 23570 0 23626 480
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25870 0 25926 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 1858 27512 1914 27568
rect 1582 24792 1638 24848
rect 1582 22072 1638 22128
rect 1490 21392 1546 21448
rect 1398 20712 1454 20768
rect 1582 20032 1638 20088
rect 1490 18672 1546 18728
rect 1398 17312 1454 17368
rect 1766 19352 1822 19408
rect 2962 26832 3018 26888
rect 2226 26152 2282 26208
rect 1950 25472 2006 25528
rect 1674 18708 1676 18728
rect 1676 18708 1728 18728
rect 1728 18708 1730 18728
rect 1674 18672 1730 18708
rect 1582 17992 1638 18048
rect 1582 15952 1638 16008
rect 1582 13912 1638 13968
rect 1674 13776 1730 13832
rect 2134 23432 2190 23488
rect 2042 18028 2044 18048
rect 2044 18028 2096 18048
rect 2096 18028 2098 18048
rect 2042 17992 2098 18028
rect 2042 16940 2044 16960
rect 2044 16940 2096 16960
rect 2096 16940 2098 16960
rect 2042 16904 2098 16940
rect 2042 16632 2098 16688
rect 2042 13640 2098 13696
rect 1858 12824 1914 12880
rect 1490 10920 1546 10976
rect 1950 9832 2006 9888
rect 2778 24112 2834 24168
rect 2410 17040 2466 17096
rect 2410 14476 2466 14512
rect 2410 14456 2412 14476
rect 2412 14456 2464 14476
rect 2464 14456 2466 14476
rect 2594 17720 2650 17776
rect 3882 22752 3938 22808
rect 3054 19896 3110 19952
rect 2594 15272 2650 15328
rect 2686 14592 2742 14648
rect 3054 13504 3110 13560
rect 2318 11756 2374 11792
rect 2318 11736 2320 11756
rect 2320 11736 2372 11756
rect 2372 11736 2374 11756
rect 1674 7520 1730 7576
rect 1582 6724 1638 6760
rect 1582 6704 1584 6724
rect 1584 6704 1636 6724
rect 1636 6704 1638 6724
rect 1490 6024 1546 6080
rect 1490 5072 1546 5128
rect 1398 3440 1454 3496
rect 846 2760 902 2816
rect 2042 8336 2098 8392
rect 1950 7248 2006 7304
rect 1950 4820 2006 4856
rect 1950 4800 1952 4820
rect 1952 4800 2004 4820
rect 2004 4800 2006 4820
rect 2134 4936 2190 4992
rect 2042 3848 2098 3904
rect 1858 3168 1914 3224
rect 1398 1672 1454 1728
rect 2594 10104 2650 10160
rect 2778 10260 2834 10296
rect 2778 10240 2780 10260
rect 2780 10240 2832 10260
rect 2832 10240 2834 10260
rect 2870 10004 2872 10024
rect 2872 10004 2924 10024
rect 2924 10004 2926 10024
rect 2870 9968 2926 10004
rect 3238 13932 3294 13968
rect 3238 13912 3240 13932
rect 3240 13912 3292 13932
rect 3292 13912 3294 13932
rect 3606 14320 3662 14376
rect 3330 12316 3332 12336
rect 3332 12316 3384 12336
rect 3384 12316 3386 12336
rect 3330 12280 3386 12316
rect 3422 12144 3478 12200
rect 3054 9152 3110 9208
rect 2870 9036 2926 9072
rect 2870 9016 2872 9036
rect 2872 9016 2924 9036
rect 2924 9016 2926 9036
rect 2594 7948 2650 7984
rect 2594 7928 2596 7948
rect 2596 7928 2648 7948
rect 2648 7928 2650 7948
rect 2686 6976 2742 7032
rect 2870 6840 2926 6896
rect 3238 10784 3294 10840
rect 3514 11872 3570 11928
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 13266 22616 13322 22672
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 12346 19896 12402 19952
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 11518 18672 11574 18728
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 7194 17992 7250 18048
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 4802 16904 4858 16960
rect 4710 13776 4766 13832
rect 4618 13640 4674 13696
rect 3514 9696 3570 9752
rect 3606 8200 3662 8256
rect 3698 7656 3754 7712
rect 3698 7384 3754 7440
rect 3606 6432 3662 6488
rect 2686 6024 2742 6080
rect 2594 5072 2650 5128
rect 2502 4800 2558 4856
rect 4066 8064 4122 8120
rect 4158 7404 4214 7440
rect 4158 7384 4160 7404
rect 4160 7384 4212 7404
rect 4212 7384 4214 7404
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 6366 15136 6422 15192
rect 4986 15000 5042 15056
rect 4802 11192 4858 11248
rect 4894 10804 4950 10840
rect 4894 10784 4896 10804
rect 4896 10784 4948 10804
rect 4948 10784 4950 10804
rect 4434 7792 4490 7848
rect 3974 5752 4030 5808
rect 3974 5636 4030 5672
rect 3974 5616 3976 5636
rect 3976 5616 4028 5636
rect 4028 5616 4030 5636
rect 3790 4120 3846 4176
rect 3422 3984 3478 4040
rect 3606 3984 3662 4040
rect 2778 3712 2834 3768
rect 2778 3032 2834 3088
rect 2318 2644 2374 2680
rect 2318 2624 2320 2644
rect 2320 2624 2372 2644
rect 2372 2624 2374 2644
rect 3146 3032 3202 3088
rect 2594 1944 2650 2000
rect 2226 992 2282 1048
rect 3790 3168 3846 3224
rect 3790 2896 3846 2952
rect 3606 2352 3662 2408
rect 4894 7112 4950 7168
rect 4618 2508 4674 2544
rect 4618 2488 4620 2508
rect 4620 2488 4672 2508
rect 4672 2488 4674 2508
rect 4526 2352 4582 2408
rect 4066 1264 4122 1320
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5078 12724 5080 12744
rect 5080 12724 5132 12744
rect 5132 12724 5134 12744
rect 5078 12688 5134 12724
rect 5998 12280 6054 12336
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5078 10956 5080 10976
rect 5080 10956 5132 10976
rect 5132 10956 5134 10976
rect 5078 10920 5134 10956
rect 5354 10532 5410 10568
rect 5354 10512 5356 10532
rect 5356 10512 5408 10532
rect 5408 10512 5410 10532
rect 5354 9832 5410 9888
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5998 9832 6054 9888
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5538 8064 5594 8120
rect 5814 8084 5870 8120
rect 5814 8064 5816 8084
rect 5816 8064 5868 8084
rect 5868 8064 5870 8084
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5630 6160 5686 6216
rect 5170 5616 5226 5672
rect 4986 1808 5042 1864
rect 5998 5480 6054 5536
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5814 5072 5870 5128
rect 5538 4800 5594 4856
rect 5814 4800 5870 4856
rect 5354 4428 5356 4448
rect 5356 4428 5408 4448
rect 5408 4428 5410 4448
rect 5354 4392 5410 4428
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5538 4120 5594 4176
rect 6734 14728 6790 14784
rect 6826 12416 6882 12472
rect 6182 11500 6184 11520
rect 6184 11500 6236 11520
rect 6236 11500 6238 11520
rect 6182 11464 6238 11500
rect 6274 10784 6330 10840
rect 6366 6976 6422 7032
rect 6274 5616 6330 5672
rect 6366 5072 6422 5128
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6642 6296 6698 6352
rect 6734 5072 6790 5128
rect 6642 4684 6698 4720
rect 6642 4664 6644 4684
rect 6644 4664 6696 4684
rect 6696 4664 6698 4684
rect 7102 13912 7158 13968
rect 7286 16632 7342 16688
rect 7194 10920 7250 10976
rect 7194 9968 7250 10024
rect 7102 7112 7158 7168
rect 6366 3848 6422 3904
rect 6274 2896 6330 2952
rect 5998 2624 6054 2680
rect 6550 2796 6552 2816
rect 6552 2796 6604 2816
rect 6604 2796 6606 2816
rect 6550 2760 6606 2796
rect 9678 17720 9734 17776
rect 8114 12552 8170 12608
rect 7562 12280 7618 12336
rect 7838 12144 7894 12200
rect 7562 11736 7618 11792
rect 7470 11328 7526 11384
rect 7378 10260 7434 10296
rect 7378 10240 7380 10260
rect 7380 10240 7432 10260
rect 7432 10240 7434 10260
rect 9402 16088 9458 16144
rect 9310 15952 9366 16008
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10598 17060 10654 17096
rect 10598 17040 10600 17060
rect 10600 17040 10652 17060
rect 10652 17040 10654 17060
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 9586 15544 9642 15600
rect 8574 15136 8630 15192
rect 8850 14864 8906 14920
rect 8850 14456 8906 14512
rect 8758 12960 8814 13016
rect 8298 11872 8354 11928
rect 7838 11192 7894 11248
rect 7562 10240 7618 10296
rect 7194 3188 7250 3224
rect 7194 3168 7196 3188
rect 7196 3168 7248 3188
rect 7248 3168 7250 3188
rect 7102 3032 7158 3088
rect 7286 3052 7342 3088
rect 7286 3032 7288 3052
rect 7288 3032 7340 3052
rect 7340 3032 7342 3052
rect 7470 9560 7526 9616
rect 7470 8472 7526 8528
rect 7654 7520 7710 7576
rect 8390 11228 8392 11248
rect 8392 11228 8444 11248
rect 8444 11228 8446 11248
rect 8390 11192 8446 11228
rect 8390 10920 8446 10976
rect 7930 8608 7986 8664
rect 8298 8780 8300 8800
rect 8300 8780 8352 8800
rect 8352 8780 8354 8800
rect 8298 8744 8354 8780
rect 8482 8472 8538 8528
rect 7470 4936 7526 4992
rect 7654 3712 7710 3768
rect 8022 7248 8078 7304
rect 7930 4120 7986 4176
rect 7930 3712 7986 3768
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6366 1944 6422 2000
rect 7562 1808 7618 1864
rect 7378 1672 7434 1728
rect 8390 5480 8446 5536
rect 8298 4936 8354 4992
rect 8298 4120 8354 4176
rect 8114 2760 8170 2816
rect 9402 13912 9458 13968
rect 9310 12416 9366 12472
rect 9310 10512 9366 10568
rect 8942 9988 8998 10024
rect 8942 9968 8944 9988
rect 8944 9968 8996 9988
rect 8996 9968 8998 9988
rect 9034 9460 9036 9480
rect 9036 9460 9088 9480
rect 9088 9460 9090 9480
rect 9034 9424 9090 9460
rect 9310 7420 9312 7440
rect 9312 7420 9364 7440
rect 9364 7420 9366 7440
rect 9310 7384 9366 7420
rect 8942 6160 8998 6216
rect 10046 14728 10102 14784
rect 9770 13776 9826 13832
rect 9586 12008 9642 12064
rect 9678 11892 9734 11928
rect 9678 11872 9680 11892
rect 9680 11872 9732 11892
rect 9732 11872 9734 11892
rect 9678 10240 9734 10296
rect 9678 7928 9734 7984
rect 9678 4664 9734 4720
rect 9586 3596 9642 3632
rect 9586 3576 9588 3596
rect 9588 3576 9640 3596
rect 9640 3576 9642 3596
rect 9034 2896 9090 2952
rect 9954 13504 10010 13560
rect 9954 12588 9956 12608
rect 9956 12588 10008 12608
rect 10008 12588 10010 12608
rect 9954 12552 10010 12588
rect 9862 11872 9918 11928
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10782 16632 10838 16688
rect 11242 16904 11298 16960
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 11058 15952 11114 16008
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10782 13232 10838 13288
rect 10782 12860 10784 12880
rect 10784 12860 10836 12880
rect 10836 12860 10838 12880
rect 10782 12824 10838 12860
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10690 12416 10746 12472
rect 10138 11872 10194 11928
rect 10046 11600 10102 11656
rect 9862 11464 9918 11520
rect 10046 11328 10102 11384
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10782 12008 10838 12064
rect 10046 10920 10102 10976
rect 10138 10784 10194 10840
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10874 10240 10930 10296
rect 11150 10104 11206 10160
rect 10874 9696 10930 9752
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10782 9324 10784 9344
rect 10784 9324 10836 9344
rect 10836 9324 10838 9344
rect 10782 9288 10838 9324
rect 9954 8472 10010 8528
rect 10046 8336 10102 8392
rect 9862 8200 9918 8256
rect 9954 3884 9956 3904
rect 9956 3884 10008 3904
rect 10008 3884 10010 3904
rect 9954 3848 10010 3884
rect 9862 3712 9918 3768
rect 10690 8200 10746 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10138 7964 10140 7984
rect 10140 7964 10192 7984
rect 10192 7964 10194 7984
rect 10138 7928 10194 7964
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10690 6840 10746 6896
rect 10506 6332 10508 6352
rect 10508 6332 10560 6352
rect 10560 6332 10562 6352
rect 10506 6296 10562 6332
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10138 5480 10194 5536
rect 10322 5208 10378 5264
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11150 9988 11206 10024
rect 11150 9968 11152 9988
rect 11152 9968 11204 9988
rect 11204 9968 11206 9988
rect 11518 12164 11574 12200
rect 11518 12144 11520 12164
rect 11520 12144 11572 12164
rect 11572 12144 11574 12164
rect 11702 11328 11758 11384
rect 11242 8336 11298 8392
rect 11242 8064 11298 8120
rect 11058 6860 11114 6896
rect 11058 6840 11060 6860
rect 11060 6840 11112 6860
rect 11112 6840 11114 6860
rect 10782 5344 10838 5400
rect 10782 4800 10838 4856
rect 10690 3984 10746 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10782 3848 10838 3904
rect 10690 3712 10746 3768
rect 11794 9832 11850 9888
rect 11702 9016 11758 9072
rect 11334 6160 11390 6216
rect 11334 5480 11390 5536
rect 10138 3440 10194 3496
rect 11334 4528 11390 4584
rect 11058 3984 11114 4040
rect 10966 3440 11022 3496
rect 10874 3304 10930 3360
rect 9954 3168 10010 3224
rect 11058 3032 11114 3088
rect 9034 2488 9090 2544
rect 8758 1944 8814 2000
rect 8574 1400 8630 1456
rect 9126 2372 9182 2408
rect 9126 2352 9128 2372
rect 9128 2352 9180 2372
rect 9180 2352 9182 2372
rect 10046 2216 10102 2272
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10230 2488 10286 2544
rect 10782 2624 10838 2680
rect 11334 3052 11390 3088
rect 11334 3032 11336 3052
rect 11336 3032 11388 3052
rect 11388 3032 11390 3052
rect 11794 7520 11850 7576
rect 11518 5072 11574 5128
rect 11702 5652 11704 5672
rect 11704 5652 11756 5672
rect 11756 5652 11758 5672
rect 11702 5616 11758 5652
rect 11610 1536 11666 1592
rect 13174 16088 13230 16144
rect 12898 15952 12954 16008
rect 12162 13368 12218 13424
rect 12254 12588 12256 12608
rect 12256 12588 12308 12608
rect 12308 12588 12310 12608
rect 12254 12552 12310 12588
rect 12714 12280 12770 12336
rect 12254 10512 12310 10568
rect 12162 10376 12218 10432
rect 11978 8472 12034 8528
rect 12162 7792 12218 7848
rect 12070 7384 12126 7440
rect 12530 9560 12586 9616
rect 12530 9288 12586 9344
rect 12438 8880 12494 8936
rect 12438 8472 12494 8528
rect 12162 4256 12218 4312
rect 12806 11872 12862 11928
rect 12806 11464 12862 11520
rect 12806 11192 12862 11248
rect 12622 5072 12678 5128
rect 12438 3848 12494 3904
rect 12254 3576 12310 3632
rect 12162 3304 12218 3360
rect 12898 9560 12954 9616
rect 12806 6976 12862 7032
rect 13174 11736 13230 11792
rect 13174 11464 13230 11520
rect 13174 10260 13230 10296
rect 13174 10240 13176 10260
rect 13176 10240 13228 10260
rect 13228 10240 13230 10260
rect 12990 8064 13046 8120
rect 13358 16088 13414 16144
rect 13358 15544 13414 15600
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 24766 27512 24822 27568
rect 24030 26832 24086 26888
rect 23662 22616 23718 22672
rect 23478 20032 23534 20088
rect 14830 19216 14886 19272
rect 23202 19216 23258 19272
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 22834 18808 22890 18864
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 22650 17992 22706 18048
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15658 17176 15714 17232
rect 13634 15428 13690 15464
rect 13634 15408 13636 15428
rect 13636 15408 13688 15428
rect 13688 15408 13690 15428
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 13634 14456 13690 14512
rect 14370 13776 14426 13832
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14738 13640 14794 13696
rect 14646 13404 14648 13424
rect 14648 13404 14700 13424
rect 14700 13404 14702 13424
rect 14646 13368 14702 13404
rect 13726 12960 13782 13016
rect 13542 12416 13598 12472
rect 13358 9424 13414 9480
rect 13450 8744 13506 8800
rect 12990 6840 13046 6896
rect 12898 5752 12954 5808
rect 12162 2932 12164 2952
rect 12164 2932 12216 2952
rect 12216 2932 12218 2952
rect 12162 2896 12218 2932
rect 12898 4392 12954 4448
rect 13358 6452 13414 6488
rect 13358 6432 13360 6452
rect 13360 6432 13412 6452
rect 13412 6432 13414 6452
rect 14002 11872 14058 11928
rect 13726 8880 13782 8936
rect 13726 8200 13782 8256
rect 13910 8336 13966 8392
rect 13726 6060 13728 6080
rect 13728 6060 13780 6080
rect 13780 6060 13782 6080
rect 13726 6024 13782 6060
rect 13634 5480 13690 5536
rect 13542 5364 13598 5400
rect 13542 5344 13544 5364
rect 13544 5344 13596 5364
rect 13596 5344 13598 5364
rect 14646 13096 14702 13152
rect 14646 12688 14702 12744
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15474 12824 15530 12880
rect 14738 12280 14794 12336
rect 14554 12008 14610 12064
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14278 9152 14334 9208
rect 13266 3848 13322 3904
rect 12898 3168 12954 3224
rect 13358 3732 13414 3768
rect 13358 3712 13360 3732
rect 13360 3712 13412 3732
rect 13412 3712 13414 3732
rect 14278 3576 14334 3632
rect 14278 3304 14334 3360
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14738 9832 14794 9888
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14830 9016 14886 9072
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14830 8336 14886 8392
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14830 6704 14886 6760
rect 15106 6704 15162 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15290 6160 15346 6216
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15014 4548 15070 4584
rect 15014 4528 15016 4548
rect 15016 4528 15068 4548
rect 15068 4528 15070 4548
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14646 3984 14702 4040
rect 14462 3712 14518 3768
rect 15290 3848 15346 3904
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15014 2624 15070 2680
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14554 1264 14610 1320
rect 17682 16904 17738 16960
rect 16210 16224 16266 16280
rect 15750 15544 15806 15600
rect 15658 15408 15714 15464
rect 15842 15000 15898 15056
rect 16118 13948 16120 13968
rect 16120 13948 16172 13968
rect 16172 13948 16174 13968
rect 15658 12552 15714 12608
rect 16118 13912 16174 13948
rect 17130 15952 17186 16008
rect 16302 14900 16304 14920
rect 16304 14900 16356 14920
rect 16356 14900 16358 14920
rect 16302 14864 16358 14900
rect 16486 14864 16542 14920
rect 16302 13948 16304 13968
rect 16304 13948 16356 13968
rect 16356 13948 16358 13968
rect 16302 13912 16358 13948
rect 16026 12688 16082 12744
rect 16118 12552 16174 12608
rect 16762 14456 16818 14512
rect 16854 14340 16910 14376
rect 16854 14320 16856 14340
rect 16856 14320 16908 14340
rect 16908 14320 16910 14340
rect 17038 14048 17094 14104
rect 16670 13776 16726 13832
rect 16762 13096 16818 13152
rect 16854 12688 16910 12744
rect 16394 12280 16450 12336
rect 16394 10648 16450 10704
rect 16854 10956 16856 10976
rect 16856 10956 16908 10976
rect 16908 10956 16910 10976
rect 16854 10920 16910 10956
rect 16670 9696 16726 9752
rect 15934 9288 15990 9344
rect 15934 8608 15990 8664
rect 15566 7112 15622 7168
rect 15474 3984 15530 4040
rect 15566 3732 15622 3768
rect 15566 3712 15568 3732
rect 15568 3712 15620 3732
rect 15620 3712 15622 3732
rect 15934 6840 15990 6896
rect 16854 7792 16910 7848
rect 16026 3848 16082 3904
rect 16210 2352 16266 2408
rect 16670 7384 16726 7440
rect 16670 6432 16726 6488
rect 16486 5244 16488 5264
rect 16488 5244 16540 5264
rect 16540 5244 16542 5264
rect 16486 5208 16542 5244
rect 17314 14356 17316 14376
rect 17316 14356 17368 14376
rect 17368 14356 17370 14376
rect 17314 14320 17370 14356
rect 17314 12960 17370 13016
rect 17222 9424 17278 9480
rect 17222 8472 17278 8528
rect 17314 7928 17370 7984
rect 17130 3984 17186 4040
rect 16854 3596 16910 3632
rect 16854 3576 16856 3596
rect 16856 3576 16908 3596
rect 16908 3576 16910 3596
rect 17038 3168 17094 3224
rect 16854 2644 16910 2680
rect 16854 2624 16856 2644
rect 16856 2624 16908 2644
rect 16908 2624 16910 2644
rect 16302 1672 16358 1728
rect 16578 1536 16634 1592
rect 17590 10648 17646 10704
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 18050 15988 18052 16008
rect 18052 15988 18104 16008
rect 18104 15988 18106 16008
rect 18050 15952 18106 15988
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 20810 15544 20866 15600
rect 18602 14456 18658 14512
rect 18510 12844 18566 12880
rect 18510 12824 18512 12844
rect 18512 12824 18564 12844
rect 18564 12824 18566 12844
rect 18510 12552 18566 12608
rect 18326 11056 18382 11112
rect 18602 11736 18658 11792
rect 18418 7520 18474 7576
rect 17958 7148 17960 7168
rect 17960 7148 18012 7168
rect 18012 7148 18014 7168
rect 17958 7112 18014 7148
rect 19062 12300 19118 12336
rect 19062 12280 19064 12300
rect 19064 12280 19116 12300
rect 19116 12280 19118 12300
rect 18970 11464 19026 11520
rect 19062 8880 19118 8936
rect 19062 8472 19118 8528
rect 17682 6840 17738 6896
rect 17498 6296 17554 6352
rect 17222 3576 17278 3632
rect 18142 3460 18198 3496
rect 18142 3440 18144 3460
rect 18144 3440 18196 3460
rect 18196 3440 18198 3460
rect 18326 3304 18382 3360
rect 17774 1944 17830 2000
rect 18878 6996 18934 7032
rect 18878 6976 18880 6996
rect 18880 6976 18932 6996
rect 18932 6976 18934 6996
rect 18970 6024 19026 6080
rect 19062 5616 19118 5672
rect 19246 11328 19302 11384
rect 19246 8356 19302 8392
rect 19246 8336 19248 8356
rect 19248 8336 19300 8356
rect 19300 8336 19302 8356
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19614 13912 19670 13968
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19522 12708 19578 12744
rect 19522 12688 19524 12708
rect 19524 12688 19576 12708
rect 19576 12688 19578 12708
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19982 11736 20038 11792
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19706 11212 19762 11248
rect 19706 11192 19708 11212
rect 19708 11192 19760 11212
rect 19760 11192 19762 11212
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19798 9968 19854 10024
rect 19982 9988 20038 10024
rect 19982 9968 19984 9988
rect 19984 9968 20036 9988
rect 20036 9968 20038 9988
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20442 13232 20498 13288
rect 21822 15272 21878 15328
rect 20810 13504 20866 13560
rect 20350 11056 20406 11112
rect 20534 11056 20590 11112
rect 20810 9560 20866 9616
rect 20718 9460 20720 9480
rect 20720 9460 20772 9480
rect 20772 9460 20774 9480
rect 20718 9424 20774 9460
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19614 7520 19670 7576
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19338 6296 19394 6352
rect 19338 6196 19340 6216
rect 19340 6196 19392 6216
rect 19392 6196 19394 6216
rect 19338 6160 19394 6196
rect 4066 312 4122 368
rect 20442 8608 20498 8664
rect 20166 7284 20168 7304
rect 20168 7284 20220 7304
rect 20220 7284 20222 7304
rect 20166 7248 20222 7284
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19614 5616 19670 5672
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19430 4800 19486 4856
rect 19430 3884 19432 3904
rect 19432 3884 19484 3904
rect 19484 3884 19486 3904
rect 19430 3848 19486 3884
rect 20074 5072 20130 5128
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19522 3032 19578 3088
rect 19246 2896 19302 2952
rect 19430 2896 19486 2952
rect 19890 2896 19946 2952
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20258 4120 20314 4176
rect 20810 5208 20866 5264
rect 20350 3712 20406 3768
rect 20810 3984 20866 4040
rect 21086 11500 21088 11520
rect 21088 11500 21140 11520
rect 21140 11500 21142 11520
rect 21086 11464 21142 11500
rect 20994 10920 21050 10976
rect 21086 10104 21142 10160
rect 21362 9172 21418 9208
rect 21362 9152 21364 9172
rect 21364 9152 21416 9172
rect 21416 9152 21418 9172
rect 20994 4120 21050 4176
rect 21270 7520 21326 7576
rect 21178 3884 21180 3904
rect 21180 3884 21232 3904
rect 21232 3884 21234 3904
rect 21178 3848 21234 3884
rect 20718 2624 20774 2680
rect 21638 13368 21694 13424
rect 21822 11600 21878 11656
rect 21822 3712 21878 3768
rect 22006 8336 22062 8392
rect 22282 13368 22338 13424
rect 22282 11500 22284 11520
rect 22284 11500 22336 11520
rect 22336 11500 22338 11520
rect 22282 11464 22338 11500
rect 22374 9832 22430 9888
rect 22190 9016 22246 9072
rect 23478 17992 23534 18048
rect 24122 26152 24178 26208
rect 22742 7928 22798 7984
rect 22834 7692 22836 7712
rect 22836 7692 22888 7712
rect 22888 7692 22890 7712
rect 22834 7656 22890 7692
rect 22650 7384 22706 7440
rect 23018 10376 23074 10432
rect 25134 25472 25190 25528
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24792 24822 24848
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24214 23432 24270 23488
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22752 24822 22808
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24582 21292 24584 21312
rect 24584 21292 24636 21312
rect 24636 21292 24638 21312
rect 24582 21256 24638 21292
rect 24674 20712 24730 20768
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 19352 24822 19408
rect 24674 18808 24730 18864
rect 24674 18672 24730 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24858 17992 24914 18048
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 23846 16124 23848 16144
rect 23848 16124 23900 16144
rect 23900 16124 23902 16144
rect 23846 16088 23902 16124
rect 23754 15308 23756 15328
rect 23756 15308 23808 15328
rect 23808 15308 23810 15328
rect 23754 15272 23810 15308
rect 23478 13504 23534 13560
rect 23938 14864 23994 14920
rect 23846 14048 23902 14104
rect 23846 13232 23902 13288
rect 23662 12960 23718 13016
rect 23662 11464 23718 11520
rect 23662 10512 23718 10568
rect 24214 17176 24270 17232
rect 24674 17040 24730 17096
rect 24214 16632 24270 16688
rect 24122 16244 24178 16280
rect 24122 16224 24124 16244
rect 24124 16224 24176 16244
rect 24176 16224 24178 16244
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24766 15952 24822 16008
rect 24674 15272 24730 15328
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24398 14900 24400 14920
rect 24400 14900 24452 14920
rect 24452 14900 24454 14920
rect 24398 14864 24454 14900
rect 24582 14320 24638 14376
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 23478 7792 23534 7848
rect 23754 10376 23810 10432
rect 23662 8336 23718 8392
rect 22374 4120 22430 4176
rect 21454 3476 21456 3496
rect 21456 3476 21508 3496
rect 21508 3476 21510 3496
rect 21270 3304 21326 3360
rect 21454 3440 21510 3476
rect 21362 3032 21418 3088
rect 21454 2624 21510 2680
rect 21086 1808 21142 1864
rect 22006 2624 22062 2680
rect 22650 3712 22706 3768
rect 23202 4120 23258 4176
rect 22650 3460 22706 3496
rect 22650 3440 22652 3460
rect 22652 3440 22704 3460
rect 22704 3440 22706 3460
rect 23018 2896 23074 2952
rect 23754 6976 23810 7032
rect 23662 5208 23718 5264
rect 23478 5072 23534 5128
rect 23662 3848 23718 3904
rect 24030 9152 24086 9208
rect 24030 7520 24086 7576
rect 24766 13948 24768 13968
rect 24768 13948 24820 13968
rect 24820 13948 24822 13968
rect 24766 13912 24822 13948
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24306 10512 24362 10568
rect 24214 10240 24270 10296
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24674 7792 24730 7848
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24858 12552 24914 12608
rect 24858 11056 24914 11112
rect 25502 24112 25558 24168
rect 25410 22072 25466 22128
rect 25226 10648 25282 10704
rect 25226 10104 25282 10160
rect 25686 21392 25742 21448
rect 25502 8472 25558 8528
rect 25226 7928 25282 7984
rect 24858 6704 24914 6760
rect 24214 5752 24270 5808
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24858 5752 24914 5808
rect 25410 6976 25466 7032
rect 24766 4392 24822 4448
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23938 3884 23940 3904
rect 23940 3884 23992 3904
rect 23992 3884 23994 3904
rect 23938 3848 23994 3884
rect 24030 3304 24086 3360
rect 24122 3168 24178 3224
rect 24122 2896 24178 2952
rect 23754 1808 23810 1864
rect 23662 992 23718 1048
rect 24582 3984 24638 4040
rect 24306 3848 24362 3904
rect 25318 4120 25374 4176
rect 24766 3576 24822 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24674 3168 24730 3224
rect 24674 2760 24730 2816
rect 24674 2388 24676 2408
rect 24676 2388 24728 2408
rect 24728 2388 24730 2408
rect 24674 2352 24730 2388
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25870 3712 25926 3768
rect 26514 3440 26570 3496
rect 26054 3068 26056 3088
rect 26056 3068 26108 3088
rect 26108 3068 26110 3088
rect 26054 3032 26110 3068
rect 27618 2760 27674 2816
rect 18970 312 19026 368
<< metal3 >>
rect 0 27570 480 27600
rect 1853 27570 1919 27573
rect 0 27568 1919 27570
rect 0 27512 1858 27568
rect 1914 27512 1919 27568
rect 0 27510 1919 27512
rect 0 27480 480 27510
rect 1853 27507 1919 27510
rect 24761 27570 24827 27573
rect 27520 27570 28000 27600
rect 24761 27568 28000 27570
rect 24761 27512 24766 27568
rect 24822 27512 28000 27568
rect 24761 27510 28000 27512
rect 24761 27507 24827 27510
rect 27520 27480 28000 27510
rect 0 26890 480 26920
rect 2957 26890 3023 26893
rect 0 26888 3023 26890
rect 0 26832 2962 26888
rect 3018 26832 3023 26888
rect 0 26830 3023 26832
rect 0 26800 480 26830
rect 2957 26827 3023 26830
rect 24025 26890 24091 26893
rect 27520 26890 28000 26920
rect 24025 26888 28000 26890
rect 24025 26832 24030 26888
rect 24086 26832 28000 26888
rect 24025 26830 28000 26832
rect 24025 26827 24091 26830
rect 27520 26800 28000 26830
rect 0 26210 480 26240
rect 2221 26210 2287 26213
rect 0 26208 2287 26210
rect 0 26152 2226 26208
rect 2282 26152 2287 26208
rect 0 26150 2287 26152
rect 0 26120 480 26150
rect 2221 26147 2287 26150
rect 24117 26210 24183 26213
rect 27520 26210 28000 26240
rect 24117 26208 28000 26210
rect 24117 26152 24122 26208
rect 24178 26152 28000 26208
rect 24117 26150 28000 26152
rect 24117 26147 24183 26150
rect 27520 26120 28000 26150
rect 10277 25600 10597 25601
rect 0 25530 480 25560
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1945 25530 2011 25533
rect 0 25528 2011 25530
rect 0 25472 1950 25528
rect 2006 25472 2011 25528
rect 0 25470 2011 25472
rect 0 25440 480 25470
rect 1945 25467 2011 25470
rect 25129 25530 25195 25533
rect 27520 25530 28000 25560
rect 25129 25528 28000 25530
rect 25129 25472 25134 25528
rect 25190 25472 28000 25528
rect 25129 25470 28000 25472
rect 25129 25467 25195 25470
rect 27520 25440 28000 25470
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 1577 24850 1643 24853
rect 0 24848 1643 24850
rect 0 24792 1582 24848
rect 1638 24792 1643 24848
rect 0 24790 1643 24792
rect 0 24760 480 24790
rect 1577 24787 1643 24790
rect 24761 24850 24827 24853
rect 27520 24850 28000 24880
rect 24761 24848 28000 24850
rect 24761 24792 24766 24848
rect 24822 24792 28000 24848
rect 24761 24790 28000 24792
rect 24761 24787 24827 24790
rect 27520 24760 28000 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24170 480 24200
rect 2773 24170 2839 24173
rect 0 24168 2839 24170
rect 0 24112 2778 24168
rect 2834 24112 2839 24168
rect 0 24110 2839 24112
rect 0 24080 480 24110
rect 2773 24107 2839 24110
rect 25497 24170 25563 24173
rect 27520 24170 28000 24200
rect 25497 24168 28000 24170
rect 25497 24112 25502 24168
rect 25558 24112 28000 24168
rect 25497 24110 28000 24112
rect 25497 24107 25563 24110
rect 27520 24080 28000 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 0 23490 480 23520
rect 2129 23490 2195 23493
rect 0 23488 2195 23490
rect 0 23432 2134 23488
rect 2190 23432 2195 23488
rect 0 23430 2195 23432
rect 0 23400 480 23430
rect 2129 23427 2195 23430
rect 24209 23490 24275 23493
rect 27520 23490 28000 23520
rect 24209 23488 28000 23490
rect 24209 23432 24214 23488
rect 24270 23432 28000 23488
rect 24209 23430 28000 23432
rect 24209 23427 24275 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 27520 23400 28000 23430
rect 19610 23359 19930 23360
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 3877 22810 3943 22813
rect 0 22808 3943 22810
rect 0 22752 3882 22808
rect 3938 22752 3943 22808
rect 0 22750 3943 22752
rect 0 22720 480 22750
rect 3877 22747 3943 22750
rect 24761 22810 24827 22813
rect 27520 22810 28000 22840
rect 24761 22808 28000 22810
rect 24761 22752 24766 22808
rect 24822 22752 28000 22808
rect 24761 22750 28000 22752
rect 24761 22747 24827 22750
rect 27520 22720 28000 22750
rect 13261 22674 13327 22677
rect 23657 22674 23723 22677
rect 13261 22672 23723 22674
rect 13261 22616 13266 22672
rect 13322 22616 23662 22672
rect 23718 22616 23723 22672
rect 13261 22614 23723 22616
rect 13261 22611 13327 22614
rect 23657 22611 23723 22614
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 0 22130 480 22160
rect 1577 22130 1643 22133
rect 0 22128 1643 22130
rect 0 22072 1582 22128
rect 1638 22072 1643 22128
rect 0 22070 1643 22072
rect 0 22040 480 22070
rect 1577 22067 1643 22070
rect 25405 22130 25471 22133
rect 27520 22130 28000 22160
rect 25405 22128 28000 22130
rect 25405 22072 25410 22128
rect 25466 22072 28000 22128
rect 25405 22070 28000 22072
rect 25405 22067 25471 22070
rect 27520 22040 28000 22070
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21450 480 21480
rect 1485 21450 1551 21453
rect 0 21448 1551 21450
rect 0 21392 1490 21448
rect 1546 21392 1551 21448
rect 0 21390 1551 21392
rect 0 21360 480 21390
rect 1485 21387 1551 21390
rect 25681 21450 25747 21453
rect 27520 21450 28000 21480
rect 25681 21448 28000 21450
rect 25681 21392 25686 21448
rect 25742 21392 28000 21448
rect 25681 21390 28000 21392
rect 25681 21387 25747 21390
rect 27520 21360 28000 21390
rect 21214 21252 21220 21316
rect 21284 21314 21290 21316
rect 24577 21314 24643 21317
rect 21284 21312 24643 21314
rect 21284 21256 24582 21312
rect 24638 21256 24643 21312
rect 21284 21254 24643 21256
rect 21284 21252 21290 21254
rect 24577 21251 24643 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 20770 480 20800
rect 1393 20770 1459 20773
rect 0 20768 1459 20770
rect 0 20712 1398 20768
rect 1454 20712 1459 20768
rect 0 20710 1459 20712
rect 0 20680 480 20710
rect 1393 20707 1459 20710
rect 24669 20770 24735 20773
rect 27520 20770 28000 20800
rect 24669 20768 28000 20770
rect 24669 20712 24674 20768
rect 24730 20712 28000 20768
rect 24669 20710 28000 20712
rect 24669 20707 24735 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 480 20030
rect 1577 20027 1643 20030
rect 23473 20090 23539 20093
rect 27520 20090 28000 20120
rect 23473 20088 28000 20090
rect 23473 20032 23478 20088
rect 23534 20032 28000 20088
rect 23473 20030 28000 20032
rect 23473 20027 23539 20030
rect 27520 20000 28000 20030
rect 3049 19954 3115 19957
rect 12341 19954 12407 19957
rect 3049 19952 12407 19954
rect 3049 19896 3054 19952
rect 3110 19896 12346 19952
rect 12402 19896 12407 19952
rect 3049 19894 12407 19896
rect 3049 19891 3115 19894
rect 12341 19891 12407 19894
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19410 480 19440
rect 1761 19410 1827 19413
rect 0 19408 1827 19410
rect 0 19352 1766 19408
rect 1822 19352 1827 19408
rect 0 19350 1827 19352
rect 0 19320 480 19350
rect 1761 19347 1827 19350
rect 24761 19410 24827 19413
rect 27520 19410 28000 19440
rect 24761 19408 28000 19410
rect 24761 19352 24766 19408
rect 24822 19352 28000 19408
rect 24761 19350 28000 19352
rect 24761 19347 24827 19350
rect 27520 19320 28000 19350
rect 14825 19274 14891 19277
rect 23197 19274 23263 19277
rect 14825 19272 23263 19274
rect 14825 19216 14830 19272
rect 14886 19216 23202 19272
rect 23258 19216 23263 19272
rect 14825 19214 23263 19216
rect 14825 19211 14891 19214
rect 23197 19211 23263 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 22829 18866 22895 18869
rect 24669 18866 24735 18869
rect 22829 18864 24735 18866
rect 22829 18808 22834 18864
rect 22890 18808 24674 18864
rect 24730 18808 24735 18864
rect 22829 18806 24735 18808
rect 22829 18803 22895 18806
rect 24669 18803 24735 18806
rect 0 18730 480 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 480 18670
rect 1485 18667 1551 18670
rect 1669 18730 1735 18733
rect 11513 18730 11579 18733
rect 1669 18728 11579 18730
rect 1669 18672 1674 18728
rect 1730 18672 11518 18728
rect 11574 18672 11579 18728
rect 1669 18670 11579 18672
rect 1669 18667 1735 18670
rect 11513 18667 11579 18670
rect 24669 18730 24735 18733
rect 27520 18730 28000 18760
rect 24669 18728 28000 18730
rect 24669 18672 24674 18728
rect 24730 18672 28000 18728
rect 24669 18670 28000 18672
rect 24669 18667 24735 18670
rect 27520 18640 28000 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 0 18050 480 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 480 17990
rect 1577 17987 1643 17990
rect 2037 18050 2103 18053
rect 7189 18050 7255 18053
rect 2037 18048 7255 18050
rect 2037 17992 2042 18048
rect 2098 17992 7194 18048
rect 7250 17992 7255 18048
rect 2037 17990 7255 17992
rect 2037 17987 2103 17990
rect 7189 17987 7255 17990
rect 22645 18050 22711 18053
rect 23473 18050 23539 18053
rect 22645 18048 23539 18050
rect 22645 17992 22650 18048
rect 22706 17992 23478 18048
rect 23534 17992 23539 18048
rect 22645 17990 23539 17992
rect 22645 17987 22711 17990
rect 23473 17987 23539 17990
rect 24853 18050 24919 18053
rect 27520 18050 28000 18080
rect 24853 18048 28000 18050
rect 24853 17992 24858 18048
rect 24914 17992 28000 18048
rect 24853 17990 28000 17992
rect 24853 17987 24919 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 2589 17778 2655 17781
rect 9673 17778 9739 17781
rect 2589 17776 9739 17778
rect 2589 17720 2594 17776
rect 2650 17720 9678 17776
rect 9734 17720 9739 17776
rect 2589 17718 9739 17720
rect 2589 17715 2655 17718
rect 9673 17715 9739 17718
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 1393 17370 1459 17373
rect 27520 17370 28000 17400
rect 0 17368 1459 17370
rect 0 17312 1398 17368
rect 1454 17312 1459 17368
rect 0 17310 1459 17312
rect 0 17280 480 17310
rect 1393 17307 1459 17310
rect 24718 17310 28000 17370
rect 15653 17234 15719 17237
rect 24209 17234 24275 17237
rect 15653 17232 24275 17234
rect 15653 17176 15658 17232
rect 15714 17176 24214 17232
rect 24270 17176 24275 17232
rect 15653 17174 24275 17176
rect 15653 17171 15719 17174
rect 24209 17171 24275 17174
rect 24718 17101 24778 17310
rect 27520 17280 28000 17310
rect 2405 17098 2471 17101
rect 10593 17098 10659 17101
rect 2405 17096 10659 17098
rect 2405 17040 2410 17096
rect 2466 17040 10598 17096
rect 10654 17040 10659 17096
rect 2405 17038 10659 17040
rect 2405 17035 2471 17038
rect 10593 17035 10659 17038
rect 24669 17096 24778 17101
rect 24669 17040 24674 17096
rect 24730 17040 24778 17096
rect 24669 17038 24778 17040
rect 24669 17035 24735 17038
rect 2037 16962 2103 16965
rect 4797 16962 4863 16965
rect 2037 16960 4863 16962
rect 2037 16904 2042 16960
rect 2098 16904 4802 16960
rect 4858 16904 4863 16960
rect 2037 16902 4863 16904
rect 2037 16899 2103 16902
rect 4797 16899 4863 16902
rect 11237 16962 11303 16965
rect 17677 16962 17743 16965
rect 11237 16960 17743 16962
rect 11237 16904 11242 16960
rect 11298 16904 17682 16960
rect 17738 16904 17743 16960
rect 11237 16902 17743 16904
rect 11237 16899 11303 16902
rect 17677 16899 17743 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16690 480 16720
rect 2037 16690 2103 16693
rect 0 16688 2103 16690
rect 0 16632 2042 16688
rect 2098 16632 2103 16688
rect 0 16630 2103 16632
rect 0 16600 480 16630
rect 2037 16627 2103 16630
rect 7281 16690 7347 16693
rect 10777 16690 10843 16693
rect 7281 16688 10843 16690
rect 7281 16632 7286 16688
rect 7342 16632 10782 16688
rect 10838 16632 10843 16688
rect 7281 16630 10843 16632
rect 7281 16627 7347 16630
rect 10777 16627 10843 16630
rect 24209 16690 24275 16693
rect 27520 16690 28000 16720
rect 24209 16688 28000 16690
rect 24209 16632 24214 16688
rect 24270 16632 28000 16688
rect 24209 16630 28000 16632
rect 24209 16627 24275 16630
rect 27520 16600 28000 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 16205 16282 16271 16285
rect 24117 16282 24183 16285
rect 16205 16280 24183 16282
rect 16205 16224 16210 16280
rect 16266 16224 24122 16280
rect 24178 16224 24183 16280
rect 16205 16222 24183 16224
rect 16205 16219 16271 16222
rect 24117 16219 24183 16222
rect 9397 16146 9463 16149
rect 13169 16146 13235 16149
rect 13353 16146 13419 16149
rect 23841 16146 23907 16149
rect 9397 16144 13419 16146
rect 9397 16088 9402 16144
rect 9458 16088 13174 16144
rect 13230 16088 13358 16144
rect 13414 16088 13419 16144
rect 9397 16086 13419 16088
rect 9397 16083 9463 16086
rect 13169 16083 13235 16086
rect 13353 16083 13419 16086
rect 13494 16144 23907 16146
rect 13494 16088 23846 16144
rect 23902 16088 23907 16144
rect 13494 16086 23907 16088
rect 0 16010 480 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 480 15950
rect 1577 15947 1643 15950
rect 9305 16010 9371 16013
rect 11053 16010 11119 16013
rect 9305 16008 11119 16010
rect 9305 15952 9310 16008
rect 9366 15952 11058 16008
rect 11114 15952 11119 16008
rect 9305 15950 11119 15952
rect 9305 15947 9371 15950
rect 11053 15947 11119 15950
rect 12893 16010 12959 16013
rect 13494 16010 13554 16086
rect 23841 16083 23907 16086
rect 12893 16008 13554 16010
rect 12893 15952 12898 16008
rect 12954 15952 13554 16008
rect 12893 15950 13554 15952
rect 17125 16010 17191 16013
rect 18045 16010 18111 16013
rect 17125 16008 18111 16010
rect 17125 15952 17130 16008
rect 17186 15952 18050 16008
rect 18106 15952 18111 16008
rect 17125 15950 18111 15952
rect 12893 15947 12959 15950
rect 17125 15947 17191 15950
rect 18045 15947 18111 15950
rect 24761 16010 24827 16013
rect 27520 16010 28000 16040
rect 24761 16008 28000 16010
rect 24761 15952 24766 16008
rect 24822 15952 28000 16008
rect 24761 15950 28000 15952
rect 24761 15947 24827 15950
rect 27520 15920 28000 15950
rect 13126 15814 15946 15874
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 9581 15602 9647 15605
rect 13126 15602 13186 15814
rect 9581 15600 13186 15602
rect 9581 15544 9586 15600
rect 9642 15544 13186 15600
rect 9581 15542 13186 15544
rect 13353 15602 13419 15605
rect 15745 15602 15811 15605
rect 13353 15600 15811 15602
rect 13353 15544 13358 15600
rect 13414 15544 15750 15600
rect 15806 15544 15811 15600
rect 13353 15542 15811 15544
rect 15886 15602 15946 15814
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 20805 15602 20871 15605
rect 15886 15600 20871 15602
rect 15886 15544 20810 15600
rect 20866 15544 20871 15600
rect 15886 15542 20871 15544
rect 9581 15539 9647 15542
rect 13353 15539 13419 15542
rect 15745 15539 15811 15542
rect 20805 15539 20871 15542
rect 13629 15466 13695 15469
rect 15653 15466 15719 15469
rect 13629 15464 15719 15466
rect 13629 15408 13634 15464
rect 13690 15408 15658 15464
rect 15714 15408 15719 15464
rect 13629 15406 15719 15408
rect 13629 15403 13695 15406
rect 15653 15403 15719 15406
rect 0 15330 480 15360
rect 2589 15330 2655 15333
rect 0 15328 2655 15330
rect 0 15272 2594 15328
rect 2650 15272 2655 15328
rect 0 15270 2655 15272
rect 0 15240 480 15270
rect 2589 15267 2655 15270
rect 21817 15330 21883 15333
rect 23749 15330 23815 15333
rect 21817 15328 23815 15330
rect 21817 15272 21822 15328
rect 21878 15272 23754 15328
rect 23810 15272 23815 15328
rect 21817 15270 23815 15272
rect 21817 15267 21883 15270
rect 23749 15267 23815 15270
rect 24669 15330 24735 15333
rect 27520 15330 28000 15360
rect 24669 15328 28000 15330
rect 24669 15272 24674 15328
rect 24730 15272 28000 15328
rect 24669 15270 28000 15272
rect 24669 15267 24735 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 27520 15240 28000 15270
rect 24277 15199 24597 15200
rect 6361 15194 6427 15197
rect 8569 15194 8635 15197
rect 6361 15192 8635 15194
rect 6361 15136 6366 15192
rect 6422 15136 8574 15192
rect 8630 15136 8635 15192
rect 6361 15134 8635 15136
rect 6361 15131 6427 15134
rect 8569 15131 8635 15134
rect 4981 15058 5047 15061
rect 15837 15058 15903 15061
rect 4981 15056 15903 15058
rect 4981 15000 4986 15056
rect 5042 15000 15842 15056
rect 15898 15000 15903 15056
rect 4981 14998 15903 15000
rect 4981 14995 5047 14998
rect 15837 14995 15903 14998
rect 8845 14922 8911 14925
rect 16297 14922 16363 14925
rect 8845 14920 16363 14922
rect 8845 14864 8850 14920
rect 8906 14864 16302 14920
rect 16358 14864 16363 14920
rect 8845 14862 16363 14864
rect 8845 14859 8911 14862
rect 16297 14859 16363 14862
rect 16481 14922 16547 14925
rect 23933 14922 23999 14925
rect 24393 14922 24459 14925
rect 16481 14920 24459 14922
rect 16481 14864 16486 14920
rect 16542 14864 23938 14920
rect 23994 14864 24398 14920
rect 24454 14864 24459 14920
rect 16481 14862 24459 14864
rect 16481 14859 16547 14862
rect 23933 14859 23999 14862
rect 24393 14859 24459 14862
rect 6729 14786 6795 14789
rect 10041 14786 10107 14789
rect 6729 14784 10107 14786
rect 6729 14728 6734 14784
rect 6790 14728 10046 14784
rect 10102 14728 10107 14784
rect 6729 14726 10107 14728
rect 6729 14723 6795 14726
rect 10041 14723 10107 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 2681 14650 2747 14653
rect 27520 14650 28000 14680
rect 0 14648 2747 14650
rect 0 14592 2686 14648
rect 2742 14592 2747 14648
rect 0 14590 2747 14592
rect 0 14560 480 14590
rect 2681 14587 2747 14590
rect 27478 14560 28000 14650
rect 2405 14514 2471 14517
rect 8845 14514 8911 14517
rect 2405 14512 8911 14514
rect 2405 14456 2410 14512
rect 2466 14456 8850 14512
rect 8906 14456 8911 14512
rect 2405 14454 8911 14456
rect 2405 14451 2471 14454
rect 8845 14451 8911 14454
rect 13629 14514 13695 14517
rect 16757 14514 16823 14517
rect 13629 14512 16823 14514
rect 13629 14456 13634 14512
rect 13690 14456 16762 14512
rect 16818 14456 16823 14512
rect 13629 14454 16823 14456
rect 13629 14451 13695 14454
rect 16757 14451 16823 14454
rect 18597 14514 18663 14517
rect 27478 14514 27538 14560
rect 18597 14512 27538 14514
rect 18597 14456 18602 14512
rect 18658 14456 27538 14512
rect 18597 14454 27538 14456
rect 18597 14451 18663 14454
rect 3601 14378 3667 14381
rect 16849 14378 16915 14381
rect 3601 14376 16915 14378
rect 3601 14320 3606 14376
rect 3662 14320 16854 14376
rect 16910 14320 16915 14376
rect 3601 14318 16915 14320
rect 3601 14315 3667 14318
rect 16849 14315 16915 14318
rect 17309 14378 17375 14381
rect 24577 14378 24643 14381
rect 17309 14376 24643 14378
rect 17309 14320 17314 14376
rect 17370 14320 24582 14376
rect 24638 14320 24643 14376
rect 17309 14318 24643 14320
rect 17309 14315 17375 14318
rect 24577 14315 24643 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 17033 14106 17099 14109
rect 23841 14106 23907 14109
rect 17033 14104 23907 14106
rect 17033 14048 17038 14104
rect 17094 14048 23846 14104
rect 23902 14048 23907 14104
rect 17033 14046 23907 14048
rect 17033 14043 17099 14046
rect 23841 14043 23907 14046
rect 0 13970 480 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 480 13910
rect 1577 13907 1643 13910
rect 3233 13970 3299 13973
rect 7097 13970 7163 13973
rect 3233 13968 7163 13970
rect 3233 13912 3238 13968
rect 3294 13912 7102 13968
rect 7158 13912 7163 13968
rect 3233 13910 7163 13912
rect 3233 13907 3299 13910
rect 7097 13907 7163 13910
rect 9397 13970 9463 13973
rect 16113 13970 16179 13973
rect 9397 13968 16179 13970
rect 9397 13912 9402 13968
rect 9458 13912 16118 13968
rect 16174 13912 16179 13968
rect 9397 13910 16179 13912
rect 9397 13907 9463 13910
rect 16113 13907 16179 13910
rect 16297 13970 16363 13973
rect 19609 13970 19675 13973
rect 16297 13968 19675 13970
rect 16297 13912 16302 13968
rect 16358 13912 19614 13968
rect 19670 13912 19675 13968
rect 16297 13910 19675 13912
rect 16297 13907 16363 13910
rect 19609 13907 19675 13910
rect 24761 13970 24827 13973
rect 27520 13970 28000 14000
rect 24761 13968 28000 13970
rect 24761 13912 24766 13968
rect 24822 13912 28000 13968
rect 24761 13910 28000 13912
rect 24761 13907 24827 13910
rect 27520 13880 28000 13910
rect 1669 13834 1735 13837
rect 4705 13834 4771 13837
rect 1669 13832 4771 13834
rect 1669 13776 1674 13832
rect 1730 13776 4710 13832
rect 4766 13776 4771 13832
rect 1669 13774 4771 13776
rect 1669 13771 1735 13774
rect 4705 13771 4771 13774
rect 9765 13834 9831 13837
rect 14365 13834 14431 13837
rect 16665 13834 16731 13837
rect 9765 13832 14431 13834
rect 9765 13776 9770 13832
rect 9826 13776 14370 13832
rect 14426 13776 14431 13832
rect 9765 13774 14431 13776
rect 9765 13771 9831 13774
rect 14365 13771 14431 13774
rect 14782 13832 16731 13834
rect 14782 13776 16670 13832
rect 16726 13776 16731 13832
rect 14782 13774 16731 13776
rect 14782 13701 14842 13774
rect 16665 13771 16731 13774
rect 2037 13698 2103 13701
rect 4613 13698 4679 13701
rect 2037 13696 4679 13698
rect 2037 13640 2042 13696
rect 2098 13640 4618 13696
rect 4674 13640 4679 13696
rect 2037 13638 4679 13640
rect 2037 13635 2103 13638
rect 4613 13635 4679 13638
rect 14733 13696 14842 13701
rect 14733 13640 14738 13696
rect 14794 13640 14842 13696
rect 14733 13638 14842 13640
rect 14733 13635 14799 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3049 13562 3115 13565
rect 9949 13562 10015 13565
rect 3049 13560 10015 13562
rect 3049 13504 3054 13560
rect 3110 13504 9954 13560
rect 10010 13504 10015 13560
rect 3049 13502 10015 13504
rect 3049 13499 3115 13502
rect 9949 13499 10015 13502
rect 20805 13562 20871 13565
rect 23473 13562 23539 13565
rect 20805 13560 23539 13562
rect 20805 13504 20810 13560
rect 20866 13504 23478 13560
rect 23534 13504 23539 13560
rect 20805 13502 23539 13504
rect 20805 13499 20871 13502
rect 23473 13499 23539 13502
rect 12157 13426 12223 13429
rect 14641 13428 14707 13429
rect 5398 13424 12223 13426
rect 5398 13368 12162 13424
rect 12218 13368 12223 13424
rect 5398 13366 12223 13368
rect 0 13290 480 13320
rect 2998 13290 3004 13292
rect 0 13230 3004 13290
rect 0 13200 480 13230
rect 2998 13228 3004 13230
rect 3068 13228 3074 13292
rect 5398 13018 5458 13366
rect 12157 13363 12223 13366
rect 14590 13364 14596 13428
rect 14660 13426 14707 13428
rect 21633 13426 21699 13429
rect 22277 13426 22343 13429
rect 14660 13424 14752 13426
rect 14702 13368 14752 13424
rect 14660 13366 14752 13368
rect 21633 13424 22343 13426
rect 21633 13368 21638 13424
rect 21694 13368 22282 13424
rect 22338 13368 22343 13424
rect 21633 13366 22343 13368
rect 14660 13364 14707 13366
rect 14641 13363 14707 13364
rect 21633 13363 21699 13366
rect 22277 13363 22343 13366
rect 10777 13290 10843 13293
rect 20437 13290 20503 13293
rect 10777 13288 20503 13290
rect 10777 13232 10782 13288
rect 10838 13232 20442 13288
rect 20498 13232 20503 13288
rect 10777 13230 20503 13232
rect 10777 13227 10843 13230
rect 20437 13227 20503 13230
rect 23841 13290 23907 13293
rect 27520 13290 28000 13320
rect 23841 13288 28000 13290
rect 23841 13232 23846 13288
rect 23902 13232 28000 13288
rect 23841 13230 28000 13232
rect 23841 13227 23907 13230
rect 27520 13200 28000 13230
rect 6678 13092 6684 13156
rect 6748 13154 6754 13156
rect 14641 13154 14707 13157
rect 6748 13152 14707 13154
rect 6748 13096 14646 13152
rect 14702 13096 14707 13152
rect 6748 13094 14707 13096
rect 6748 13092 6754 13094
rect 14641 13091 14707 13094
rect 16757 13154 16823 13157
rect 21214 13154 21220 13156
rect 16757 13152 21220 13154
rect 16757 13096 16762 13152
rect 16818 13096 21220 13152
rect 16757 13094 21220 13096
rect 16757 13091 16823 13094
rect 21214 13092 21220 13094
rect 21284 13092 21290 13156
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 1350 12958 5458 13018
rect 8753 13018 8819 13021
rect 13721 13018 13787 13021
rect 17309 13018 17375 13021
rect 23657 13018 23723 13021
rect 8753 13016 13787 13018
rect 8753 12960 8758 13016
rect 8814 12960 13726 13016
rect 13782 12960 13787 13016
rect 8753 12958 13787 12960
rect 0 12610 480 12640
rect 1350 12610 1410 12958
rect 8753 12955 8819 12958
rect 13721 12955 13787 12958
rect 15334 13016 23723 13018
rect 15334 12960 17314 13016
rect 17370 12960 23662 13016
rect 23718 12960 23723 13016
rect 15334 12958 23723 12960
rect 1853 12882 1919 12885
rect 10777 12882 10843 12885
rect 15334 12882 15394 12958
rect 17309 12955 17375 12958
rect 23657 12955 23723 12958
rect 1853 12880 10843 12882
rect 1853 12824 1858 12880
rect 1914 12824 10782 12880
rect 10838 12824 10843 12880
rect 1853 12822 10843 12824
rect 1853 12819 1919 12822
rect 10777 12819 10843 12822
rect 10918 12822 15394 12882
rect 15469 12882 15535 12885
rect 18505 12882 18571 12885
rect 15469 12880 18571 12882
rect 15469 12824 15474 12880
rect 15530 12824 18510 12880
rect 18566 12824 18571 12880
rect 15469 12822 18571 12824
rect 5073 12746 5139 12749
rect 10918 12746 10978 12822
rect 15469 12819 15535 12822
rect 18505 12819 18571 12822
rect 5073 12744 10978 12746
rect 5073 12688 5078 12744
rect 5134 12688 10978 12744
rect 5073 12686 10978 12688
rect 14641 12746 14707 12749
rect 16021 12746 16087 12749
rect 14641 12744 16087 12746
rect 14641 12688 14646 12744
rect 14702 12688 16026 12744
rect 16082 12688 16087 12744
rect 14641 12686 16087 12688
rect 5073 12683 5139 12686
rect 14641 12683 14707 12686
rect 16021 12683 16087 12686
rect 16849 12746 16915 12749
rect 19517 12746 19583 12749
rect 16849 12744 19583 12746
rect 16849 12688 16854 12744
rect 16910 12688 19522 12744
rect 19578 12688 19583 12744
rect 16849 12686 19583 12688
rect 16849 12683 16915 12686
rect 19517 12683 19583 12686
rect 0 12550 1410 12610
rect 8109 12610 8175 12613
rect 9949 12610 10015 12613
rect 8109 12608 10015 12610
rect 8109 12552 8114 12608
rect 8170 12552 9954 12608
rect 10010 12552 10015 12608
rect 8109 12550 10015 12552
rect 0 12520 480 12550
rect 8109 12547 8175 12550
rect 9949 12547 10015 12550
rect 12249 12610 12315 12613
rect 15653 12610 15719 12613
rect 12249 12608 15719 12610
rect 12249 12552 12254 12608
rect 12310 12552 15658 12608
rect 15714 12552 15719 12608
rect 12249 12550 15719 12552
rect 12249 12547 12315 12550
rect 15653 12547 15719 12550
rect 16113 12610 16179 12613
rect 18505 12610 18571 12613
rect 16113 12608 18571 12610
rect 16113 12552 16118 12608
rect 16174 12552 18510 12608
rect 18566 12552 18571 12608
rect 16113 12550 18571 12552
rect 16113 12547 16179 12550
rect 18505 12547 18571 12550
rect 24853 12610 24919 12613
rect 27520 12610 28000 12640
rect 24853 12608 28000 12610
rect 24853 12552 24858 12608
rect 24914 12552 28000 12608
rect 24853 12550 28000 12552
rect 24853 12547 24919 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 6821 12474 6887 12477
rect 9305 12474 9371 12477
rect 6821 12472 9371 12474
rect 6821 12416 6826 12472
rect 6882 12416 9310 12472
rect 9366 12416 9371 12472
rect 6821 12414 9371 12416
rect 6821 12411 6887 12414
rect 9305 12411 9371 12414
rect 10685 12474 10751 12477
rect 13537 12474 13603 12477
rect 10685 12472 13603 12474
rect 10685 12416 10690 12472
rect 10746 12416 13542 12472
rect 13598 12416 13603 12472
rect 10685 12414 13603 12416
rect 10685 12411 10751 12414
rect 13537 12411 13603 12414
rect 3325 12338 3391 12341
rect 5993 12338 6059 12341
rect 3325 12336 6059 12338
rect 3325 12280 3330 12336
rect 3386 12280 5998 12336
rect 6054 12280 6059 12336
rect 3325 12278 6059 12280
rect 3325 12275 3391 12278
rect 5993 12275 6059 12278
rect 7557 12338 7623 12341
rect 12709 12338 12775 12341
rect 14733 12338 14799 12341
rect 7557 12336 14799 12338
rect 7557 12280 7562 12336
rect 7618 12280 12714 12336
rect 12770 12280 14738 12336
rect 14794 12280 14799 12336
rect 7557 12278 14799 12280
rect 7557 12275 7623 12278
rect 12709 12275 12775 12278
rect 14733 12275 14799 12278
rect 16389 12338 16455 12341
rect 19057 12338 19123 12341
rect 16389 12336 19123 12338
rect 16389 12280 16394 12336
rect 16450 12280 19062 12336
rect 19118 12280 19123 12336
rect 16389 12278 19123 12280
rect 16389 12275 16455 12278
rect 19057 12275 19123 12278
rect 3417 12202 3483 12205
rect 7833 12202 7899 12205
rect 11513 12202 11579 12205
rect 3417 12200 6056 12202
rect 3417 12144 3422 12200
rect 3478 12144 6056 12200
rect 3417 12142 6056 12144
rect 3417 12139 3483 12142
rect 5996 12066 6056 12142
rect 7833 12200 11579 12202
rect 7833 12144 7838 12200
rect 7894 12144 11518 12200
rect 11574 12144 11579 12200
rect 7833 12142 11579 12144
rect 7833 12139 7899 12142
rect 11513 12139 11579 12142
rect 9581 12066 9647 12069
rect 10777 12066 10843 12069
rect 14549 12066 14615 12069
rect 5996 12064 10426 12066
rect 5996 12008 9586 12064
rect 9642 12008 10426 12064
rect 5996 12006 10426 12008
rect 9581 12003 9647 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 3509 11930 3575 11933
rect 0 11928 3575 11930
rect 0 11872 3514 11928
rect 3570 11872 3575 11928
rect 0 11870 3575 11872
rect 0 11840 480 11870
rect 3509 11867 3575 11870
rect 8293 11930 8359 11933
rect 9673 11930 9739 11933
rect 8293 11928 9739 11930
rect 8293 11872 8298 11928
rect 8354 11872 9678 11928
rect 9734 11872 9739 11928
rect 8293 11870 9739 11872
rect 8293 11867 8359 11870
rect 9673 11867 9739 11870
rect 9857 11930 9923 11933
rect 10133 11930 10199 11933
rect 9857 11928 10199 11930
rect 9857 11872 9862 11928
rect 9918 11872 10138 11928
rect 10194 11872 10199 11928
rect 9857 11870 10199 11872
rect 10366 11930 10426 12006
rect 10777 12064 14615 12066
rect 10777 12008 10782 12064
rect 10838 12008 14554 12064
rect 14610 12008 14615 12064
rect 10777 12006 14615 12008
rect 10777 12003 10843 12006
rect 14549 12003 14615 12006
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 10910 11930 10916 11932
rect 10366 11870 10916 11930
rect 9857 11867 9923 11870
rect 10133 11867 10199 11870
rect 10910 11868 10916 11870
rect 10980 11868 10986 11932
rect 12801 11930 12867 11933
rect 13997 11930 14063 11933
rect 27520 11930 28000 11960
rect 12801 11928 14063 11930
rect 12801 11872 12806 11928
rect 12862 11872 14002 11928
rect 14058 11872 14063 11928
rect 12801 11870 14063 11872
rect 12801 11867 12867 11870
rect 13997 11867 14063 11870
rect 24902 11870 28000 11930
rect 2313 11794 2379 11797
rect 7557 11794 7623 11797
rect 2313 11792 7623 11794
rect 2313 11736 2318 11792
rect 2374 11736 7562 11792
rect 7618 11736 7623 11792
rect 2313 11734 7623 11736
rect 2313 11731 2379 11734
rect 7557 11731 7623 11734
rect 13169 11794 13235 11797
rect 18597 11794 18663 11797
rect 13169 11792 18663 11794
rect 13169 11736 13174 11792
rect 13230 11736 18602 11792
rect 18658 11736 18663 11792
rect 13169 11734 18663 11736
rect 13169 11731 13235 11734
rect 18597 11731 18663 11734
rect 19977 11794 20043 11797
rect 24902 11794 24962 11870
rect 27520 11840 28000 11870
rect 19977 11792 24962 11794
rect 19977 11736 19982 11792
rect 20038 11736 24962 11792
rect 19977 11734 24962 11736
rect 19977 11731 20043 11734
rect 10041 11658 10107 11661
rect 21817 11658 21883 11661
rect 10041 11656 21883 11658
rect 10041 11600 10046 11656
rect 10102 11600 21822 11656
rect 21878 11600 21883 11656
rect 10041 11598 21883 11600
rect 10041 11595 10107 11598
rect 21817 11595 21883 11598
rect 6177 11522 6243 11525
rect 9857 11522 9923 11525
rect 12801 11522 12867 11525
rect 6177 11520 9923 11522
rect 6177 11464 6182 11520
rect 6238 11464 9862 11520
rect 9918 11464 9923 11520
rect 6177 11462 9923 11464
rect 6177 11459 6243 11462
rect 9857 11459 9923 11462
rect 10688 11520 12867 11522
rect 10688 11464 12806 11520
rect 12862 11464 12867 11520
rect 10688 11462 12867 11464
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 7465 11386 7531 11389
rect 10041 11386 10107 11389
rect 7465 11384 10107 11386
rect 7465 11328 7470 11384
rect 7526 11328 10046 11384
rect 10102 11328 10107 11384
rect 7465 11326 10107 11328
rect 7465 11323 7531 11326
rect 10041 11323 10107 11326
rect 0 11250 480 11280
rect 4797 11250 4863 11253
rect 7833 11250 7899 11253
rect 0 11216 2744 11250
rect 4797 11248 7899 11250
rect 0 11190 2836 11216
rect 0 11160 480 11190
rect 2684 11156 2836 11190
rect 4797 11192 4802 11248
rect 4858 11192 7838 11248
rect 7894 11192 7899 11248
rect 4797 11190 7899 11192
rect 4797 11187 4863 11190
rect 7833 11187 7899 11190
rect 8385 11250 8451 11253
rect 10688 11250 10748 11462
rect 12801 11459 12867 11462
rect 13169 11522 13235 11525
rect 18965 11522 19031 11525
rect 13169 11520 19031 11522
rect 13169 11464 13174 11520
rect 13230 11464 18970 11520
rect 19026 11464 19031 11520
rect 13169 11462 19031 11464
rect 13169 11459 13235 11462
rect 18965 11459 19031 11462
rect 21081 11522 21147 11525
rect 22277 11522 22343 11525
rect 21081 11520 22343 11522
rect 21081 11464 21086 11520
rect 21142 11464 22282 11520
rect 22338 11464 22343 11520
rect 21081 11462 22343 11464
rect 21081 11459 21147 11462
rect 22277 11459 22343 11462
rect 23657 11522 23723 11525
rect 23657 11520 23858 11522
rect 23657 11464 23662 11520
rect 23718 11464 23858 11520
rect 23657 11462 23858 11464
rect 23657 11459 23723 11462
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 11697 11386 11763 11389
rect 19241 11386 19307 11389
rect 11697 11384 19307 11386
rect 11697 11328 11702 11384
rect 11758 11328 19246 11384
rect 19302 11328 19307 11384
rect 11697 11326 19307 11328
rect 11697 11323 11763 11326
rect 19241 11323 19307 11326
rect 8385 11248 10748 11250
rect 8385 11192 8390 11248
rect 8446 11192 10748 11248
rect 8385 11190 10748 11192
rect 12801 11250 12867 11253
rect 19701 11250 19767 11253
rect 12801 11248 19767 11250
rect 12801 11192 12806 11248
rect 12862 11192 19706 11248
rect 19762 11192 19767 11248
rect 12801 11190 19767 11192
rect 23798 11250 23858 11462
rect 27520 11250 28000 11280
rect 23798 11190 28000 11250
rect 8385 11187 8451 11190
rect 12801 11187 12867 11190
rect 19701 11187 19767 11190
rect 27520 11160 28000 11190
rect 2776 11114 2836 11156
rect 18321 11114 18387 11117
rect 20345 11114 20411 11117
rect 2776 11112 20411 11114
rect 2776 11056 18326 11112
rect 18382 11056 20350 11112
rect 20406 11056 20411 11112
rect 2776 11054 20411 11056
rect 18321 11051 18387 11054
rect 20345 11051 20411 11054
rect 20529 11114 20595 11117
rect 24853 11114 24919 11117
rect 20529 11112 24919 11114
rect 20529 11056 20534 11112
rect 20590 11056 24858 11112
rect 24914 11056 24919 11112
rect 20529 11054 24919 11056
rect 20529 11051 20595 11054
rect 24853 11051 24919 11054
rect 1485 10978 1551 10981
rect 5073 10978 5139 10981
rect 1485 10976 5139 10978
rect 1485 10920 1490 10976
rect 1546 10920 5078 10976
rect 5134 10920 5139 10976
rect 1485 10918 5139 10920
rect 1485 10915 1551 10918
rect 5073 10915 5139 10918
rect 7189 10978 7255 10981
rect 8385 10978 8451 10981
rect 10041 10978 10107 10981
rect 7189 10976 10107 10978
rect 7189 10920 7194 10976
rect 7250 10920 8390 10976
rect 8446 10920 10046 10976
rect 10102 10920 10107 10976
rect 7189 10918 10107 10920
rect 7189 10915 7255 10918
rect 8385 10915 8451 10918
rect 10041 10915 10107 10918
rect 16849 10978 16915 10981
rect 20989 10978 21055 10981
rect 16849 10976 21055 10978
rect 16849 10920 16854 10976
rect 16910 10920 20994 10976
rect 21050 10920 21055 10976
rect 16849 10918 21055 10920
rect 16849 10915 16915 10918
rect 20989 10915 21055 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 3233 10842 3299 10845
rect 4889 10842 4955 10845
rect 3233 10840 4955 10842
rect 3233 10784 3238 10840
rect 3294 10784 4894 10840
rect 4950 10784 4955 10840
rect 3233 10782 4955 10784
rect 3233 10779 3299 10782
rect 4889 10779 4955 10782
rect 6269 10842 6335 10845
rect 10133 10842 10199 10845
rect 6269 10840 10199 10842
rect 6269 10784 6274 10840
rect 6330 10784 10138 10840
rect 10194 10784 10199 10840
rect 6269 10782 10199 10784
rect 6269 10779 6335 10782
rect 10133 10779 10199 10782
rect 16389 10706 16455 10709
rect 17585 10706 17651 10709
rect 25221 10706 25287 10709
rect 7606 10704 25287 10706
rect 7606 10648 16394 10704
rect 16450 10648 17590 10704
rect 17646 10648 25226 10704
rect 25282 10648 25287 10704
rect 7606 10646 25287 10648
rect 0 10570 480 10600
rect 5349 10572 5415 10573
rect 3918 10570 3924 10572
rect 0 10510 3924 10570
rect 0 10480 480 10510
rect 3918 10508 3924 10510
rect 3988 10508 3994 10572
rect 5349 10570 5396 10572
rect 5304 10568 5396 10570
rect 5304 10512 5354 10568
rect 5304 10510 5396 10512
rect 5349 10508 5396 10510
rect 5460 10508 5466 10572
rect 5349 10507 5415 10508
rect 7606 10434 7666 10646
rect 16389 10643 16455 10646
rect 17585 10643 17651 10646
rect 25221 10643 25287 10646
rect 9305 10570 9371 10573
rect 12249 10570 12315 10573
rect 23657 10570 23723 10573
rect 9305 10568 12315 10570
rect 9305 10512 9310 10568
rect 9366 10512 12254 10568
rect 12310 10512 12315 10568
rect 9305 10510 12315 10512
rect 9305 10507 9371 10510
rect 12249 10507 12315 10510
rect 17174 10568 23723 10570
rect 17174 10512 23662 10568
rect 23718 10512 23723 10568
rect 17174 10510 23723 10512
rect 1534 10374 7666 10434
rect 12157 10434 12223 10437
rect 17174 10434 17234 10510
rect 23657 10507 23723 10510
rect 24301 10570 24367 10573
rect 27520 10570 28000 10600
rect 24301 10568 28000 10570
rect 24301 10512 24306 10568
rect 24362 10512 28000 10568
rect 24301 10510 28000 10512
rect 24301 10507 24367 10510
rect 27520 10480 28000 10510
rect 12157 10432 17234 10434
rect 12157 10376 12162 10432
rect 12218 10376 17234 10432
rect 12157 10374 17234 10376
rect 23013 10434 23079 10437
rect 23749 10434 23815 10437
rect 23013 10432 23815 10434
rect 23013 10376 23018 10432
rect 23074 10376 23754 10432
rect 23810 10376 23815 10432
rect 23013 10374 23815 10376
rect 0 9890 480 9920
rect 1534 9890 1594 10374
rect 12157 10371 12223 10374
rect 23013 10371 23079 10374
rect 23749 10371 23815 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 2773 10298 2839 10301
rect 7373 10298 7439 10301
rect 2773 10296 7439 10298
rect 2773 10240 2778 10296
rect 2834 10240 7378 10296
rect 7434 10240 7439 10296
rect 2773 10238 7439 10240
rect 2773 10235 2839 10238
rect 7373 10235 7439 10238
rect 7557 10298 7623 10301
rect 9673 10298 9739 10301
rect 7557 10296 9739 10298
rect 7557 10240 7562 10296
rect 7618 10240 9678 10296
rect 9734 10240 9739 10296
rect 7557 10238 9739 10240
rect 7557 10235 7623 10238
rect 9673 10235 9739 10238
rect 10869 10298 10935 10301
rect 13169 10298 13235 10301
rect 24209 10298 24275 10301
rect 10869 10296 19442 10298
rect 10869 10240 10874 10296
rect 10930 10240 13174 10296
rect 13230 10240 19442 10296
rect 10869 10238 19442 10240
rect 10869 10235 10935 10238
rect 13169 10235 13235 10238
rect 2589 10162 2655 10165
rect 11145 10162 11211 10165
rect 2589 10160 11211 10162
rect 2589 10104 2594 10160
rect 2650 10104 11150 10160
rect 11206 10104 11211 10160
rect 2589 10102 11211 10104
rect 19382 10162 19442 10238
rect 23614 10296 24275 10298
rect 23614 10240 24214 10296
rect 24270 10240 24275 10296
rect 23614 10238 24275 10240
rect 21081 10162 21147 10165
rect 23614 10162 23674 10238
rect 24209 10235 24275 10238
rect 25221 10162 25287 10165
rect 19382 10160 23674 10162
rect 19382 10104 21086 10160
rect 21142 10104 23674 10160
rect 19382 10102 23674 10104
rect 23798 10160 25287 10162
rect 23798 10104 25226 10160
rect 25282 10104 25287 10160
rect 23798 10102 25287 10104
rect 2589 10099 2655 10102
rect 11145 10099 11211 10102
rect 21081 10099 21147 10102
rect 2865 10026 2931 10029
rect 7189 10026 7255 10029
rect 8937 10026 9003 10029
rect 2865 10024 9003 10026
rect 2865 9968 2870 10024
rect 2926 9968 7194 10024
rect 7250 9968 8942 10024
rect 8998 9968 9003 10024
rect 2865 9966 9003 9968
rect 2865 9963 2931 9966
rect 7189 9963 7255 9966
rect 8937 9963 9003 9966
rect 11145 10026 11211 10029
rect 19793 10026 19859 10029
rect 11145 10024 19859 10026
rect 11145 9968 11150 10024
rect 11206 9968 19798 10024
rect 19854 9968 19859 10024
rect 11145 9966 19859 9968
rect 11145 9963 11211 9966
rect 19750 9963 19859 9966
rect 19977 10026 20043 10029
rect 23798 10026 23858 10102
rect 25221 10099 25287 10102
rect 19977 10024 23858 10026
rect 19977 9968 19982 10024
rect 20038 9968 23858 10024
rect 19977 9966 23858 9968
rect 23982 9966 24778 10026
rect 19977 9963 20043 9966
rect 0 9830 1594 9890
rect 1945 9890 2011 9893
rect 5349 9890 5415 9893
rect 1945 9888 5415 9890
rect 1945 9832 1950 9888
rect 2006 9832 5354 9888
rect 5410 9832 5415 9888
rect 1945 9830 5415 9832
rect 0 9800 480 9830
rect 1945 9827 2011 9830
rect 5349 9827 5415 9830
rect 5993 9890 6059 9893
rect 11789 9890 11855 9893
rect 14733 9890 14799 9893
rect 5993 9888 14799 9890
rect 5993 9832 5998 9888
rect 6054 9832 11794 9888
rect 11850 9832 14738 9888
rect 14794 9832 14799 9888
rect 5993 9830 14799 9832
rect 19750 9890 19810 9963
rect 22369 9890 22435 9893
rect 19750 9888 22435 9890
rect 19750 9832 22374 9888
rect 22430 9832 22435 9888
rect 19750 9830 22435 9832
rect 5993 9827 6059 9830
rect 11789 9827 11855 9830
rect 14733 9827 14799 9830
rect 22369 9827 22435 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 3509 9754 3575 9757
rect 10869 9754 10935 9757
rect 16665 9756 16731 9757
rect 3509 9752 5458 9754
rect 3509 9696 3514 9752
rect 3570 9696 5458 9752
rect 3509 9694 5458 9696
rect 3509 9691 3575 9694
rect 5398 9618 5458 9694
rect 5996 9752 10935 9754
rect 5996 9696 10874 9752
rect 10930 9696 10935 9752
rect 5996 9694 10935 9696
rect 5996 9618 6056 9694
rect 10869 9691 10935 9694
rect 16614 9692 16620 9756
rect 16684 9754 16731 9756
rect 23982 9754 24042 9966
rect 24718 9890 24778 9966
rect 27520 9890 28000 9920
rect 24718 9830 28000 9890
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9830
rect 24277 9759 24597 9760
rect 16684 9752 24042 9754
rect 16726 9696 24042 9752
rect 16684 9694 24042 9696
rect 16684 9692 16731 9694
rect 16665 9691 16731 9692
rect 5398 9558 6056 9618
rect 7465 9618 7531 9621
rect 12525 9618 12591 9621
rect 7465 9616 12591 9618
rect 7465 9560 7470 9616
rect 7526 9560 12530 9616
rect 12586 9560 12591 9616
rect 7465 9558 12591 9560
rect 7465 9555 7531 9558
rect 12525 9555 12591 9558
rect 12893 9618 12959 9621
rect 20805 9618 20871 9621
rect 12893 9616 20871 9618
rect 12893 9560 12898 9616
rect 12954 9560 20810 9616
rect 20866 9560 20871 9616
rect 12893 9558 20871 9560
rect 12893 9555 12959 9558
rect 20805 9555 20871 9558
rect 9029 9482 9095 9485
rect 13353 9482 13419 9485
rect 9029 9480 13419 9482
rect 9029 9424 9034 9480
rect 9090 9424 13358 9480
rect 13414 9424 13419 9480
rect 9029 9422 13419 9424
rect 9029 9419 9095 9422
rect 13353 9419 13419 9422
rect 17217 9482 17283 9485
rect 20713 9482 20779 9485
rect 17217 9480 20779 9482
rect 17217 9424 17222 9480
rect 17278 9424 20718 9480
rect 20774 9424 20779 9480
rect 17217 9422 20779 9424
rect 17217 9419 17283 9422
rect 20713 9419 20779 9422
rect 10777 9348 10843 9349
rect 10726 9284 10732 9348
rect 10796 9346 10843 9348
rect 12525 9346 12591 9349
rect 15929 9346 15995 9349
rect 10796 9344 10888 9346
rect 10838 9288 10888 9344
rect 10796 9286 10888 9288
rect 12525 9344 15995 9346
rect 12525 9288 12530 9344
rect 12586 9288 15934 9344
rect 15990 9288 15995 9344
rect 12525 9286 15995 9288
rect 10796 9284 10843 9286
rect 10777 9283 10843 9284
rect 12525 9283 12591 9286
rect 15929 9283 15995 9286
rect 10277 9280 10597 9281
rect 0 9210 480 9240
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3049 9210 3115 9213
rect 14273 9212 14339 9213
rect 0 9208 3115 9210
rect 0 9152 3054 9208
rect 3110 9152 3115 9208
rect 0 9150 3115 9152
rect 0 9120 480 9150
rect 3049 9147 3115 9150
rect 14222 9148 14228 9212
rect 14292 9210 14339 9212
rect 14292 9208 14384 9210
rect 14334 9152 14384 9208
rect 14292 9150 14384 9152
rect 14292 9148 14339 9150
rect 21214 9148 21220 9212
rect 21284 9210 21290 9212
rect 21357 9210 21423 9213
rect 21284 9208 21423 9210
rect 21284 9152 21362 9208
rect 21418 9152 21423 9208
rect 21284 9150 21423 9152
rect 21284 9148 21290 9150
rect 14273 9147 14339 9148
rect 21357 9147 21423 9150
rect 24025 9210 24091 9213
rect 27520 9210 28000 9240
rect 24025 9208 28000 9210
rect 24025 9152 24030 9208
rect 24086 9152 28000 9208
rect 24025 9150 28000 9152
rect 24025 9147 24091 9150
rect 27520 9120 28000 9150
rect 2865 9074 2931 9077
rect 11697 9074 11763 9077
rect 2865 9072 11763 9074
rect 2865 9016 2870 9072
rect 2926 9016 11702 9072
rect 11758 9016 11763 9072
rect 2865 9014 11763 9016
rect 2865 9011 2931 9014
rect 11697 9011 11763 9014
rect 14825 9074 14891 9077
rect 22185 9074 22251 9077
rect 14825 9072 22251 9074
rect 14825 9016 14830 9072
rect 14886 9016 22190 9072
rect 22246 9016 22251 9072
rect 14825 9014 22251 9016
rect 14825 9011 14891 9014
rect 22185 9011 22251 9014
rect 11094 8876 11100 8940
rect 11164 8938 11170 8940
rect 12433 8938 12499 8941
rect 11164 8936 12499 8938
rect 11164 8880 12438 8936
rect 12494 8880 12499 8936
rect 11164 8878 12499 8880
rect 11164 8876 11170 8878
rect 12433 8875 12499 8878
rect 13721 8938 13787 8941
rect 19057 8938 19123 8941
rect 13721 8936 19123 8938
rect 13721 8880 13726 8936
rect 13782 8880 19062 8936
rect 19118 8880 19123 8936
rect 13721 8878 19123 8880
rect 13721 8875 13787 8878
rect 19057 8875 19123 8878
rect 8293 8802 8359 8805
rect 13445 8802 13511 8805
rect 8293 8800 13511 8802
rect 8293 8744 8298 8800
rect 8354 8744 13450 8800
rect 13506 8744 13511 8800
rect 8293 8742 13511 8744
rect 8293 8739 8359 8742
rect 13445 8739 13511 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 7925 8666 7991 8669
rect 15929 8666 15995 8669
rect 20437 8666 20503 8669
rect 7925 8664 12266 8666
rect 7925 8608 7930 8664
rect 7986 8608 12266 8664
rect 7925 8606 12266 8608
rect 7925 8603 7991 8606
rect 0 8530 480 8560
rect 7465 8530 7531 8533
rect 8477 8530 8543 8533
rect 0 8528 7531 8530
rect 0 8472 7470 8528
rect 7526 8472 7531 8528
rect 0 8470 7531 8472
rect 0 8440 480 8470
rect 7465 8467 7531 8470
rect 7974 8528 8543 8530
rect 7974 8472 8482 8528
rect 8538 8472 8543 8528
rect 7974 8470 8543 8472
rect 2037 8394 2103 8397
rect 7974 8394 8034 8470
rect 8477 8467 8543 8470
rect 9949 8530 10015 8533
rect 11973 8530 12039 8533
rect 9949 8528 12039 8530
rect 9949 8472 9954 8528
rect 10010 8472 11978 8528
rect 12034 8472 12039 8528
rect 9949 8470 12039 8472
rect 9949 8467 10015 8470
rect 11973 8467 12039 8470
rect 2037 8392 8034 8394
rect 2037 8336 2042 8392
rect 2098 8336 8034 8392
rect 2037 8334 8034 8336
rect 10041 8394 10107 8397
rect 11237 8394 11303 8397
rect 10041 8392 11303 8394
rect 10041 8336 10046 8392
rect 10102 8336 11242 8392
rect 11298 8336 11303 8392
rect 10041 8334 11303 8336
rect 12206 8394 12266 8606
rect 15929 8664 20503 8666
rect 15929 8608 15934 8664
rect 15990 8608 20442 8664
rect 20498 8608 20503 8664
rect 15929 8606 20503 8608
rect 15929 8603 15995 8606
rect 20437 8603 20503 8606
rect 12433 8530 12499 8533
rect 17217 8530 17283 8533
rect 12433 8528 17283 8530
rect 12433 8472 12438 8528
rect 12494 8472 17222 8528
rect 17278 8472 17283 8528
rect 12433 8470 17283 8472
rect 12433 8467 12499 8470
rect 17217 8467 17283 8470
rect 19057 8530 19123 8533
rect 25497 8530 25563 8533
rect 27520 8530 28000 8560
rect 19057 8528 25563 8530
rect 19057 8472 19062 8528
rect 19118 8472 25502 8528
rect 25558 8472 25563 8528
rect 19057 8470 25563 8472
rect 19057 8467 19123 8470
rect 25497 8467 25563 8470
rect 25638 8470 28000 8530
rect 13905 8394 13971 8397
rect 14825 8394 14891 8397
rect 12206 8392 14891 8394
rect 12206 8336 13910 8392
rect 13966 8336 14830 8392
rect 14886 8336 14891 8392
rect 12206 8334 14891 8336
rect 2037 8331 2103 8334
rect 10041 8331 10107 8334
rect 11237 8331 11303 8334
rect 13905 8331 13971 8334
rect 14825 8331 14891 8334
rect 19241 8394 19307 8397
rect 22001 8394 22067 8397
rect 19241 8392 22067 8394
rect 19241 8336 19246 8392
rect 19302 8336 22006 8392
rect 22062 8336 22067 8392
rect 19241 8334 22067 8336
rect 19241 8331 19307 8334
rect 22001 8331 22067 8334
rect 23657 8394 23723 8397
rect 25638 8394 25698 8470
rect 27520 8440 28000 8470
rect 23657 8392 25698 8394
rect 23657 8336 23662 8392
rect 23718 8336 25698 8392
rect 23657 8334 25698 8336
rect 23657 8331 23723 8334
rect 3601 8258 3667 8261
rect 9857 8258 9923 8261
rect 3601 8256 9923 8258
rect 3601 8200 3606 8256
rect 3662 8200 9862 8256
rect 9918 8200 9923 8256
rect 3601 8198 9923 8200
rect 3601 8195 3667 8198
rect 9857 8195 9923 8198
rect 10685 8258 10751 8261
rect 13721 8258 13787 8261
rect 10685 8256 13787 8258
rect 10685 8200 10690 8256
rect 10746 8200 13726 8256
rect 13782 8200 13787 8256
rect 10685 8198 13787 8200
rect 10685 8195 10751 8198
rect 13721 8195 13787 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 4061 8122 4127 8125
rect 5533 8122 5599 8125
rect 5809 8122 5875 8125
rect 4061 8120 5875 8122
rect 4061 8064 4066 8120
rect 4122 8064 5538 8120
rect 5594 8064 5814 8120
rect 5870 8064 5875 8120
rect 4061 8062 5875 8064
rect 4061 8059 4127 8062
rect 5533 8059 5599 8062
rect 5809 8059 5875 8062
rect 11237 8122 11303 8125
rect 12985 8122 13051 8125
rect 11237 8120 13051 8122
rect 11237 8064 11242 8120
rect 11298 8064 12990 8120
rect 13046 8064 13051 8120
rect 11237 8062 13051 8064
rect 11237 8059 11303 8062
rect 12985 8059 13051 8062
rect 2589 7986 2655 7989
rect 9673 7986 9739 7989
rect 2589 7984 9739 7986
rect 2589 7928 2594 7984
rect 2650 7928 9678 7984
rect 9734 7928 9739 7984
rect 2589 7926 9739 7928
rect 2589 7923 2655 7926
rect 9673 7923 9739 7926
rect 10133 7986 10199 7989
rect 17309 7986 17375 7989
rect 10133 7984 17375 7986
rect 10133 7928 10138 7984
rect 10194 7928 17314 7984
rect 17370 7928 17375 7984
rect 10133 7926 17375 7928
rect 10133 7923 10199 7926
rect 17309 7923 17375 7926
rect 22737 7986 22803 7989
rect 25221 7986 25287 7989
rect 22737 7984 25287 7986
rect 22737 7928 22742 7984
rect 22798 7928 25226 7984
rect 25282 7928 25287 7984
rect 22737 7926 25287 7928
rect 22737 7923 22803 7926
rect 25221 7923 25287 7926
rect 0 7850 480 7880
rect 4429 7850 4495 7853
rect 12157 7850 12223 7853
rect 0 7848 4495 7850
rect 0 7792 4434 7848
rect 4490 7792 4495 7848
rect 0 7790 4495 7792
rect 0 7760 480 7790
rect 4429 7787 4495 7790
rect 5398 7848 12223 7850
rect 5398 7792 12162 7848
rect 12218 7792 12223 7848
rect 5398 7790 12223 7792
rect 3693 7714 3759 7717
rect 5398 7714 5458 7790
rect 12157 7787 12223 7790
rect 16849 7850 16915 7853
rect 23473 7850 23539 7853
rect 16849 7848 23539 7850
rect 16849 7792 16854 7848
rect 16910 7792 23478 7848
rect 23534 7792 23539 7848
rect 16849 7790 23539 7792
rect 16849 7787 16915 7790
rect 23473 7787 23539 7790
rect 24669 7850 24735 7853
rect 27520 7850 28000 7880
rect 24669 7848 28000 7850
rect 24669 7792 24674 7848
rect 24730 7792 28000 7848
rect 24669 7790 28000 7792
rect 24669 7787 24735 7790
rect 27520 7760 28000 7790
rect 22829 7714 22895 7717
rect 3693 7712 5458 7714
rect 3693 7656 3698 7712
rect 3754 7656 5458 7712
rect 3693 7654 5458 7656
rect 19934 7712 22895 7714
rect 19934 7656 22834 7712
rect 22890 7656 22895 7712
rect 19934 7654 22895 7656
rect 3693 7651 3759 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 1669 7578 1735 7581
rect 7649 7578 7715 7581
rect 11789 7578 11855 7581
rect 1669 7576 4170 7578
rect 1669 7520 1674 7576
rect 1730 7520 4170 7576
rect 1669 7518 4170 7520
rect 1669 7515 1735 7518
rect 4110 7445 4170 7518
rect 7649 7576 11855 7578
rect 7649 7520 7654 7576
rect 7710 7520 11794 7576
rect 11850 7520 11855 7576
rect 7649 7518 11855 7520
rect 7649 7515 7715 7518
rect 11789 7515 11855 7518
rect 18413 7578 18479 7581
rect 19609 7578 19675 7581
rect 19934 7578 19994 7654
rect 22829 7651 22895 7654
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 18413 7576 19994 7578
rect 18413 7520 18418 7576
rect 18474 7520 19614 7576
rect 19670 7520 19994 7576
rect 18413 7518 19994 7520
rect 21265 7578 21331 7581
rect 24025 7578 24091 7581
rect 21265 7576 24091 7578
rect 21265 7520 21270 7576
rect 21326 7520 24030 7576
rect 24086 7520 24091 7576
rect 21265 7518 24091 7520
rect 18413 7515 18479 7518
rect 19609 7515 19675 7518
rect 21265 7515 21331 7518
rect 24025 7515 24091 7518
rect 3693 7442 3759 7445
rect 1534 7440 3759 7442
rect 1534 7384 3698 7440
rect 3754 7384 3759 7440
rect 1534 7382 3759 7384
rect 4110 7442 4219 7445
rect 9305 7442 9371 7445
rect 12065 7442 12131 7445
rect 4110 7440 8218 7442
rect 4110 7384 4158 7440
rect 4214 7384 8218 7440
rect 4110 7382 8218 7384
rect 0 7170 480 7200
rect 1534 7170 1594 7382
rect 3693 7379 3759 7382
rect 4153 7379 4219 7382
rect 1945 7306 2011 7309
rect 8017 7306 8083 7309
rect 1945 7304 8083 7306
rect 1945 7248 1950 7304
rect 2006 7248 8022 7304
rect 8078 7248 8083 7304
rect 1945 7246 8083 7248
rect 8158 7306 8218 7382
rect 9305 7440 12131 7442
rect 9305 7384 9310 7440
rect 9366 7384 12070 7440
rect 12126 7384 12131 7440
rect 9305 7382 12131 7384
rect 9305 7379 9371 7382
rect 12065 7379 12131 7382
rect 16665 7442 16731 7445
rect 22645 7442 22711 7445
rect 16665 7440 22711 7442
rect 16665 7384 16670 7440
rect 16726 7384 22650 7440
rect 22706 7384 22711 7440
rect 16665 7382 22711 7384
rect 16665 7379 16731 7382
rect 22645 7379 22711 7382
rect 20161 7306 20227 7309
rect 8158 7304 20227 7306
rect 8158 7248 20166 7304
rect 20222 7248 20227 7304
rect 8158 7246 20227 7248
rect 1945 7243 2011 7246
rect 8017 7243 8083 7246
rect 20161 7243 20227 7246
rect 0 7110 1594 7170
rect 4889 7170 4955 7173
rect 7097 7170 7163 7173
rect 4889 7168 7163 7170
rect 4889 7112 4894 7168
rect 4950 7112 7102 7168
rect 7158 7112 7163 7168
rect 4889 7110 7163 7112
rect 0 7080 480 7110
rect 4889 7107 4955 7110
rect 7097 7107 7163 7110
rect 15561 7170 15627 7173
rect 17953 7170 18019 7173
rect 27520 7170 28000 7200
rect 15561 7168 18019 7170
rect 15561 7112 15566 7168
rect 15622 7112 17958 7168
rect 18014 7112 18019 7168
rect 15561 7110 18019 7112
rect 15561 7107 15627 7110
rect 17953 7107 18019 7110
rect 20118 7110 28000 7170
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2681 7034 2747 7037
rect 6361 7034 6427 7037
rect 2681 7032 6427 7034
rect 2681 6976 2686 7032
rect 2742 6976 6366 7032
rect 6422 6976 6427 7032
rect 2681 6974 6427 6976
rect 2681 6971 2747 6974
rect 6361 6971 6427 6974
rect 12801 7034 12867 7037
rect 18873 7034 18939 7037
rect 12801 7032 18939 7034
rect 12801 6976 12806 7032
rect 12862 6976 18878 7032
rect 18934 6976 18939 7032
rect 12801 6974 18939 6976
rect 12801 6971 12867 6974
rect 18873 6971 18939 6974
rect 2865 6898 2931 6901
rect 10685 6900 10751 6901
rect 10685 6898 10732 6900
rect 2865 6896 10732 6898
rect 10796 6898 10802 6900
rect 11053 6898 11119 6901
rect 12985 6898 13051 6901
rect 15929 6898 15995 6901
rect 2865 6840 2870 6896
rect 2926 6840 10690 6896
rect 2865 6838 10732 6840
rect 2865 6835 2931 6838
rect 10685 6836 10732 6838
rect 10796 6838 10878 6898
rect 11053 6896 15995 6898
rect 11053 6840 11058 6896
rect 11114 6840 12990 6896
rect 13046 6840 15934 6896
rect 15990 6840 15995 6896
rect 11053 6838 15995 6840
rect 10796 6836 10802 6838
rect 10685 6835 10751 6836
rect 11053 6835 11119 6838
rect 12985 6835 13051 6838
rect 15929 6835 15995 6838
rect 17677 6898 17743 6901
rect 20118 6898 20178 7110
rect 27520 7080 28000 7110
rect 23749 7034 23815 7037
rect 25405 7034 25471 7037
rect 23749 7032 25471 7034
rect 23749 6976 23754 7032
rect 23810 6976 25410 7032
rect 25466 6976 25471 7032
rect 23749 6974 25471 6976
rect 23749 6971 23815 6974
rect 25405 6971 25471 6974
rect 17677 6896 20178 6898
rect 17677 6840 17682 6896
rect 17738 6840 20178 6896
rect 17677 6838 20178 6840
rect 17677 6835 17743 6838
rect 1577 6762 1643 6765
rect 14825 6762 14891 6765
rect 1577 6760 14891 6762
rect 1577 6704 1582 6760
rect 1638 6704 14830 6760
rect 14886 6704 14891 6760
rect 1577 6702 14891 6704
rect 1577 6699 1643 6702
rect 14825 6699 14891 6702
rect 15101 6762 15167 6765
rect 24853 6762 24919 6765
rect 15101 6760 24919 6762
rect 15101 6704 15106 6760
rect 15162 6704 24858 6760
rect 24914 6704 24919 6760
rect 15101 6702 24919 6704
rect 15101 6699 15167 6702
rect 24853 6699 24919 6702
rect 19336 6566 23536 6626
rect 5610 6560 5930 6561
rect 0 6490 480 6520
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 3601 6490 3667 6493
rect 13353 6492 13419 6493
rect 0 6488 3667 6490
rect 0 6432 3606 6488
rect 3662 6432 3667 6488
rect 0 6430 3667 6432
rect 0 6400 480 6430
rect 3601 6427 3667 6430
rect 13302 6428 13308 6492
rect 13372 6490 13419 6492
rect 16665 6490 16731 6493
rect 19336 6490 19396 6566
rect 13372 6488 13464 6490
rect 13414 6432 13464 6488
rect 13372 6430 13464 6432
rect 16665 6488 19396 6490
rect 16665 6432 16670 6488
rect 16726 6432 19396 6488
rect 16665 6430 19396 6432
rect 13372 6428 13419 6430
rect 13353 6427 13419 6428
rect 16665 6427 16731 6430
rect 6637 6354 6703 6357
rect 10501 6354 10567 6357
rect 6637 6352 10567 6354
rect 6637 6296 6642 6352
rect 6698 6296 10506 6352
rect 10562 6296 10567 6352
rect 6637 6294 10567 6296
rect 6637 6291 6703 6294
rect 10501 6291 10567 6294
rect 17493 6354 17559 6357
rect 19333 6354 19399 6357
rect 17493 6352 19399 6354
rect 17493 6296 17498 6352
rect 17554 6296 19338 6352
rect 19394 6296 19399 6352
rect 17493 6294 19399 6296
rect 23476 6354 23536 6566
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 27520 6490 28000 6520
rect 24672 6430 28000 6490
rect 24672 6354 24732 6430
rect 27520 6400 28000 6430
rect 23476 6294 24732 6354
rect 17493 6291 17559 6294
rect 19333 6291 19399 6294
rect 5625 6218 5691 6221
rect 8937 6218 9003 6221
rect 5625 6216 9003 6218
rect 5625 6160 5630 6216
rect 5686 6160 8942 6216
rect 8998 6160 9003 6216
rect 5625 6158 9003 6160
rect 5625 6155 5691 6158
rect 8937 6155 9003 6158
rect 11329 6218 11395 6221
rect 15285 6218 15351 6221
rect 19333 6218 19399 6221
rect 11329 6216 19399 6218
rect 11329 6160 11334 6216
rect 11390 6160 15290 6216
rect 15346 6160 19338 6216
rect 19394 6160 19399 6216
rect 11329 6158 19399 6160
rect 11329 6155 11395 6158
rect 15285 6155 15351 6158
rect 19333 6155 19399 6158
rect 1485 6082 1551 6085
rect 2681 6082 2747 6085
rect 13721 6082 13787 6085
rect 18965 6082 19031 6085
rect 1485 6080 7666 6082
rect 1485 6024 1490 6080
rect 1546 6024 2686 6080
rect 2742 6024 7666 6080
rect 1485 6022 7666 6024
rect 1485 6019 1551 6022
rect 2681 6019 2747 6022
rect 0 5810 480 5840
rect 3969 5810 4035 5813
rect 0 5808 4035 5810
rect 0 5752 3974 5808
rect 4030 5752 4035 5808
rect 0 5750 4035 5752
rect 7606 5810 7666 6022
rect 13721 6080 19031 6082
rect 13721 6024 13726 6080
rect 13782 6024 18970 6080
rect 19026 6024 19031 6080
rect 13721 6022 19031 6024
rect 13721 6019 13787 6022
rect 18965 6019 19031 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 10688 5886 17234 5946
rect 10688 5810 10748 5886
rect 12893 5810 12959 5813
rect 7606 5750 10748 5810
rect 10918 5808 12959 5810
rect 10918 5752 12898 5808
rect 12954 5752 12959 5808
rect 10918 5750 12959 5752
rect 17174 5810 17234 5886
rect 24209 5810 24275 5813
rect 17174 5808 24275 5810
rect 17174 5752 24214 5808
rect 24270 5752 24275 5808
rect 17174 5750 24275 5752
rect 0 5720 480 5750
rect 3969 5747 4035 5750
rect 3969 5674 4035 5677
rect 5165 5674 5231 5677
rect 6269 5674 6335 5677
rect 10918 5674 10978 5750
rect 12893 5747 12959 5750
rect 24209 5747 24275 5750
rect 24853 5810 24919 5813
rect 27520 5810 28000 5840
rect 24853 5808 28000 5810
rect 24853 5752 24858 5808
rect 24914 5752 28000 5808
rect 24853 5750 28000 5752
rect 24853 5747 24919 5750
rect 27520 5720 28000 5750
rect 3969 5672 6335 5674
rect 3969 5616 3974 5672
rect 4030 5616 5170 5672
rect 5226 5616 6274 5672
rect 6330 5616 6335 5672
rect 3969 5614 6335 5616
rect 3969 5611 4035 5614
rect 5165 5611 5231 5614
rect 6269 5611 6335 5614
rect 6456 5614 10978 5674
rect 11697 5674 11763 5677
rect 19057 5674 19123 5677
rect 19609 5674 19675 5677
rect 11697 5672 19675 5674
rect 11697 5616 11702 5672
rect 11758 5616 19062 5672
rect 19118 5616 19614 5672
rect 19670 5616 19675 5672
rect 11697 5614 19675 5616
rect 5993 5538 6059 5541
rect 6456 5538 6516 5614
rect 11697 5611 11763 5614
rect 19057 5611 19123 5614
rect 19609 5611 19675 5614
rect 5993 5536 6516 5538
rect 5993 5480 5998 5536
rect 6054 5480 6516 5536
rect 5993 5478 6516 5480
rect 8385 5538 8451 5541
rect 10133 5538 10199 5541
rect 11329 5538 11395 5541
rect 8385 5536 11395 5538
rect 8385 5480 8390 5536
rect 8446 5480 10138 5536
rect 10194 5480 11334 5536
rect 11390 5480 11395 5536
rect 8385 5478 11395 5480
rect 5993 5475 6059 5478
rect 8385 5475 8451 5478
rect 10133 5475 10199 5478
rect 11329 5475 11395 5478
rect 12934 5476 12940 5540
rect 13004 5538 13010 5540
rect 13629 5538 13695 5541
rect 13004 5536 13695 5538
rect 13004 5480 13634 5536
rect 13690 5480 13695 5536
rect 13004 5478 13695 5480
rect 13004 5476 13010 5478
rect 13629 5475 13695 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 10777 5402 10843 5405
rect 13537 5402 13603 5405
rect 10777 5400 13603 5402
rect 10777 5344 10782 5400
rect 10838 5344 13542 5400
rect 13598 5344 13603 5400
rect 10777 5342 13603 5344
rect 10777 5339 10843 5342
rect 13537 5339 13603 5342
rect 10317 5266 10383 5269
rect 16481 5266 16547 5269
rect 10317 5264 16547 5266
rect 10317 5208 10322 5264
rect 10378 5208 16486 5264
rect 16542 5208 16547 5264
rect 10317 5206 16547 5208
rect 10317 5203 10383 5206
rect 16481 5203 16547 5206
rect 20805 5266 20871 5269
rect 23657 5266 23723 5269
rect 20805 5264 23723 5266
rect 20805 5208 20810 5264
rect 20866 5208 23662 5264
rect 23718 5208 23723 5264
rect 20805 5206 23723 5208
rect 20805 5203 20871 5206
rect 23657 5203 23723 5206
rect 0 5130 480 5160
rect 1485 5130 1551 5133
rect 0 5128 1551 5130
rect 0 5072 1490 5128
rect 1546 5072 1551 5128
rect 0 5070 1551 5072
rect 0 5040 480 5070
rect 1485 5067 1551 5070
rect 2589 5130 2655 5133
rect 5809 5130 5875 5133
rect 2589 5128 5875 5130
rect 2589 5072 2594 5128
rect 2650 5072 5814 5128
rect 5870 5072 5875 5128
rect 2589 5070 5875 5072
rect 2589 5067 2655 5070
rect 5809 5067 5875 5070
rect 6361 5130 6427 5133
rect 6494 5130 6500 5132
rect 6361 5128 6500 5130
rect 6361 5072 6366 5128
rect 6422 5072 6500 5128
rect 6361 5070 6500 5072
rect 6361 5067 6427 5070
rect 6494 5068 6500 5070
rect 6564 5068 6570 5132
rect 6729 5130 6795 5133
rect 11513 5130 11579 5133
rect 6729 5128 11579 5130
rect 6729 5072 6734 5128
rect 6790 5072 11518 5128
rect 11574 5072 11579 5128
rect 6729 5070 11579 5072
rect 6729 5067 6795 5070
rect 11513 5067 11579 5070
rect 12617 5130 12683 5133
rect 20069 5130 20135 5133
rect 12617 5128 20135 5130
rect 12617 5072 12622 5128
rect 12678 5072 20074 5128
rect 20130 5072 20135 5128
rect 12617 5070 20135 5072
rect 12617 5067 12683 5070
rect 20069 5067 20135 5070
rect 23473 5130 23539 5133
rect 27520 5130 28000 5160
rect 23473 5128 28000 5130
rect 23473 5072 23478 5128
rect 23534 5072 28000 5128
rect 23473 5070 28000 5072
rect 23473 5067 23539 5070
rect 27520 5040 28000 5070
rect 2129 4994 2195 4997
rect 7465 4994 7531 4997
rect 8293 4994 8359 4997
rect 2129 4992 8359 4994
rect 2129 4936 2134 4992
rect 2190 4936 7470 4992
rect 7526 4936 8298 4992
rect 8354 4936 8359 4992
rect 2129 4934 8359 4936
rect 2129 4931 2195 4934
rect 7465 4931 7531 4934
rect 8293 4931 8359 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 1945 4858 2011 4861
rect 2497 4858 2563 4861
rect 5533 4858 5599 4861
rect 1945 4856 5599 4858
rect 1945 4800 1950 4856
rect 2006 4800 2502 4856
rect 2558 4800 5538 4856
rect 5594 4800 5599 4856
rect 1945 4798 5599 4800
rect 1945 4795 2011 4798
rect 2497 4795 2563 4798
rect 5533 4795 5599 4798
rect 5809 4858 5875 4861
rect 10777 4858 10843 4861
rect 19425 4858 19491 4861
rect 5809 4856 6194 4858
rect 5809 4800 5814 4856
rect 5870 4800 6194 4856
rect 5809 4798 6194 4800
rect 5809 4795 5875 4798
rect 0 4450 480 4480
rect 5349 4450 5415 4453
rect 0 4448 5415 4450
rect 0 4392 5354 4448
rect 5410 4392 5415 4448
rect 0 4390 5415 4392
rect 6134 4450 6194 4798
rect 10777 4856 19491 4858
rect 10777 4800 10782 4856
rect 10838 4800 19430 4856
rect 19486 4800 19491 4856
rect 10777 4798 19491 4800
rect 10777 4795 10843 4798
rect 19425 4795 19491 4798
rect 6637 4722 6703 4725
rect 9673 4722 9739 4725
rect 6637 4720 9739 4722
rect 6637 4664 6642 4720
rect 6698 4664 9678 4720
rect 9734 4664 9739 4720
rect 6637 4662 9739 4664
rect 6637 4659 6703 4662
rect 9673 4659 9739 4662
rect 11329 4586 11395 4589
rect 15009 4586 15075 4589
rect 11329 4584 15075 4586
rect 11329 4528 11334 4584
rect 11390 4528 15014 4584
rect 15070 4528 15075 4584
rect 11329 4526 15075 4528
rect 11329 4523 11395 4526
rect 15009 4523 15075 4526
rect 12893 4450 12959 4453
rect 6134 4448 12959 4450
rect 6134 4392 12898 4448
rect 12954 4392 12959 4448
rect 6134 4390 12959 4392
rect 0 4360 480 4390
rect 5349 4387 5415 4390
rect 12893 4387 12959 4390
rect 24761 4450 24827 4453
rect 27520 4450 28000 4480
rect 24761 4448 28000 4450
rect 24761 4392 24766 4448
rect 24822 4392 28000 4448
rect 24761 4390 28000 4392
rect 24761 4387 24827 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 10910 4252 10916 4316
rect 10980 4314 10986 4316
rect 12157 4314 12223 4317
rect 10980 4312 12223 4314
rect 10980 4256 12162 4312
rect 12218 4256 12223 4312
rect 10980 4254 12223 4256
rect 10980 4252 10986 4254
rect 12157 4251 12223 4254
rect 3785 4178 3851 4181
rect 5533 4178 5599 4181
rect 7925 4178 7991 4181
rect 3785 4176 7991 4178
rect 3785 4120 3790 4176
rect 3846 4120 5538 4176
rect 5594 4120 7930 4176
rect 7986 4120 7991 4176
rect 3785 4118 7991 4120
rect 3785 4115 3851 4118
rect 5533 4115 5599 4118
rect 7925 4115 7991 4118
rect 8293 4178 8359 4181
rect 20253 4178 20319 4181
rect 8293 4176 20319 4178
rect 8293 4120 8298 4176
rect 8354 4120 20258 4176
rect 20314 4120 20319 4176
rect 8293 4118 20319 4120
rect 8293 4115 8359 4118
rect 20253 4115 20319 4118
rect 20989 4178 21055 4181
rect 22369 4178 22435 4181
rect 20989 4176 22435 4178
rect 20989 4120 20994 4176
rect 21050 4120 22374 4176
rect 22430 4120 22435 4176
rect 20989 4118 22435 4120
rect 20989 4115 21055 4118
rect 22369 4115 22435 4118
rect 23197 4178 23263 4181
rect 25313 4178 25379 4181
rect 23197 4176 25379 4178
rect 23197 4120 23202 4176
rect 23258 4120 25318 4176
rect 25374 4120 25379 4176
rect 23197 4118 25379 4120
rect 23197 4115 23263 4118
rect 25313 4115 25379 4118
rect 3417 4042 3483 4045
rect 1350 4040 3483 4042
rect 1350 3984 3422 4040
rect 3478 3984 3483 4040
rect 1350 3982 3483 3984
rect 0 3770 480 3800
rect 1350 3770 1410 3982
rect 3417 3979 3483 3982
rect 3601 4042 3667 4045
rect 10685 4042 10751 4045
rect 3601 4040 10751 4042
rect 3601 3984 3606 4040
rect 3662 3984 10690 4040
rect 10746 3984 10751 4040
rect 3601 3982 10751 3984
rect 3601 3979 3667 3982
rect 10685 3979 10751 3982
rect 11053 4042 11119 4045
rect 14641 4042 14707 4045
rect 11053 4040 14707 4042
rect 11053 3984 11058 4040
rect 11114 3984 14646 4040
rect 14702 3984 14707 4040
rect 11053 3982 14707 3984
rect 11053 3979 11119 3982
rect 14641 3979 14707 3982
rect 15469 4042 15535 4045
rect 17125 4042 17191 4045
rect 15469 4040 17191 4042
rect 15469 3984 15474 4040
rect 15530 3984 17130 4040
rect 17186 3984 17191 4040
rect 15469 3982 17191 3984
rect 15469 3979 15535 3982
rect 17125 3979 17191 3982
rect 20805 4042 20871 4045
rect 24577 4042 24643 4045
rect 20805 4040 24643 4042
rect 20805 3984 20810 4040
rect 20866 3984 24582 4040
rect 24638 3984 24643 4040
rect 20805 3982 24643 3984
rect 20805 3979 20871 3982
rect 24577 3979 24643 3982
rect 2037 3908 2103 3909
rect 2037 3906 2084 3908
rect 1992 3904 2084 3906
rect 1992 3848 2042 3904
rect 1992 3846 2084 3848
rect 2037 3844 2084 3846
rect 2148 3844 2154 3908
rect 6361 3906 6427 3909
rect 9949 3906 10015 3909
rect 6361 3904 10015 3906
rect 6361 3848 6366 3904
rect 6422 3848 9954 3904
rect 10010 3848 10015 3904
rect 6361 3846 10015 3848
rect 2037 3843 2103 3844
rect 6361 3843 6427 3846
rect 9949 3843 10015 3846
rect 10777 3906 10843 3909
rect 12433 3906 12499 3909
rect 10777 3904 12499 3906
rect 10777 3848 10782 3904
rect 10838 3848 12438 3904
rect 12494 3848 12499 3904
rect 10777 3846 12499 3848
rect 10777 3843 10843 3846
rect 12433 3843 12499 3846
rect 13261 3906 13327 3909
rect 15285 3906 15351 3909
rect 13261 3904 15351 3906
rect 13261 3848 13266 3904
rect 13322 3848 15290 3904
rect 15346 3848 15351 3904
rect 13261 3846 15351 3848
rect 13261 3843 13327 3846
rect 15285 3843 15351 3846
rect 16021 3906 16087 3909
rect 19425 3906 19491 3909
rect 16021 3904 19491 3906
rect 16021 3848 16026 3904
rect 16082 3848 19430 3904
rect 19486 3848 19491 3904
rect 16021 3846 19491 3848
rect 16021 3843 16087 3846
rect 19425 3843 19491 3846
rect 21173 3906 21239 3909
rect 23657 3906 23723 3909
rect 21173 3904 23723 3906
rect 21173 3848 21178 3904
rect 21234 3848 23662 3904
rect 23718 3848 23723 3904
rect 21173 3846 23723 3848
rect 21173 3843 21239 3846
rect 23657 3843 23723 3846
rect 23790 3844 23796 3908
rect 23860 3906 23866 3908
rect 23933 3906 23999 3909
rect 23860 3904 23999 3906
rect 23860 3848 23938 3904
rect 23994 3848 23999 3904
rect 23860 3846 23999 3848
rect 23860 3844 23866 3846
rect 23933 3843 23999 3846
rect 24301 3906 24367 3909
rect 24301 3904 26066 3906
rect 24301 3848 24306 3904
rect 24362 3848 26066 3904
rect 24301 3846 26066 3848
rect 24301 3843 24367 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3710 1410 3770
rect 2773 3770 2839 3773
rect 7649 3770 7715 3773
rect 2773 3768 7715 3770
rect 2773 3712 2778 3768
rect 2834 3712 7654 3768
rect 7710 3712 7715 3768
rect 2773 3710 7715 3712
rect 0 3680 480 3710
rect 2773 3707 2839 3710
rect 7649 3707 7715 3710
rect 7925 3770 7991 3773
rect 9857 3770 9923 3773
rect 7925 3768 9923 3770
rect 7925 3712 7930 3768
rect 7986 3712 9862 3768
rect 9918 3712 9923 3768
rect 7925 3710 9923 3712
rect 7925 3707 7991 3710
rect 9857 3707 9923 3710
rect 10685 3770 10751 3773
rect 13353 3770 13419 3773
rect 10685 3768 13419 3770
rect 10685 3712 10690 3768
rect 10746 3712 13358 3768
rect 13414 3712 13419 3768
rect 10685 3710 13419 3712
rect 10685 3707 10751 3710
rect 13353 3707 13419 3710
rect 14457 3770 14523 3773
rect 15561 3770 15627 3773
rect 14457 3768 15627 3770
rect 14457 3712 14462 3768
rect 14518 3712 15566 3768
rect 15622 3712 15627 3768
rect 14457 3710 15627 3712
rect 14457 3707 14523 3710
rect 15561 3707 15627 3710
rect 20345 3770 20411 3773
rect 21817 3770 21883 3773
rect 20345 3768 21883 3770
rect 20345 3712 20350 3768
rect 20406 3712 21822 3768
rect 21878 3712 21883 3768
rect 20345 3710 21883 3712
rect 20345 3707 20411 3710
rect 21817 3707 21883 3710
rect 22645 3770 22711 3773
rect 25865 3770 25931 3773
rect 22645 3768 25931 3770
rect 22645 3712 22650 3768
rect 22706 3712 25870 3768
rect 25926 3712 25931 3768
rect 22645 3710 25931 3712
rect 26006 3770 26066 3846
rect 27520 3770 28000 3800
rect 26006 3710 28000 3770
rect 22645 3707 22711 3710
rect 25865 3707 25931 3710
rect 27520 3680 28000 3710
rect 9581 3634 9647 3637
rect 12249 3634 12315 3637
rect 9581 3632 12315 3634
rect 9581 3576 9586 3632
rect 9642 3576 12254 3632
rect 12310 3576 12315 3632
rect 9581 3574 12315 3576
rect 9581 3571 9647 3574
rect 12249 3571 12315 3574
rect 14273 3634 14339 3637
rect 16849 3634 16915 3637
rect 14273 3632 16915 3634
rect 14273 3576 14278 3632
rect 14334 3576 16854 3632
rect 16910 3576 16915 3632
rect 14273 3574 16915 3576
rect 14273 3571 14339 3574
rect 16849 3571 16915 3574
rect 17217 3634 17283 3637
rect 24761 3634 24827 3637
rect 17217 3632 24827 3634
rect 17217 3576 17222 3632
rect 17278 3576 24766 3632
rect 24822 3576 24827 3632
rect 17217 3574 24827 3576
rect 17217 3571 17283 3574
rect 24761 3571 24827 3574
rect 1393 3498 1459 3501
rect 10133 3498 10199 3501
rect 1393 3496 10199 3498
rect 1393 3440 1398 3496
rect 1454 3440 10138 3496
rect 10194 3440 10199 3496
rect 1393 3438 10199 3440
rect 1393 3435 1459 3438
rect 10133 3435 10199 3438
rect 10961 3498 11027 3501
rect 18137 3498 18203 3501
rect 21449 3498 21515 3501
rect 10961 3496 15394 3498
rect 10961 3440 10966 3496
rect 11022 3440 15394 3496
rect 10961 3438 15394 3440
rect 10961 3435 11027 3438
rect 10869 3362 10935 3365
rect 12157 3362 12223 3365
rect 14273 3362 14339 3365
rect 10869 3360 11898 3362
rect 10869 3304 10874 3360
rect 10930 3304 11898 3360
rect 10869 3302 11898 3304
rect 10869 3299 10935 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 1853 3226 1919 3229
rect 3785 3226 3851 3229
rect 1853 3224 3851 3226
rect 1853 3168 1858 3224
rect 1914 3168 3790 3224
rect 3846 3168 3851 3224
rect 1853 3166 3851 3168
rect 1853 3163 1919 3166
rect 3785 3163 3851 3166
rect 6862 3164 6868 3228
rect 6932 3226 6938 3228
rect 7189 3226 7255 3229
rect 6932 3224 7255 3226
rect 6932 3168 7194 3224
rect 7250 3168 7255 3224
rect 6932 3166 7255 3168
rect 6932 3164 6938 3166
rect 7189 3163 7255 3166
rect 9949 3226 10015 3229
rect 11838 3226 11898 3302
rect 12157 3360 14339 3362
rect 12157 3304 12162 3360
rect 12218 3304 14278 3360
rect 14334 3304 14339 3360
rect 12157 3302 14339 3304
rect 15334 3362 15394 3438
rect 18137 3496 21515 3498
rect 18137 3440 18142 3496
rect 18198 3440 21454 3496
rect 21510 3440 21515 3496
rect 18137 3438 21515 3440
rect 18137 3435 18203 3438
rect 21449 3435 21515 3438
rect 22645 3498 22711 3501
rect 26509 3498 26575 3501
rect 22645 3496 26575 3498
rect 22645 3440 22650 3496
rect 22706 3440 26514 3496
rect 26570 3440 26575 3496
rect 22645 3438 26575 3440
rect 22645 3435 22711 3438
rect 26509 3435 26575 3438
rect 18321 3362 18387 3365
rect 15334 3360 18387 3362
rect 15334 3304 18326 3360
rect 18382 3304 18387 3360
rect 15334 3302 18387 3304
rect 12157 3299 12223 3302
rect 14273 3299 14339 3302
rect 18321 3299 18387 3302
rect 21265 3362 21331 3365
rect 24025 3362 24091 3365
rect 21265 3360 24091 3362
rect 21265 3304 21270 3360
rect 21326 3304 24030 3360
rect 24086 3304 24091 3360
rect 21265 3302 24091 3304
rect 21265 3299 21331 3302
rect 24025 3299 24091 3302
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 12893 3226 12959 3229
rect 9949 3224 11714 3226
rect 9949 3168 9954 3224
rect 10010 3168 11714 3224
rect 9949 3166 11714 3168
rect 11838 3224 12959 3226
rect 11838 3168 12898 3224
rect 12954 3168 12959 3224
rect 11838 3166 12959 3168
rect 9949 3163 10015 3166
rect 0 3090 480 3120
rect 2773 3090 2839 3093
rect 0 3088 2839 3090
rect 0 3032 2778 3088
rect 2834 3032 2839 3088
rect 0 3030 2839 3032
rect 0 3000 480 3030
rect 2773 3027 2839 3030
rect 3141 3090 3207 3093
rect 7097 3090 7163 3093
rect 3141 3088 7163 3090
rect 3141 3032 3146 3088
rect 3202 3032 7102 3088
rect 7158 3032 7163 3088
rect 3141 3030 7163 3032
rect 3141 3027 3207 3030
rect 7097 3027 7163 3030
rect 7281 3090 7347 3093
rect 11053 3090 11119 3093
rect 7281 3088 11119 3090
rect 7281 3032 7286 3088
rect 7342 3032 11058 3088
rect 11114 3032 11119 3088
rect 7281 3030 11119 3032
rect 7281 3027 7347 3030
rect 11053 3027 11119 3030
rect 11329 3090 11395 3093
rect 11462 3090 11468 3092
rect 11329 3088 11468 3090
rect 11329 3032 11334 3088
rect 11390 3032 11468 3088
rect 11329 3030 11468 3032
rect 11329 3027 11395 3030
rect 11462 3028 11468 3030
rect 11532 3028 11538 3092
rect 11654 3090 11714 3166
rect 12893 3163 12959 3166
rect 17033 3226 17099 3229
rect 24117 3226 24183 3229
rect 17033 3224 24183 3226
rect 17033 3168 17038 3224
rect 17094 3168 24122 3224
rect 24178 3168 24183 3224
rect 17033 3166 24183 3168
rect 17033 3163 17099 3166
rect 24117 3163 24183 3166
rect 24669 3226 24735 3229
rect 24669 3224 26250 3226
rect 24669 3168 24674 3224
rect 24730 3168 26250 3224
rect 24669 3166 26250 3168
rect 24669 3163 24735 3166
rect 19517 3090 19583 3093
rect 11654 3088 19583 3090
rect 11654 3032 19522 3088
rect 19578 3032 19583 3088
rect 11654 3030 19583 3032
rect 19517 3027 19583 3030
rect 21357 3090 21423 3093
rect 26049 3090 26115 3093
rect 21357 3088 26115 3090
rect 21357 3032 21362 3088
rect 21418 3032 26054 3088
rect 26110 3032 26115 3088
rect 21357 3030 26115 3032
rect 26190 3090 26250 3166
rect 27520 3090 28000 3120
rect 26190 3030 28000 3090
rect 21357 3027 21423 3030
rect 26049 3027 26115 3030
rect 27520 3000 28000 3030
rect 3785 2954 3851 2957
rect 6269 2954 6335 2957
rect 3785 2952 6335 2954
rect 3785 2896 3790 2952
rect 3846 2896 6274 2952
rect 6330 2896 6335 2952
rect 3785 2894 6335 2896
rect 3785 2891 3851 2894
rect 6269 2891 6335 2894
rect 9029 2954 9095 2957
rect 12157 2954 12223 2957
rect 9029 2952 12223 2954
rect 9029 2896 9034 2952
rect 9090 2896 12162 2952
rect 12218 2896 12223 2952
rect 9029 2894 12223 2896
rect 9029 2891 9095 2894
rect 12157 2891 12223 2894
rect 19241 2954 19307 2957
rect 19425 2954 19491 2957
rect 19241 2952 19491 2954
rect 19241 2896 19246 2952
rect 19302 2896 19430 2952
rect 19486 2896 19491 2952
rect 19241 2894 19491 2896
rect 19241 2891 19307 2894
rect 19425 2891 19491 2894
rect 19885 2954 19951 2957
rect 23013 2954 23079 2957
rect 19885 2952 23079 2954
rect 19885 2896 19890 2952
rect 19946 2896 23018 2952
rect 23074 2896 23079 2952
rect 19885 2894 23079 2896
rect 19885 2891 19951 2894
rect 23013 2891 23079 2894
rect 24117 2954 24183 2957
rect 24117 2952 26434 2954
rect 24117 2896 24122 2952
rect 24178 2896 26434 2952
rect 24117 2894 26434 2896
rect 24117 2891 24183 2894
rect 841 2818 907 2821
rect 6545 2818 6611 2821
rect 8109 2818 8175 2821
rect 24669 2818 24735 2821
rect 841 2816 8175 2818
rect 841 2760 846 2816
rect 902 2760 6550 2816
rect 6606 2760 8114 2816
rect 8170 2760 8175 2816
rect 841 2758 8175 2760
rect 841 2755 907 2758
rect 6545 2755 6611 2758
rect 8109 2755 8175 2758
rect 23430 2816 24735 2818
rect 23430 2760 24674 2816
rect 24730 2760 24735 2816
rect 23430 2758 24735 2760
rect 26374 2818 26434 2894
rect 27613 2818 27679 2821
rect 26374 2816 27679 2818
rect 26374 2760 27618 2816
rect 27674 2760 27679 2816
rect 26374 2758 27679 2760
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 2313 2682 2379 2685
rect 5993 2682 6059 2685
rect 2313 2680 6059 2682
rect 2313 2624 2318 2680
rect 2374 2624 5998 2680
rect 6054 2624 6059 2680
rect 2313 2622 6059 2624
rect 2313 2619 2379 2622
rect 5993 2619 6059 2622
rect 10777 2682 10843 2685
rect 11094 2682 11100 2684
rect 10777 2680 11100 2682
rect 10777 2624 10782 2680
rect 10838 2624 11100 2680
rect 10777 2622 11100 2624
rect 10777 2619 10843 2622
rect 11094 2620 11100 2622
rect 11164 2620 11170 2684
rect 15009 2682 15075 2685
rect 16849 2682 16915 2685
rect 15009 2680 16915 2682
rect 15009 2624 15014 2680
rect 15070 2624 16854 2680
rect 16910 2624 16915 2680
rect 15009 2622 16915 2624
rect 15009 2619 15075 2622
rect 16849 2619 16915 2622
rect 20713 2682 20779 2685
rect 21449 2682 21515 2685
rect 22001 2682 22067 2685
rect 20713 2680 22067 2682
rect 20713 2624 20718 2680
rect 20774 2624 21454 2680
rect 21510 2624 22006 2680
rect 22062 2624 22067 2680
rect 20713 2622 22067 2624
rect 20713 2619 20779 2622
rect 21449 2619 21515 2622
rect 22001 2619 22067 2622
rect 4613 2546 4679 2549
rect 9029 2546 9095 2549
rect 4613 2544 9095 2546
rect 4613 2488 4618 2544
rect 4674 2488 9034 2544
rect 9090 2488 9095 2544
rect 4613 2486 9095 2488
rect 4613 2483 4679 2486
rect 9029 2483 9095 2486
rect 10225 2546 10291 2549
rect 23430 2546 23490 2758
rect 24669 2755 24735 2758
rect 27613 2755 27679 2758
rect 10225 2544 23490 2546
rect 10225 2488 10230 2544
rect 10286 2488 23490 2544
rect 10225 2486 23490 2488
rect 10225 2483 10291 2486
rect 0 2410 480 2440
rect 3601 2410 3667 2413
rect 0 2408 3667 2410
rect 0 2352 3606 2408
rect 3662 2352 3667 2408
rect 0 2350 3667 2352
rect 0 2320 480 2350
rect 3601 2347 3667 2350
rect 4521 2410 4587 2413
rect 9121 2410 9187 2413
rect 16205 2410 16271 2413
rect 4521 2408 9187 2410
rect 4521 2352 4526 2408
rect 4582 2352 9126 2408
rect 9182 2352 9187 2408
rect 4521 2350 9187 2352
rect 4521 2347 4587 2350
rect 9121 2347 9187 2350
rect 14230 2408 16271 2410
rect 14230 2352 16210 2408
rect 16266 2352 16271 2408
rect 14230 2350 16271 2352
rect 10041 2274 10107 2277
rect 14230 2274 14290 2350
rect 16205 2347 16271 2350
rect 24669 2410 24735 2413
rect 27520 2410 28000 2440
rect 24669 2408 28000 2410
rect 24669 2352 24674 2408
rect 24730 2352 28000 2408
rect 24669 2350 28000 2352
rect 24669 2347 24735 2350
rect 27520 2320 28000 2350
rect 10041 2272 14290 2274
rect 10041 2216 10046 2272
rect 10102 2216 14290 2272
rect 10041 2214 14290 2216
rect 10041 2211 10107 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 2589 2002 2655 2005
rect 6361 2002 6427 2005
rect 2589 2000 6427 2002
rect 2589 1944 2594 2000
rect 2650 1944 6366 2000
rect 6422 1944 6427 2000
rect 2589 1942 6427 1944
rect 2589 1939 2655 1942
rect 6361 1939 6427 1942
rect 8753 2002 8819 2005
rect 17769 2002 17835 2005
rect 8753 2000 17835 2002
rect 8753 1944 8758 2000
rect 8814 1944 17774 2000
rect 17830 1944 17835 2000
rect 8753 1942 17835 1944
rect 8753 1939 8819 1942
rect 17769 1939 17835 1942
rect 4981 1866 5047 1869
rect 1166 1864 5047 1866
rect 1166 1808 4986 1864
rect 5042 1808 5047 1864
rect 1166 1806 5047 1808
rect 0 1730 480 1760
rect 1166 1730 1226 1806
rect 4981 1803 5047 1806
rect 7557 1866 7623 1869
rect 21081 1866 21147 1869
rect 23749 1866 23815 1869
rect 7557 1864 23815 1866
rect 7557 1808 7562 1864
rect 7618 1808 21086 1864
rect 21142 1808 23754 1864
rect 23810 1808 23815 1864
rect 7557 1806 23815 1808
rect 7557 1803 7623 1806
rect 21081 1803 21147 1806
rect 23749 1803 23815 1806
rect 0 1670 1226 1730
rect 1393 1730 1459 1733
rect 7373 1730 7439 1733
rect 16297 1730 16363 1733
rect 27520 1730 28000 1760
rect 1393 1728 16363 1730
rect 1393 1672 1398 1728
rect 1454 1672 7378 1728
rect 7434 1672 16302 1728
rect 16358 1672 16363 1728
rect 1393 1670 16363 1672
rect 0 1640 480 1670
rect 1393 1667 1459 1670
rect 7373 1667 7439 1670
rect 16297 1667 16363 1670
rect 26926 1670 28000 1730
rect 11605 1594 11671 1597
rect 16573 1594 16639 1597
rect 26926 1594 26986 1670
rect 27520 1640 28000 1670
rect 11605 1592 16639 1594
rect 11605 1536 11610 1592
rect 11666 1536 16578 1592
rect 16634 1536 16639 1592
rect 11605 1534 16639 1536
rect 11605 1531 11671 1534
rect 16573 1531 16639 1534
rect 17174 1534 26986 1594
rect 8569 1458 8635 1461
rect 17174 1458 17234 1534
rect 8569 1456 17234 1458
rect 8569 1400 8574 1456
rect 8630 1400 17234 1456
rect 8569 1398 17234 1400
rect 8569 1395 8635 1398
rect 4061 1322 4127 1325
rect 14549 1322 14615 1325
rect 4061 1320 14615 1322
rect 4061 1264 4066 1320
rect 4122 1264 14554 1320
rect 14610 1264 14615 1320
rect 4061 1262 14615 1264
rect 4061 1259 4127 1262
rect 14549 1259 14615 1262
rect 0 1050 480 1080
rect 2221 1050 2287 1053
rect 0 1048 2287 1050
rect 0 992 2226 1048
rect 2282 992 2287 1048
rect 0 990 2287 992
rect 0 960 480 990
rect 2221 987 2287 990
rect 23657 1050 23723 1053
rect 27520 1050 28000 1080
rect 23657 1048 28000 1050
rect 23657 992 23662 1048
rect 23718 992 28000 1048
rect 23657 990 28000 992
rect 23657 987 23723 990
rect 27520 960 28000 990
rect 0 370 480 400
rect 4061 370 4127 373
rect 0 368 4127 370
rect 0 312 4066 368
rect 4122 312 4127 368
rect 0 310 4127 312
rect 0 280 480 310
rect 4061 307 4127 310
rect 18965 370 19031 373
rect 27520 370 28000 400
rect 18965 368 28000 370
rect 18965 312 18970 368
rect 19026 312 28000 368
rect 18965 310 28000 312
rect 18965 307 19031 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 21220 21252 21284 21316
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 3004 13228 3068 13292
rect 14596 13424 14660 13428
rect 14596 13368 14646 13424
rect 14646 13368 14660 13424
rect 14596 13364 14660 13368
rect 6684 13092 6748 13156
rect 21220 13092 21284 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10916 11868 10980 11932
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 3924 10508 3988 10572
rect 5396 10568 5460 10572
rect 5396 10512 5410 10568
rect 5410 10512 5460 10568
rect 5396 10508 5460 10512
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 16620 9752 16684 9756
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 16620 9696 16670 9752
rect 16670 9696 16684 9752
rect 16620 9692 16684 9696
rect 10732 9344 10796 9348
rect 10732 9288 10782 9344
rect 10782 9288 10796 9344
rect 10732 9284 10796 9288
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 14228 9208 14292 9212
rect 14228 9152 14278 9208
rect 14278 9152 14292 9208
rect 14228 9148 14292 9152
rect 21220 9148 21284 9212
rect 11100 8876 11164 8940
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 10732 6896 10796 6900
rect 10732 6840 10746 6896
rect 10746 6840 10796 6896
rect 10732 6836 10796 6840
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 13308 6488 13372 6492
rect 13308 6432 13358 6488
rect 13358 6432 13372 6488
rect 13308 6428 13372 6432
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 12940 5476 13004 5540
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 6500 5068 6564 5132
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10916 4252 10980 4316
rect 2084 3904 2148 3908
rect 2084 3848 2098 3904
rect 2098 3848 2148 3904
rect 2084 3844 2148 3848
rect 23796 3844 23860 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 6868 3164 6932 3228
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 11468 3028 11532 3092
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 11100 2620 11164 2684
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 3003 13292 3069 13293
rect 3003 13228 3004 13292
rect 3068 13228 3069 13292
rect 3003 13227 3069 13228
rect 2086 3909 2146 13142
rect 3006 9298 3066 13227
rect 5610 13088 5931 14112
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 6683 13156 6749 13157
rect 6683 13092 6684 13156
rect 6748 13092 6749 13156
rect 6683 13091 6749 13092
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 3923 10572 3989 10573
rect 3923 10508 3924 10572
rect 3988 10508 3989 10572
rect 3923 10507 3989 10508
rect 3926 6578 3986 10507
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 6686 5810 6746 13091
rect 10277 12544 10597 13568
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14595 13428 14661 13429
rect 14595 13378 14596 13428
rect 14660 13378 14661 13428
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 10915 11932 10981 11933
rect 10915 11868 10916 11932
rect 10980 11868 10981 11932
rect 10915 11867 10981 11868
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10731 9348 10797 9349
rect 10731 9284 10732 9348
rect 10796 9284 10797 9348
rect 10731 9283 10797 9284
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10734 6901 10794 9283
rect 10731 6900 10797 6901
rect 10731 6836 10732 6900
rect 10796 6836 10797 6900
rect 10731 6835 10797 6836
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 6686 5750 6930 5810
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 2083 3908 2149 3909
rect 2083 3844 2084 3908
rect 2148 3844 2149 3908
rect 2083 3843 2149 3844
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 6870 3229 6930 5750
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10918 4317 10978 11867
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 21219 21316 21285 21317
rect 21219 21252 21220 21316
rect 21284 21252 21285 21316
rect 21219 21251 21285 21252
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 21222 13157 21282 21251
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 21219 13156 21285 13157
rect 21219 13092 21220 13156
rect 21284 13092 21285 13156
rect 21219 13091 21285 13092
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 11099 8940 11165 8941
rect 11099 8876 11100 8940
rect 11164 8876 11165 8940
rect 11099 8875 11165 8876
rect 10915 4316 10981 4317
rect 10915 4252 10916 4316
rect 10980 4252 10981 4316
rect 10915 4251 10981 4252
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 6867 3228 6933 3229
rect 6867 3164 6868 3228
rect 6932 3164 6933 3228
rect 6867 3163 6933 3164
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 11102 2685 11162 8875
rect 14944 8736 15264 9760
rect 16622 9757 16682 10422
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 16619 9756 16685 9757
rect 16619 9692 16620 9756
rect 16684 9692 16685 9756
rect 16619 9691 16685 9692
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 12939 5540 13005 5541
rect 12939 5476 12940 5540
rect 13004 5476 13005 5540
rect 12939 5475 13005 5476
rect 12942 5218 13002 5475
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 11099 2684 11165 2685
rect 11099 2620 11100 2684
rect 11164 2620 11165 2684
rect 11099 2619 11165 2620
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 21222 9213 21282 13091
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 21219 9212 21285 9213
rect 21219 9148 21220 9212
rect 21284 9148 21285 9212
rect 21219 9147 21285 9148
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 23795 3908 23861 3909
rect 23795 3844 23796 3908
rect 23860 3844 23861 3908
rect 23795 3843 23861 3844
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 23798 3178 23858 3843
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 1998 13142 2234 13378
rect 5310 10572 5546 10658
rect 5310 10508 5396 10572
rect 5396 10508 5460 10572
rect 5460 10508 5546 10572
rect 2918 9062 3154 9298
rect 5310 10422 5546 10508
rect 3838 6342 4074 6578
rect 14510 13364 14596 13378
rect 14596 13364 14660 13378
rect 14660 13364 14746 13378
rect 14510 13142 14746 13364
rect 6414 5132 6650 5218
rect 6414 5068 6500 5132
rect 6500 5068 6564 5132
rect 6564 5068 6650 5132
rect 6414 4982 6650 5068
rect 16534 10422 16770 10658
rect 14142 9212 14378 9298
rect 14142 9148 14228 9212
rect 14228 9148 14292 9212
rect 14292 9148 14378 9212
rect 14142 9062 14378 9148
rect 13222 6492 13458 6578
rect 13222 6428 13308 6492
rect 13308 6428 13372 6492
rect 13372 6428 13458 6492
rect 13222 6342 13458 6428
rect 12854 4982 13090 5218
rect 11382 3092 11618 3178
rect 11382 3028 11468 3092
rect 11468 3028 11532 3092
rect 11532 3028 11618 3092
rect 11382 2942 11618 3028
rect 23710 2942 23946 3178
<< metal5 >>
rect 1956 13378 14788 13420
rect 1956 13142 1998 13378
rect 2234 13142 14510 13378
rect 14746 13142 14788 13378
rect 1956 13100 14788 13142
rect 5268 10658 16812 10700
rect 5268 10422 5310 10658
rect 5546 10422 16534 10658
rect 16770 10422 16812 10658
rect 5268 10380 16812 10422
rect 2876 9298 14420 9340
rect 2876 9062 2918 9298
rect 3154 9062 14142 9298
rect 14378 9062 14420 9298
rect 2876 9020 14420 9062
rect 3796 6578 13500 6620
rect 3796 6342 3838 6578
rect 4074 6342 13222 6578
rect 13458 6342 13500 6578
rect 3796 6300 13500 6342
rect 6372 5218 13132 5260
rect 6372 4982 6414 5218
rect 6650 4982 12854 5218
rect 13090 4982 13132 5218
rect 6372 4940 13132 4982
rect 11340 3178 23988 3220
rect 11340 2942 11382 3178
rect 11618 2942 23710 3178
rect 23946 2942 23988 3178
rect 11340 2900 23988 2942
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_17
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_1_24 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_21
timestamp 1586364061
transform 1 0 3036 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _125_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_103
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _127_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_conb_1  _034_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_203
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_206
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_210
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_235
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_241
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23920 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24196 0 -1 2720
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24104 0 1 2720
box -38 -48 1786 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_260
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_264 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_0_276
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_273
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 130 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_98
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _122_
timestamp 1586364061
transform 1 0 9752 0 -1 3808
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_39.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_37.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_179
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _116_
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_35.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_236
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_240
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 1786 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_67
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_111
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_119
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_39.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_139
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_177
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_37.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_35.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_209
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_230
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24104 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_259
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_263
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_267
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_271 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_26
timestamp 1586364061
transform 1 0 3496 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_49
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_53
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_66
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_70
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_73
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _124_
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_101
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_188
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_192
timestamp 1586364061
transform 1 0 18768 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_31.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20976 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_225
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_229
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24656 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_264 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_272
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_26
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_81
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_85
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _121_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_144
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_148
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_203
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_207
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_249
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_261
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_265
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_conb_1  _038_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_26
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_22
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_45
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_111
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _058_
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_122
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  _123_
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_129
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 1786 592
use scs8hd_buf_2  _126_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_164
timestamp 1586364061
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_buf_2  _119_
timestamp 1586364061
transform 1 0 18124 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_189
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_189
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 1786 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 21068 0 -1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_225
timestamp 1586364061
transform 1 0 21804 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_221
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21620 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_31.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_254
timestamp 1586364061
transform 1 0 24472 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_248
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 24288 0 -1 5984
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24656 0 -1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 1786 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_265
timestamp 1586364061
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_273
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_track_3.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_35
timestamp 1586364061
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_73
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_101
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_124
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_181
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_234
timestamp 1586364061
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_238
timestamp 1586364061
transform 1 0 23000 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23736 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 23184 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_242
timestamp 1586364061
transform 1 0 23368 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_265
timestamp 1586364061
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 1786 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_30
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_106
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_conb_1  _057_
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_161
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 406 592
use scs8hd_buf_2  _118_
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_209
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_226
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_270
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_25
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_101
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_172
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_176
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 17664 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_234
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_238
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_244
timestamp 1586364061
transform 1 0 23552 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 1786 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_8
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_146
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23920 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 26036 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_273
timestamp 1586364061
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use scs8hd_conb_1  _066_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_51
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_173
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_2  _120_
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 406 592
use scs8hd_mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22356 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_229
timestamp 1586364061
transform 1 0 22172 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_233
timestamp 1586364061
transform 1 0 22540 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_238
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_242
timestamp 1586364061
transform 1 0 23368 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_265
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_60
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_65
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_122
timestamp 1586364061
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _056_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_165
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_161
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_195
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_207
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_203
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_215
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _117_
timestamp 1586364061
transform 1 0 20516 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_223
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_219
timestamp 1586364061
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_233
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_229
timestamp 1586364061
transform 1 0 22172 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 1786 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_270
timestamp 1586364061
transform 1 0 25944 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_60
timestamp 1586364061
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_67
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_148
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_152
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18124 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_261
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_266
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_buf_1  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_58
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_73
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_100
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_123
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_140
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 774 592
use scs8hd_conb_1  _061_
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_181
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_234
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_238
timestamp 1586364061
transform 1 0 23000 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_257
timestamp 1586364061
transform 1 0 24748 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_8
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_21
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_25
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_133
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _060_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_194
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_238
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_264
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_37
timestamp 1586364061
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_157
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_165
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_169
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _062_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_218
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_222
timestamp 1586364061
transform 1 0 21528 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_245
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_249
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 406 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_31
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_48
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_114
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_39.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 16192 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_174
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_178
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_183
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18676 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_200
timestamp 1586364061
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_conb_1  _059_
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 314 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _063_
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_221
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_buf_1  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 406 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12972 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_131
timestamp 1586364061
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 406 592
use scs8hd_mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_35.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 314 592
use scs8hd_buf_1  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_212
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_27.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_249
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_263
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_22_76
timestamp 1586364061
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_112
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_116
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_133
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_1  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_192
timestamp 1586364061
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_37.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_203
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_218
timestamp 1586364061
transform 1 0 21160 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_31.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_230
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_236
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23552 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _083_
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_20
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_26
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_70
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 406 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_157
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_161
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_buf_1  mux_bottom_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_187
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_191
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_195
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 130 592
use scs8hd_buf_1  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20148 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_199
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_203
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_210
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_226
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_249
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_48
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_101
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_124
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  mux_right_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_167
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _067_
timestamp 1586364061
transform 1 0 22540 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_8  FILLER_24_236
timestamp 1586364061
transform 1 0 22816 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  mux_bottom_track_29.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23552 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_247
timestamp 1586364061
transform 1 0 23828 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_buf_1  mux_left_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_129
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_142
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_146
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_169
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 774 592
use scs8hd_buf_1  mux_bottom_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_181
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _064_
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_25_227
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 590 592
use scs8hd_decap_8  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 774 592
use scs8hd_conb_1  _065_
timestamp 1586364061
transform 1 0 24196 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_249
timestamp 1586364061
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_254
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_270
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_85
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_99
timestamp 1586364061
transform 1 0 10212 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_90
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10304 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_173
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_172
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_185
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_197
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_209
timestamp 1586364061
transform 1 0 20332 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_1  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23552 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_243
timestamp 1586364061
transform 1 0 23460 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_271
timestamp 1586364061
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_259
timestamp 1586364061
transform 1 0 24932 0 -1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_99
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 10304 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_154
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_166
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_99
timestamp 1586364061
transform 1 0 10212 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_114
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 590 592
use scs8hd_mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_131
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_136
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 314 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_17
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_41
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_left_track_33.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_33.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_131
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_165
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_177
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_buf_1  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_133
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_136
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_148
timestamp 1586364061
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_18
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 406 592
use scs8hd_buf_1  mux_left_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_46
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_131
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_165
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_259
timestamp 1586364061
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_271
timestamp 1586364061
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 24564 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_259
timestamp 1586364061
transform 1 0 24932 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_271
timestamp 1586364061
transform 1 0 26036 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_1  mux_right_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24104 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_248
timestamp 1586364061
transform 1 0 23920 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_252
timestamp 1586364061
transform 1 0 24288 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2594 0 2650 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3790 0 3846 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 4342 0 4398 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 ccff_head
port 8 nsew default input
rlabel metal2 s 23202 27520 23258 28000 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 960 480 1080 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 1640 480 1760 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 2320 480 2440 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 24080 480 24200 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 25440 480 25560 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 26120 480 26240 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 26800 480 26920 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 15240 480 15360 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 280 28000 400 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 9120 28000 9240 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 13200 28000 13320 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 960 28000 1080 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 1640 28000 1760 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 2320 28000 2440 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 3000 28000 3120 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 5040 28000 5160 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 5720 28000 5840 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 6400 28000 6520 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 22040 28000 22160 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 22720 28000 22840 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 23400 28000 23520 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 24080 28000 24200 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 25440 28000 25560 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 26120 28000 26240 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 26800 28000 26920 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 15240 28000 15360 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 17280 28000 17400 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 18640 28000 18760 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 19320 28000 19440 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 22374 0 22430 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 23018 0 23074 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 25870 0 25926 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 19522 0 19578 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 21270 0 21326 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal3 s 0 27480 480 27600 6 left_top_grid_pin_1_
port 130 nsew default input
rlabel metal2 s 4618 27520 4674 28000 6 prog_clk
port 131 nsew default input
rlabel metal3 s 27520 27480 28000 27600 6 right_top_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
