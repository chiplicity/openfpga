magic
tech sky130A
magscale 1 2
timestamp 1608764133
<< checkpaint >>
rect -1260 -1260 18260 21260
<< locali >>
rect 7573 4063 7607 4233
rect 11713 4063 11747 4233
rect 7941 2907 7975 3009
<< viali >>
rect 4721 15657 4755 15691
rect 4537 15521 4571 15555
rect 3985 15113 4019 15147
rect 5549 15113 5583 15147
rect 3801 14909 3835 14943
rect 5365 14909 5399 14943
rect 4445 14841 4479 14875
rect 4721 14773 4755 14807
rect 6009 14773 6043 14807
rect 2789 14569 2823 14603
rect 7297 14569 7331 14603
rect 9873 14569 9907 14603
rect 6285 14433 6319 14467
rect 7113 14433 7147 14467
rect 9689 14433 9723 14467
rect 6101 14229 6135 14263
rect 14657 14025 14691 14059
rect 2789 13957 2823 13991
rect 3249 13957 3283 13991
rect 3893 13889 3927 13923
rect 3157 13821 3191 13855
rect 6285 13821 6319 13855
rect 9781 13821 9815 13855
rect 14473 13821 14507 13855
rect 15025 13821 15059 13855
rect 7205 13685 7239 13719
rect 4353 13345 4387 13379
rect 4609 13345 4643 13379
rect 5733 13141 5767 13175
rect 7481 13141 7515 13175
rect 7757 13141 7791 13175
rect 4629 12937 4663 12971
rect 5089 12937 5123 12971
rect 7481 12801 7515 12835
rect 7665 12801 7699 12835
rect 7389 12733 7423 12767
rect 7021 12597 7055 12631
rect 8125 12597 8159 12631
rect 6101 12257 6135 12291
rect 7389 12053 7423 12087
rect 8125 12053 8159 12087
rect 7573 11849 7607 11883
rect 9137 11849 9171 11883
rect 7757 11713 7791 11747
rect 8024 11645 8058 11679
rect 6193 11509 6227 11543
rect 3801 11305 3835 11339
rect 7113 11305 7147 11339
rect 8677 11305 8711 11339
rect 10149 11305 10183 11339
rect 8953 11237 8987 11271
rect 2948 11169 2982 11203
rect 6101 11169 6135 11203
rect 6745 11169 6779 11203
rect 7297 11169 7331 11203
rect 7553 11169 7587 11203
rect 10057 11169 10091 11203
rect 6193 11101 6227 11135
rect 6377 11101 6411 11135
rect 10241 11101 10275 11135
rect 5733 11033 5767 11067
rect 9689 11033 9723 11067
rect 3019 10965 3053 10999
rect 10701 10965 10735 10999
rect 2973 10761 3007 10795
rect 3525 10761 3559 10795
rect 6193 10761 6227 10795
rect 9689 10761 9723 10795
rect 6469 10693 6503 10727
rect 9781 10693 9815 10727
rect 11161 10693 11195 10727
rect 3801 10625 3835 10659
rect 10333 10625 10367 10659
rect 11345 10625 11379 10659
rect 6653 10557 6687 10591
rect 7573 10557 7607 10591
rect 9321 10557 9355 10591
rect 3893 10489 3927 10523
rect 4813 10489 4847 10523
rect 5825 10489 5859 10523
rect 7113 10489 7147 10523
rect 7840 10489 7874 10523
rect 10149 10489 10183 10523
rect 7481 10421 7515 10455
rect 8953 10421 8987 10455
rect 10241 10421 10275 10455
rect 10793 10421 10827 10455
rect 7205 10217 7239 10251
rect 8677 10217 8711 10251
rect 8953 10217 8987 10251
rect 9413 10217 9447 10251
rect 10149 10217 10183 10251
rect 1593 10149 1627 10183
rect 2513 10149 2547 10183
rect 6101 10081 6135 10115
rect 7297 10081 7331 10115
rect 7564 10081 7598 10115
rect 10057 10081 10091 10115
rect 1501 10013 1535 10047
rect 6193 10013 6227 10047
rect 6377 10013 6411 10047
rect 10241 10013 10275 10047
rect 10701 10013 10735 10047
rect 5733 9877 5767 9911
rect 6837 9877 6871 9911
rect 9689 9877 9723 9911
rect 6193 9673 6227 9707
rect 10425 9673 10459 9707
rect 6929 9605 6963 9639
rect 8309 9605 8343 9639
rect 9505 9605 9539 9639
rect 7573 9537 7607 9571
rect 9137 9537 9171 9571
rect 10793 9537 10827 9571
rect 6653 9469 6687 9503
rect 7297 9469 7331 9503
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 7389 9401 7423 9435
rect 8033 9401 8067 9435
rect 1593 9333 1627 9367
rect 1961 9333 1995 9367
rect 5825 9333 5859 9367
rect 8493 9333 8527 9367
rect 10057 9333 10091 9367
rect 7297 9129 7331 9163
rect 7665 9129 7699 9163
rect 8769 9129 8803 9163
rect 7757 9061 7791 9095
rect 8401 9061 8435 9095
rect 7205 8993 7239 9027
rect 12449 8993 12483 9027
rect 7941 8925 7975 8959
rect 12633 8925 12667 8959
rect 7389 8585 7423 8619
rect 7757 8585 7791 8619
rect 8033 8585 8067 8619
rect 8217 8517 8251 8551
rect 8861 8449 8895 8483
rect 9229 8449 9263 8483
rect 8677 8381 8711 8415
rect 8585 8313 8619 8347
rect 12725 8313 12759 8347
rect 8585 8041 8619 8075
rect 4169 7497 4203 7531
rect 3341 7293 3375 7327
rect 3617 7225 3651 7259
rect 5089 6409 5123 6443
rect 9781 6409 9815 6443
rect 9321 6341 9355 6375
rect 4905 6205 4939 6239
rect 7481 6205 7515 6239
rect 9137 6205 9171 6239
rect 8125 6137 8159 6171
rect 5549 6069 5583 6103
rect 7665 6069 7699 6103
rect 7205 5865 7239 5899
rect 9873 5865 9907 5899
rect 12173 5865 12207 5899
rect 4077 5729 4111 5763
rect 5181 5729 5215 5763
rect 7021 5729 7055 5763
rect 8125 5729 8159 5763
rect 9689 5729 9723 5763
rect 10793 5729 10827 5763
rect 11989 5729 12023 5763
rect 10977 5593 11011 5627
rect 4261 5525 4295 5559
rect 4629 5525 4663 5559
rect 5365 5525 5399 5559
rect 8309 5525 8343 5559
rect 9137 5525 9171 5559
rect 4169 5321 4203 5355
rect 5273 5321 5307 5355
rect 5825 5321 5859 5355
rect 12633 5321 12667 5355
rect 7021 5253 7055 5287
rect 7849 5253 7883 5287
rect 6285 5185 6319 5219
rect 10793 5185 10827 5219
rect 4537 5117 4571 5151
rect 5641 5117 5675 5151
rect 6837 5117 6871 5151
rect 7941 5117 7975 5151
rect 9045 5117 9079 5151
rect 10149 5117 10183 5151
rect 11253 5117 11287 5151
rect 12449 5117 12483 5151
rect 11897 5049 11931 5083
rect 4721 4981 4755 5015
rect 7481 4981 7515 5015
rect 8125 4981 8159 5015
rect 8585 4981 8619 5015
rect 8953 4981 8987 5015
rect 9229 4981 9263 5015
rect 9781 4981 9815 5015
rect 10333 4981 10367 5015
rect 11161 4981 11195 5015
rect 11437 4981 11471 5015
rect 12265 4981 12299 5015
rect 13093 4981 13127 5015
rect 8033 4777 8067 4811
rect 10149 4777 10183 4811
rect 12633 4777 12667 4811
rect 4813 4641 4847 4675
rect 5917 4641 5951 4675
rect 7849 4641 7883 4675
rect 9965 4641 9999 4675
rect 11069 4641 11103 4675
rect 12449 4641 12483 4675
rect 13553 4641 13587 4675
rect 4997 4437 5031 4471
rect 6101 4437 6135 4471
rect 11253 4437 11287 4471
rect 13737 4437 13771 4471
rect 4905 4233 4939 4267
rect 6009 4233 6043 4267
rect 7481 4233 7515 4267
rect 7573 4233 7607 4267
rect 10793 4233 10827 4267
rect 11161 4233 11195 4267
rect 11713 4233 11747 4267
rect 11897 4233 11931 4267
rect 13645 4233 13679 4267
rect 7849 4097 7883 4131
rect 9689 4097 9723 4131
rect 6837 4029 6871 4063
rect 7573 4029 7607 4063
rect 7947 4029 7981 4063
rect 9045 4029 9079 4063
rect 10149 4029 10183 4063
rect 11253 4029 11287 4063
rect 11713 4029 11747 4063
rect 12265 4029 12299 4063
rect 12449 4029 12483 4063
rect 7021 3893 7055 3927
rect 8125 3893 8159 3927
rect 8585 3893 8619 3927
rect 9229 3893 9263 3927
rect 10057 3893 10091 3927
rect 10333 3893 10367 3927
rect 11437 3893 11471 3927
rect 12633 3893 12667 3927
rect 13093 3893 13127 3927
rect 10425 3689 10459 3723
rect 6837 3553 6871 3587
rect 8125 3553 8159 3587
rect 10241 3553 10275 3587
rect 11535 3553 11569 3587
rect 8309 3417 8343 3451
rect 7021 3349 7055 3383
rect 11713 3349 11747 3383
rect 8125 3145 8159 3179
rect 11621 3145 11655 3179
rect 7941 3009 7975 3043
rect 7113 2873 7147 2907
rect 7941 2873 7975 2907
rect 10333 2805 10367 2839
<< metal1 >>
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 9858 17008 9864 17060
rect 9916 17048 9922 17060
rect 10962 17048 10968 17060
rect 9916 17020 10968 17048
rect 9916 17008 9922 17020
rect 10962 17008 10968 17020
rect 11020 17008 11026 17060
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 4890 16396 4896 16448
rect 4948 16436 4954 16448
rect 9306 16436 9312 16448
rect 4948 16408 9312 16436
rect 4948 16396 4954 16408
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9674 16396 9680 16448
rect 9732 16436 9738 16448
rect 11790 16436 11796 16448
rect 9732 16408 11796 16436
rect 9732 16396 9738 16408
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 9674 16164 9680 16176
rect 7984 16136 9680 16164
rect 7984 16124 7990 16136
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 8846 16096 8852 16108
rect 6696 16068 8852 16096
rect 6696 16056 6702 16068
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 12618 16096 12624 16108
rect 9640 16068 12624 16096
rect 9640 16056 9646 16068
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 9122 15988 9128 16040
rect 9180 16028 9186 16040
rect 12158 16028 12164 16040
rect 9180 16000 12164 16028
rect 9180 15988 9186 16000
rect 12158 15988 12164 16000
rect 12216 15988 12222 16040
rect 3694 15920 3700 15972
rect 3752 15960 3758 15972
rect 4062 15960 4068 15972
rect 3752 15932 4068 15960
rect 3752 15920 3758 15932
rect 4062 15920 4068 15932
rect 4120 15920 4126 15972
rect 5534 15920 5540 15972
rect 5592 15960 5598 15972
rect 8202 15960 8208 15972
rect 5592 15932 8208 15960
rect 5592 15920 5598 15932
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 8662 15920 8668 15972
rect 8720 15960 8726 15972
rect 9674 15960 9680 15972
rect 8720 15932 9680 15960
rect 8720 15920 8726 15932
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 1854 15852 1860 15904
rect 1912 15892 1918 15904
rect 5626 15892 5632 15904
rect 1912 15864 5632 15892
rect 1912 15852 1918 15864
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 9950 15892 9956 15904
rect 8904 15864 9956 15892
rect 8904 15852 8910 15864
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 11330 15892 11336 15904
rect 10468 15864 11336 15892
rect 10468 15852 10474 15864
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 1452 15660 4721 15688
rect 1452 15648 1458 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 10134 15688 10140 15700
rect 6512 15660 10140 15688
rect 6512 15648 6518 15660
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 10318 15648 10324 15700
rect 10376 15688 10382 15700
rect 15470 15688 15476 15700
rect 10376 15660 15476 15688
rect 10376 15648 10382 15660
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 1026 15580 1032 15632
rect 1084 15620 1090 15632
rect 1084 15592 2820 15620
rect 1084 15580 1090 15592
rect 2792 15484 2820 15592
rect 3786 15580 3792 15632
rect 3844 15620 3850 15632
rect 4062 15620 4068 15632
rect 3844 15592 4068 15620
rect 3844 15580 3850 15592
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 5074 15620 5080 15632
rect 4264 15592 5080 15620
rect 4264 15484 4292 15592
rect 5074 15580 5080 15592
rect 5132 15580 5138 15632
rect 8018 15580 8024 15632
rect 8076 15620 8082 15632
rect 10686 15620 10692 15632
rect 8076 15592 10692 15620
rect 8076 15580 8082 15592
rect 10686 15580 10692 15592
rect 10744 15580 10750 15632
rect 13630 15580 13636 15632
rect 13688 15620 13694 15632
rect 16758 15620 16764 15632
rect 13688 15592 16764 15620
rect 13688 15580 13694 15592
rect 16758 15580 16764 15592
rect 16816 15580 16822 15632
rect 4522 15552 4528 15564
rect 4483 15524 4528 15552
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 6270 15512 6276 15564
rect 6328 15552 6334 15564
rect 9950 15552 9956 15564
rect 6328 15524 9956 15552
rect 6328 15512 6334 15524
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 10134 15512 10140 15564
rect 10192 15552 10198 15564
rect 12710 15552 12716 15564
rect 10192 15524 12716 15552
rect 10192 15512 10198 15524
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 2792 15456 4292 15484
rect 7558 15444 7564 15496
rect 7616 15484 7622 15496
rect 9582 15484 9588 15496
rect 7616 15456 9588 15484
rect 7616 15444 7622 15456
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 15930 15484 15936 15496
rect 11756 15456 15936 15484
rect 11756 15444 11762 15456
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 2222 15376 2228 15428
rect 2280 15416 2286 15428
rect 5534 15416 5540 15428
rect 2280 15388 5540 15416
rect 2280 15376 2286 15388
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 11422 15376 11428 15428
rect 11480 15416 11486 15428
rect 14274 15416 14280 15428
rect 11480 15388 14280 15416
rect 11480 15376 11486 15388
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 6730 15348 6736 15360
rect 4764 15320 6736 15348
rect 4764 15308 4770 15320
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 9582 15348 9588 15360
rect 7248 15320 9588 15348
rect 7248 15308 7254 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 566 15104 572 15156
rect 624 15144 630 15156
rect 3973 15147 4031 15153
rect 3973 15144 3985 15147
rect 624 15116 3985 15144
rect 624 15104 630 15116
rect 3973 15113 3985 15116
rect 4019 15113 4031 15147
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 3973 15107 4031 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 5353 14943 5411 14949
rect 3835 14912 4476 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4448 14881 4476 14912
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5399 14912 6040 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 4433 14875 4491 14881
rect 4433 14841 4445 14875
rect 4479 14872 4491 14875
rect 5810 14872 5816 14884
rect 4479 14844 5816 14872
rect 4479 14841 4491 14844
rect 4433 14835 4491 14841
rect 5810 14832 5816 14844
rect 5868 14832 5874 14884
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 6012 14813 6040 14912
rect 4709 14807 4767 14813
rect 4709 14804 4721 14807
rect 4580 14776 4721 14804
rect 4580 14764 4586 14776
rect 4709 14773 4721 14776
rect 4755 14773 4767 14807
rect 4709 14767 4767 14773
rect 5997 14807 6055 14813
rect 5997 14773 6009 14807
rect 6043 14804 6055 14807
rect 9674 14804 9680 14816
rect 6043 14776 9680 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 198 14560 204 14612
rect 256 14600 262 14612
rect 2590 14600 2596 14612
rect 256 14572 2596 14600
rect 256 14560 262 14572
rect 2590 14560 2596 14572
rect 2648 14600 2654 14612
rect 2777 14603 2835 14609
rect 2777 14600 2789 14603
rect 2648 14572 2789 14600
rect 2648 14560 2654 14572
rect 2777 14569 2789 14572
rect 2823 14569 2835 14603
rect 2777 14563 2835 14569
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 6788 14572 7297 14600
rect 6788 14560 6794 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 7285 14563 7343 14569
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 9640 14572 9873 14600
rect 9640 14560 9646 14572
rect 9861 14569 9873 14572
rect 9907 14569 9919 14603
rect 9861 14563 9919 14569
rect 6270 14464 6276 14476
rect 6231 14436 6276 14464
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 7098 14464 7104 14476
rect 7059 14436 7104 14464
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 10042 14464 10048 14476
rect 9723 14436 10048 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 6089 14263 6147 14269
rect 6089 14260 6101 14263
rect 5592 14232 6101 14260
rect 5592 14220 5598 14232
rect 6089 14229 6101 14232
rect 6135 14229 6147 14263
rect 6089 14223 6147 14229
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 13780 14028 14657 14056
rect 13780 14016 13786 14028
rect 14645 14025 14657 14028
rect 14691 14025 14703 14059
rect 14645 14019 14703 14025
rect 2590 13948 2596 14000
rect 2648 13988 2654 14000
rect 2777 13991 2835 13997
rect 2777 13988 2789 13991
rect 2648 13960 2789 13988
rect 2648 13948 2654 13960
rect 2777 13957 2789 13960
rect 2823 13957 2835 13991
rect 2777 13951 2835 13957
rect 2958 13948 2964 14000
rect 3016 13988 3022 14000
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 3016 13960 3249 13988
rect 3016 13948 3022 13960
rect 3237 13957 3249 13960
rect 3283 13957 3295 13991
rect 3237 13951 3295 13957
rect 3881 13923 3939 13929
rect 3881 13920 3893 13923
rect 3160 13892 3893 13920
rect 3160 13861 3188 13892
rect 3881 13889 3893 13892
rect 3927 13920 3939 13923
rect 9122 13920 9128 13932
rect 3927 13892 9128 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13821 3203 13855
rect 6270 13852 6276 13864
rect 6231 13824 6276 13852
rect 3145 13815 3203 13821
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10042 13852 10048 13864
rect 9815 13824 10048 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10042 13812 10048 13824
rect 10100 13812 10106 13864
rect 13078 13812 13084 13864
rect 13136 13852 13142 13864
rect 14461 13855 14519 13861
rect 14461 13852 14473 13855
rect 13136 13824 14473 13852
rect 13136 13812 13142 13824
rect 14461 13821 14473 13824
rect 14507 13852 14519 13855
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 14507 13824 15025 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 15013 13821 15025 13824
rect 15059 13821 15071 13855
rect 15013 13815 15071 13821
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 7156 13688 7205 13716
rect 7156 13676 7162 13688
rect 7193 13685 7205 13688
rect 7239 13716 7251 13719
rect 9214 13716 9220 13728
rect 7239 13688 9220 13716
rect 7239 13685 7251 13688
rect 7193 13679 7251 13685
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 5534 13444 5540 13456
rect 4356 13416 5540 13444
rect 4356 13385 4384 13416
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13345 4399 13379
rect 4597 13379 4655 13385
rect 4597 13376 4609 13379
rect 4341 13339 4399 13345
rect 4448 13348 4609 13376
rect 3970 13268 3976 13320
rect 4028 13308 4034 13320
rect 4448 13308 4476 13348
rect 4597 13345 4609 13348
rect 4643 13345 4655 13379
rect 4597 13339 4655 13345
rect 4028 13280 4476 13308
rect 4028 13268 4034 13280
rect 5721 13175 5779 13181
rect 5721 13141 5733 13175
rect 5767 13172 5779 13175
rect 6914 13172 6920 13184
rect 5767 13144 6920 13172
rect 5767 13141 5779 13144
rect 5721 13135 5779 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7742 13172 7748 13184
rect 7703 13144 7748 13172
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 3970 12928 3976 12980
rect 4028 12968 4034 12980
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 4028 12940 4629 12968
rect 4028 12928 4034 12940
rect 4617 12937 4629 12940
rect 4663 12937 4675 12971
rect 4617 12931 4675 12937
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5534 12968 5540 12980
rect 5123 12940 5540 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7466 12832 7472 12844
rect 7248 12804 7472 12832
rect 7248 12792 7254 12804
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 7699 12804 8156 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 7374 12764 7380 12776
rect 7287 12736 7380 12764
rect 7374 12724 7380 12736
rect 7432 12764 7438 12776
rect 7742 12764 7748 12776
rect 7432 12736 7748 12764
rect 7432 12724 7438 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7742 12628 7748 12640
rect 7156 12600 7748 12628
rect 7156 12588 7162 12600
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 8128 12637 8156 12804
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8662 12628 8668 12640
rect 8159 12600 8668 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 13722 12628 13728 12640
rect 9180 12600 13728 12628
rect 9180 12588 9186 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 6730 12424 6736 12436
rect 6420 12396 6736 12424
rect 6420 12384 6426 12396
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 4522 12316 4528 12368
rect 4580 12356 4586 12368
rect 4706 12356 4712 12368
rect 4580 12328 4712 12356
rect 4580 12316 4586 12328
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 6086 12288 6092 12300
rect 6047 12260 6092 12288
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6270 12044 6276 12096
rect 6328 12084 6334 12096
rect 6822 12084 6828 12096
rect 6328 12056 6828 12084
rect 6328 12044 6334 12056
rect 6822 12044 6828 12056
rect 6880 12084 6886 12096
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 6880 12056 7389 12084
rect 6880 12044 6886 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 8076 12056 8125 12084
rect 8076 12044 8082 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 7561 11883 7619 11889
rect 7561 11880 7573 11883
rect 5592 11852 7573 11880
rect 5592 11840 5598 11852
rect 7561 11849 7573 11852
rect 7607 11849 7619 11883
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 7561 11843 7619 11849
rect 7576 11744 7604 11843
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 7745 11747 7803 11753
rect 7745 11744 7757 11747
rect 7576 11716 7757 11744
rect 7745 11713 7757 11716
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 8018 11685 8024 11688
rect 8012 11676 8024 11685
rect 7979 11648 8024 11676
rect 8012 11639 8024 11648
rect 8018 11636 8024 11639
rect 8076 11636 8082 11688
rect 6086 11568 6092 11620
rect 6144 11568 6150 11620
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 8110 11608 8116 11620
rect 7708 11580 8116 11608
rect 7708 11568 7714 11580
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10134 11608 10140 11620
rect 9916 11580 10140 11608
rect 9916 11568 9922 11580
rect 10134 11568 10140 11580
rect 10192 11568 10198 11620
rect 6104 11540 6132 11568
rect 6181 11543 6239 11549
rect 6181 11540 6193 11543
rect 6104 11512 6193 11540
rect 6181 11509 6193 11512
rect 6227 11540 6239 11543
rect 11146 11540 11152 11552
rect 6227 11512 11152 11540
rect 6227 11509 6239 11512
rect 6181 11503 6239 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 6880 11308 7113 11336
rect 6880 11296 6886 11308
rect 7101 11305 7113 11308
rect 7147 11305 7159 11339
rect 8662 11336 8668 11348
rect 8623 11308 8668 11336
rect 7101 11299 7159 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 10137 11339 10195 11345
rect 10137 11336 10149 11339
rect 9732 11308 10149 11336
rect 9732 11296 9738 11308
rect 10137 11305 10149 11308
rect 10183 11336 10195 11339
rect 10410 11336 10416 11348
rect 10183 11308 10416 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 7650 11268 7656 11280
rect 7300 11240 7656 11268
rect 2958 11209 2964 11212
rect 2936 11203 2964 11209
rect 2936 11169 2948 11203
rect 2936 11163 2964 11169
rect 2958 11160 2964 11163
rect 3016 11160 3022 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 5592 11172 6101 11200
rect 5592 11160 5598 11172
rect 6089 11169 6101 11172
rect 6135 11200 6147 11203
rect 6638 11200 6644 11212
rect 6135 11172 6644 11200
rect 6135 11169 6147 11172
rect 6089 11163 6147 11169
rect 6638 11160 6644 11172
rect 6696 11200 6702 11212
rect 7300 11209 7328 11240
rect 7650 11228 7656 11240
rect 7708 11268 7714 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 7708 11240 8953 11268
rect 7708 11228 7714 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 8941 11231 8999 11237
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 6696 11172 6745 11200
rect 6696 11160 6702 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 6733 11163 6791 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7541 11203 7599 11209
rect 7541 11200 7553 11203
rect 7285 11163 7343 11169
rect 7392 11172 7553 11200
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 6178 11132 6184 11144
rect 5868 11104 6184 11132
rect 5868 11092 5874 11104
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11132 6423 11135
rect 6914 11132 6920 11144
rect 6411 11104 6920 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 6914 11092 6920 11104
rect 6972 11132 6978 11144
rect 7392 11132 7420 11172
rect 7541 11169 7553 11172
rect 7587 11169 7599 11203
rect 7541 11163 7599 11169
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11200 10103 11203
rect 10410 11200 10416 11212
rect 10091 11172 10416 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 6972 11104 7420 11132
rect 6972 11092 6978 11104
rect 7300 11076 7328 11104
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 8720 11104 10241 11132
rect 8720 11092 8726 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 5721 11067 5779 11073
rect 5721 11033 5733 11067
rect 5767 11064 5779 11067
rect 7190 11064 7196 11076
rect 5767 11036 7196 11064
rect 5767 11033 5779 11036
rect 5721 11027 5779 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7282 11024 7288 11076
rect 7340 11024 7346 11076
rect 9677 11067 9735 11073
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 9766 11064 9772 11076
rect 9723 11036 9772 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 3007 10999 3065 11005
rect 3007 10965 3019 10999
rect 3053 10996 3065 10999
rect 3326 10996 3332 11008
rect 3053 10968 3332 10996
rect 3053 10965 3065 10968
rect 3007 10959 3065 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 10226 10996 10232 11008
rect 9916 10968 10232 10996
rect 9916 10956 9922 10968
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 10689 10999 10747 11005
rect 10689 10996 10701 10999
rect 10652 10968 10701 10996
rect 10652 10956 10658 10968
rect 10689 10965 10701 10968
rect 10735 10965 10747 10999
rect 10689 10959 10747 10965
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 2958 10792 2964 10804
rect 2919 10764 2964 10792
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3384 10764 3525 10792
rect 3384 10752 3390 10764
rect 3513 10761 3525 10764
rect 3559 10792 3571 10795
rect 3878 10792 3884 10804
rect 3559 10764 3884 10792
rect 3559 10761 3571 10764
rect 3513 10755 3571 10761
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 6178 10792 6184 10804
rect 6091 10764 6184 10792
rect 6178 10752 6184 10764
rect 6236 10792 6242 10804
rect 9674 10792 9680 10804
rect 6236 10764 8616 10792
rect 9635 10764 9680 10792
rect 6236 10752 6242 10764
rect 8588 10736 8616 10764
rect 9674 10752 9680 10764
rect 9732 10792 9738 10804
rect 9858 10792 9864 10804
rect 9732 10764 9864 10792
rect 9732 10752 9738 10764
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 6457 10727 6515 10733
rect 6457 10693 6469 10727
rect 6503 10724 6515 10727
rect 6503 10696 7604 10724
rect 6503 10693 6515 10696
rect 6457 10687 6515 10693
rect 3786 10656 3792 10668
rect 3747 10628 3792 10656
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 6822 10588 6828 10600
rect 6687 10560 6828 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7576 10597 7604 10696
rect 8570 10684 8576 10736
rect 8628 10684 8634 10736
rect 9398 10684 9404 10736
rect 9456 10724 9462 10736
rect 9769 10727 9827 10733
rect 9769 10724 9781 10727
rect 9456 10696 9781 10724
rect 9456 10684 9462 10696
rect 9769 10693 9781 10696
rect 9815 10693 9827 10727
rect 11149 10727 11207 10733
rect 11149 10724 11161 10727
rect 9769 10687 9827 10693
rect 10336 10696 11161 10724
rect 10336 10665 10364 10696
rect 11149 10693 11161 10696
rect 11195 10693 11207 10727
rect 11149 10687 11207 10693
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 8772 10628 10333 10656
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 7650 10588 7656 10600
rect 7607 10560 7656 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 3878 10480 3884 10532
rect 3936 10520 3942 10532
rect 4798 10520 4804 10532
rect 3936 10492 3981 10520
rect 4759 10492 4804 10520
rect 3936 10480 3942 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10520 5871 10523
rect 7101 10523 7159 10529
rect 5859 10492 7052 10520
rect 5859 10489 5871 10492
rect 5813 10483 5871 10489
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 2958 10452 2964 10464
rect 1636 10424 2964 10452
rect 1636 10412 1642 10424
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 7024 10452 7052 10492
rect 7101 10489 7113 10523
rect 7147 10520 7159 10523
rect 7828 10523 7886 10529
rect 7828 10520 7840 10523
rect 7147 10492 7840 10520
rect 7147 10489 7159 10492
rect 7101 10483 7159 10489
rect 7828 10489 7840 10492
rect 7874 10520 7886 10523
rect 8662 10520 8668 10532
rect 7874 10492 8668 10520
rect 7874 10489 7886 10492
rect 7828 10483 7886 10489
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 7282 10452 7288 10464
rect 7024 10424 7288 10452
rect 7282 10412 7288 10424
rect 7340 10452 7346 10464
rect 7466 10452 7472 10464
rect 7340 10424 7472 10452
rect 7340 10412 7346 10424
rect 7466 10412 7472 10424
rect 7524 10452 7530 10464
rect 8772 10452 8800 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 10468 10628 11345 10656
rect 10468 10616 10474 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 10428 10588 10456 10616
rect 9355 10560 10456 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 10137 10523 10195 10529
rect 10137 10489 10149 10523
rect 10183 10520 10195 10523
rect 10594 10520 10600 10532
rect 10183 10492 10600 10520
rect 10183 10489 10195 10492
rect 10137 10483 10195 10489
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 8938 10452 8944 10464
rect 7524 10424 8800 10452
rect 8899 10424 8944 10452
rect 7524 10412 7530 10424
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10410 10452 10416 10464
rect 10284 10424 10416 10452
rect 10284 10412 10290 10424
rect 10410 10412 10416 10424
rect 10468 10452 10474 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10468 10424 10793 10452
rect 10468 10412 10474 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 7193 10251 7251 10257
rect 7193 10217 7205 10251
rect 7239 10248 7251 10251
rect 7282 10248 7288 10260
rect 7239 10220 7288 10248
rect 7239 10217 7251 10220
rect 7193 10211 7251 10217
rect 7282 10208 7288 10220
rect 7340 10248 7346 10260
rect 7650 10248 7656 10260
rect 7340 10220 7656 10248
rect 7340 10208 7346 10220
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8076 10220 8677 10248
rect 8076 10208 8082 10220
rect 8665 10217 8677 10220
rect 8711 10217 8723 10251
rect 8665 10211 8723 10217
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8812 10220 8953 10248
rect 8812 10208 8818 10220
rect 8941 10217 8953 10220
rect 8987 10248 8999 10251
rect 9122 10248 9128 10260
rect 8987 10220 9128 10248
rect 8987 10217 8999 10220
rect 8941 10211 8999 10217
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9398 10248 9404 10260
rect 9359 10220 9404 10248
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10318 10248 10324 10260
rect 10183 10220 10324 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 1578 10180 1584 10192
rect 1539 10152 1584 10180
rect 1578 10140 1584 10152
rect 1636 10140 1642 10192
rect 2501 10183 2559 10189
rect 2501 10149 2513 10183
rect 2547 10180 2559 10183
rect 2774 10180 2780 10192
rect 2547 10152 2780 10180
rect 2547 10149 2559 10152
rect 2501 10143 2559 10149
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 4798 10140 4804 10192
rect 4856 10180 4862 10192
rect 13078 10180 13084 10192
rect 4856 10152 13084 10180
rect 4856 10140 4862 10152
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 7282 10112 7288 10124
rect 6135 10084 6868 10112
rect 7243 10084 7288 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 1946 10044 1952 10056
rect 1535 10016 1952 10044
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5868 10016 6193 10044
rect 5868 10004 5874 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6362 10044 6368 10056
rect 6323 10016 6368 10044
rect 6181 10007 6239 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 5718 9908 5724 9920
rect 5679 9880 5724 9908
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 6840 9917 6868 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7552 10115 7610 10121
rect 7552 10081 7564 10115
rect 7598 10112 7610 10115
rect 8938 10112 8944 10124
rect 7598 10084 8944 10112
rect 7598 10081 7610 10084
rect 7552 10075 7610 10081
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 10042 10112 10048 10124
rect 10003 10084 10048 10112
rect 10042 10072 10048 10084
rect 10100 10072 10106 10124
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10044 10287 10047
rect 10689 10047 10747 10053
rect 10689 10044 10701 10047
rect 10275 10016 10701 10044
rect 10275 10013 10287 10016
rect 10229 10007 10287 10013
rect 10689 10013 10701 10016
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 9122 9936 9128 9988
rect 9180 9976 9186 9988
rect 10244 9976 10272 10007
rect 9180 9948 10272 9976
rect 9180 9936 9186 9948
rect 6825 9911 6883 9917
rect 6825 9877 6837 9911
rect 6871 9908 6883 9911
rect 6914 9908 6920 9920
rect 6871 9880 6920 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 9674 9908 9680 9920
rect 9635 9880 9680 9908
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 10226 9868 10232 9920
rect 10284 9908 10290 9920
rect 10594 9908 10600 9920
rect 10284 9880 10600 9908
rect 10284 9868 10290 9880
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 5166 9704 5172 9716
rect 4396 9676 5172 9704
rect 4396 9664 4402 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 6181 9707 6239 9713
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 6362 9704 6368 9716
rect 6227 9676 6368 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 6362 9664 6368 9676
rect 6420 9704 6426 9716
rect 8018 9704 8024 9716
rect 6420 9676 8024 9704
rect 6420 9664 6426 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 10376 9676 10425 9704
rect 10376 9664 10382 9676
rect 10413 9673 10425 9676
rect 10459 9673 10471 9707
rect 10413 9667 10471 9673
rect 6917 9639 6975 9645
rect 6917 9605 6929 9639
rect 6963 9636 6975 9639
rect 7374 9636 7380 9648
rect 6963 9608 7380 9636
rect 6963 9605 6975 9608
rect 6917 9599 6975 9605
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 7524 9608 8309 9636
rect 7524 9596 7530 9608
rect 7576 9577 7604 9608
rect 8297 9605 8309 9608
rect 8343 9605 8355 9639
rect 9214 9636 9220 9648
rect 8297 9599 8355 9605
rect 8864 9608 9220 9636
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 7607 9540 7641 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 6638 9500 6644 9512
rect 6551 9472 6644 9500
rect 6638 9460 6644 9472
rect 6696 9500 6702 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 6696 9472 7297 9500
rect 6696 9460 6702 9472
rect 7285 9469 7297 9472
rect 7331 9500 7343 9503
rect 8754 9500 8760 9512
rect 7331 9472 8760 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 8864 9509 8892 9608
rect 9214 9596 9220 9608
rect 9272 9636 9278 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 9272 9608 9505 9636
rect 9272 9596 9278 9608
rect 9493 9605 9505 9608
rect 9539 9636 9551 9639
rect 12894 9636 12900 9648
rect 9539 9608 12900 9636
rect 9539 9605 9551 9608
rect 9493 9599 9551 9605
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 9122 9568 9128 9580
rect 9083 9540 9128 9568
rect 9122 9528 9128 9540
rect 9180 9568 9186 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 9180 9540 10793 9568
rect 9180 9528 9186 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9398 9500 9404 9512
rect 8987 9472 9404 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 7377 9435 7435 9441
rect 7377 9432 7389 9435
rect 4764 9404 7389 9432
rect 4764 9392 4770 9404
rect 7377 9401 7389 9404
rect 7423 9432 7435 9435
rect 8021 9435 8079 9441
rect 8021 9432 8033 9435
rect 7423 9404 8033 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 8021 9401 8033 9404
rect 8067 9432 8079 9435
rect 9490 9432 9496 9444
rect 8067 9404 9496 9432
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1946 9364 1952 9376
rect 1907 9336 1952 9364
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 5810 9364 5816 9376
rect 5771 9336 5816 9364
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 10042 9364 10048 9376
rect 10003 9336 10048 9364
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 5868 9132 7297 9160
rect 5868 9120 5874 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7285 9123 7343 9129
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7653 9163 7711 9169
rect 7653 9160 7665 9163
rect 7432 9132 7665 9160
rect 7432 9120 7438 9132
rect 7653 9129 7665 9132
rect 7699 9160 7711 9163
rect 8478 9160 8484 9172
rect 7699 9132 8484 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 9674 9160 9680 9172
rect 8803 9132 9680 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 7006 9052 7012 9104
rect 7064 9092 7070 9104
rect 7745 9095 7803 9101
rect 7745 9092 7757 9095
rect 7064 9064 7757 9092
rect 7064 9052 7070 9064
rect 7745 9061 7757 9064
rect 7791 9092 7803 9095
rect 8018 9092 8024 9104
rect 7791 9064 8024 9092
rect 7791 9061 7803 9064
rect 7745 9055 7803 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 8389 9095 8447 9101
rect 8389 9061 8401 9095
rect 8435 9092 8447 9095
rect 8938 9092 8944 9104
rect 8435 9064 8944 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7282 9024 7288 9036
rect 7239 8996 7288 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 7892 8928 7941 8956
rect 7892 8916 7898 8928
rect 7929 8925 7941 8928
rect 7975 8956 7987 8959
rect 8404 8956 8432 9055
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 12437 9027 12495 9033
rect 12437 8993 12449 9027
rect 12483 9024 12495 9027
rect 12710 9024 12716 9036
rect 12483 8996 12716 9024
rect 12483 8993 12495 8996
rect 12437 8987 12495 8993
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 7975 8928 8432 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 11204 8928 12633 8956
rect 11204 8916 11210 8928
rect 12621 8925 12633 8928
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 7834 8616 7840 8628
rect 7791 8588 7840 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 6972 8520 8217 8548
rect 6972 8508 6978 8520
rect 8205 8517 8217 8520
rect 8251 8517 8263 8551
rect 8205 8511 8263 8517
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 8938 8480 8944 8492
rect 8895 8452 8944 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 8938 8440 8944 8452
rect 8996 8480 9002 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 8996 8452 9229 8480
rect 8996 8440 9002 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 9674 8412 9680 8424
rect 8711 8384 9680 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 8570 8344 8576 8356
rect 8483 8316 8576 8344
rect 8570 8304 8576 8316
rect 8628 8344 8634 8356
rect 9766 8344 9772 8356
rect 8628 8316 9772 8344
rect 8628 8304 8634 8316
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 12710 8344 12716 8356
rect 12671 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 9122 8276 9128 8288
rect 8904 8248 9128 8276
rect 8904 8236 8910 8248
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 8570 8072 8576 8084
rect 8531 8044 8576 8072
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 4157 7531 4215 7537
rect 4157 7497 4169 7531
rect 4203 7528 4215 7531
rect 5718 7528 5724 7540
rect 4203 7500 5724 7528
rect 4203 7497 4215 7500
rect 4157 7491 4215 7497
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 4172 7324 4200 7491
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 3375 7296 4200 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3605 7259 3663 7265
rect 3605 7256 3617 7259
rect 3016 7228 3617 7256
rect 3016 7216 3022 7228
rect 3605 7225 3617 7228
rect 3651 7225 3663 7259
rect 3605 7219 3663 7225
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 5074 6440 5080 6452
rect 5035 6412 5080 6440
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 9858 6440 9864 6452
rect 9815 6412 9864 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 7006 6332 7012 6384
rect 7064 6372 7070 6384
rect 9309 6375 9367 6381
rect 9309 6372 9321 6375
rect 7064 6344 9321 6372
rect 7064 6332 7070 6344
rect 9309 6341 9321 6344
rect 9355 6341 9367 6375
rect 9309 6335 9367 6341
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6236 4951 6239
rect 7469 6239 7527 6245
rect 4939 6208 5580 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 5552 6109 5580 6208
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9784 6236 9812 6403
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10042 6332 10048 6384
rect 10100 6372 10106 6384
rect 15470 6372 15476 6384
rect 10100 6344 15476 6372
rect 10100 6332 10106 6344
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 9171 6208 9812 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 7484 6168 7512 6199
rect 8113 6171 8171 6177
rect 8113 6168 8125 6171
rect 7484 6140 8125 6168
rect 8113 6137 8125 6140
rect 8159 6168 8171 6171
rect 10318 6168 10324 6180
rect 8159 6140 10324 6168
rect 8159 6137 8171 6140
rect 8113 6131 8171 6137
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 5537 6103 5595 6109
rect 5537 6069 5549 6103
rect 5583 6100 5595 6103
rect 6362 6100 6368 6112
rect 5583 6072 6368 6100
rect 5583 6069 5595 6072
rect 5537 6063 5595 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 7650 6100 7656 6112
rect 7611 6072 7656 6100
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 3200 5868 7205 5896
rect 3200 5856 3206 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 8260 5868 9873 5896
rect 8260 5856 8266 5868
rect 9861 5865 9873 5868
rect 9907 5865 9919 5899
rect 9861 5859 9919 5865
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 10744 5868 12173 5896
rect 10744 5856 10750 5868
rect 12161 5865 12173 5868
rect 12207 5865 12219 5899
rect 12161 5859 12219 5865
rect 5534 5828 5540 5840
rect 4172 5800 5540 5828
rect 4172 5772 4200 5800
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4154 5760 4160 5772
rect 4111 5732 4160 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5760 5227 5763
rect 6638 5760 6644 5772
rect 5215 5732 6644 5760
rect 5215 5729 5227 5732
rect 5169 5723 5227 5729
rect 5552 5704 5580 5732
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7834 5760 7840 5772
rect 7055 5732 7840 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5760 8171 5763
rect 9030 5760 9036 5772
rect 8159 5732 9036 5760
rect 8159 5729 8171 5732
rect 8113 5723 8171 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 9766 5760 9772 5772
rect 9723 5732 9772 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11238 5760 11244 5772
rect 10827 5732 11244 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 11977 5763 12035 5769
rect 11977 5729 11989 5763
rect 12023 5760 12035 5763
rect 12250 5760 12256 5772
rect 12023 5732 12256 5760
rect 12023 5729 12035 5732
rect 11977 5723 12035 5729
rect 12250 5720 12256 5732
rect 12308 5720 12314 5772
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 10226 5692 10232 5704
rect 7668 5664 10232 5692
rect 7668 5624 7696 5664
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10686 5652 10692 5704
rect 10744 5692 10750 5704
rect 12802 5692 12808 5704
rect 10744 5664 12808 5692
rect 10744 5652 10750 5664
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 4632 5596 7696 5624
rect 4246 5556 4252 5568
rect 4207 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4522 5516 4528 5568
rect 4580 5556 4586 5568
rect 4632 5565 4660 5596
rect 7742 5584 7748 5636
rect 7800 5624 7806 5636
rect 10965 5627 11023 5633
rect 10965 5624 10977 5627
rect 7800 5596 10977 5624
rect 7800 5584 7806 5596
rect 10965 5593 10977 5596
rect 11011 5593 11023 5627
rect 10965 5587 11023 5593
rect 4617 5559 4675 5565
rect 4617 5556 4629 5559
rect 4580 5528 4629 5556
rect 4580 5516 4586 5528
rect 4617 5525 4629 5528
rect 4663 5525 4675 5559
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 4617 5519 4675 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 8297 5559 8355 5565
rect 8297 5556 8309 5559
rect 7340 5528 8309 5556
rect 7340 5516 7346 5528
rect 8297 5525 8309 5528
rect 8343 5525 8355 5559
rect 8297 5519 8355 5525
rect 9125 5559 9183 5565
rect 9125 5525 9137 5559
rect 9171 5556 9183 5559
rect 9306 5556 9312 5568
rect 9171 5528 9312 5556
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 4154 5352 4160 5364
rect 4115 5324 4160 5352
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5261 5355 5319 5361
rect 5261 5321 5273 5355
rect 5307 5352 5319 5355
rect 5534 5352 5540 5364
rect 5307 5324 5540 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5684 5324 5825 5352
rect 5684 5312 5690 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 8168 5324 12633 5352
rect 8168 5312 8174 5324
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 12621 5315 12679 5321
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 7009 5287 7067 5293
rect 7009 5284 7021 5287
rect 2740 5256 7021 5284
rect 2740 5244 2746 5256
rect 7009 5253 7021 5256
rect 7055 5253 7067 5287
rect 7834 5284 7840 5296
rect 7747 5256 7840 5284
rect 7009 5247 7067 5253
rect 7834 5244 7840 5256
rect 7892 5284 7898 5296
rect 10502 5284 10508 5296
rect 7892 5256 10508 5284
rect 7892 5244 7898 5256
rect 10502 5244 10508 5256
rect 10560 5244 10566 5296
rect 6273 5219 6331 5225
rect 6273 5216 6285 5219
rect 5644 5188 6285 5216
rect 4522 5148 4528 5160
rect 4483 5120 4528 5148
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5644 5157 5672 5188
rect 6273 5185 6285 5188
rect 6319 5216 6331 5219
rect 9858 5216 9864 5228
rect 6319 5188 9864 5216
rect 6319 5185 6331 5188
rect 6273 5179 6331 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5216 10839 5219
rect 11790 5216 11796 5228
rect 10827 5188 11796 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5117 5687 5151
rect 5629 5111 5687 5117
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7466 5148 7472 5160
rect 6871 5120 7472 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 9033 5151 9091 5157
rect 7975 5120 8616 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 4062 5040 4068 5092
rect 4120 5080 4126 5092
rect 4120 5052 8156 5080
rect 4120 5040 4126 5052
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 7466 5012 7472 5024
rect 7427 4984 7472 5012
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 8128 5021 8156 5052
rect 8588 5021 8616 5120
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 9306 5148 9312 5160
rect 9079 5120 9312 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 10137 5151 10195 5157
rect 10137 5117 10149 5151
rect 10183 5148 10195 5151
rect 10796 5148 10824 5179
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 10183 5120 10824 5148
rect 11241 5151 11299 5157
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 11241 5117 11253 5151
rect 11287 5117 11299 5151
rect 11241 5111 11299 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12483 5120 13124 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 11256 5080 11284 5111
rect 11885 5083 11943 5089
rect 11885 5080 11897 5083
rect 11256 5052 11897 5080
rect 11885 5049 11897 5052
rect 11931 5080 11943 5083
rect 12986 5080 12992 5092
rect 11931 5052 12992 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 8573 5015 8631 5021
rect 8573 4981 8585 5015
rect 8619 5012 8631 5015
rect 8754 5012 8760 5024
rect 8619 4984 8760 5012
rect 8619 4981 8631 4984
rect 8573 4975 8631 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 8941 5015 8999 5021
rect 8941 4981 8953 5015
rect 8987 5012 8999 5015
rect 9030 5012 9036 5024
rect 8987 4984 9036 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 9214 5012 9220 5024
rect 9175 4984 9220 5012
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9766 5012 9772 5024
rect 9727 4984 9772 5012
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 10318 5012 10324 5024
rect 10279 4984 10324 5012
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11238 5012 11244 5024
rect 11195 4984 11244 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 11425 5015 11483 5021
rect 11425 5012 11437 5015
rect 11388 4984 11437 5012
rect 11388 4972 11394 4984
rect 11425 4981 11437 4984
rect 11471 4981 11483 5015
rect 12250 5012 12256 5024
rect 12211 4984 12256 5012
rect 11425 4975 11483 4981
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 13096 5021 13124 5120
rect 13081 5015 13139 5021
rect 13081 4981 13093 5015
rect 13127 5012 13139 5015
rect 15930 5012 15936 5024
rect 13127 4984 15936 5012
rect 13127 4981 13139 4984
rect 13081 4975 13139 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 8021 4811 8079 4817
rect 8021 4808 8033 4811
rect 4028 4780 8033 4808
rect 4028 4768 4034 4780
rect 8021 4777 8033 4780
rect 8067 4777 8079 4811
rect 8021 4771 8079 4777
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 10008 4780 10149 4808
rect 10008 4768 10014 4780
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 12618 4808 12624 4820
rect 12579 4780 12624 4808
rect 10137 4771 10195 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 9214 4740 9220 4752
rect 5224 4712 9220 4740
rect 5224 4700 5230 4712
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 13814 4740 13820 4752
rect 10836 4712 13820 4740
rect 10836 4700 10842 4712
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 4890 4672 4896 4684
rect 4847 4644 4896 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4672 5963 4675
rect 5994 4672 6000 4684
rect 5951 4644 6000 4672
rect 5951 4641 5963 4644
rect 5905 4635 5963 4641
rect 5994 4632 6000 4644
rect 6052 4672 6058 4684
rect 6454 4672 6460 4684
rect 6052 4644 6460 4672
rect 6052 4632 6058 4644
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4672 7895 4675
rect 8662 4672 8668 4684
rect 7883 4644 8668 4672
rect 7883 4641 7895 4644
rect 7837 4635 7895 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10042 4672 10048 4684
rect 9999 4644 10048 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 11057 4675 11115 4681
rect 11057 4641 11069 4675
rect 11103 4672 11115 4675
rect 11422 4672 11428 4684
rect 11103 4644 11428 4672
rect 11103 4641 11115 4644
rect 11057 4635 11115 4641
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4672 12495 4675
rect 12710 4672 12716 4684
rect 12483 4644 12716 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 13630 4672 13636 4684
rect 13587 4644 13636 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 11330 4604 11336 4616
rect 6788 4576 11336 4604
rect 6788 4564 6794 4576
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 10318 4536 10324 4548
rect 5500 4508 10324 4536
rect 5500 4496 5506 4508
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 16206 4536 16212 4548
rect 12492 4508 16212 4536
rect 12492 4496 12498 4508
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 4982 4468 4988 4480
rect 4943 4440 4988 4468
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 6086 4468 6092 4480
rect 6047 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10594 4468 10600 4480
rect 10008 4440 10600 4468
rect 10008 4428 10014 4440
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 11241 4471 11299 4477
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 11330 4468 11336 4480
rect 11287 4440 11336 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 13722 4468 13728 4480
rect 13683 4440 13728 4468
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 4890 4264 4896 4276
rect 4851 4236 4896 4264
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5994 4264 6000 4276
rect 5955 4236 6000 4264
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 7469 4267 7527 4273
rect 7469 4233 7481 4267
rect 7515 4264 7527 4267
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7515 4236 7573 4264
rect 7515 4233 7527 4236
rect 7469 4227 7527 4233
rect 7561 4233 7573 4236
rect 7607 4264 7619 4267
rect 10134 4264 10140 4276
rect 7607 4236 10140 4264
rect 7607 4233 7619 4236
rect 7561 4227 7619 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10778 4264 10784 4276
rect 10739 4236 10784 4264
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 11149 4267 11207 4273
rect 11149 4233 11161 4267
rect 11195 4264 11207 4267
rect 11422 4264 11428 4276
rect 11195 4236 11428 4264
rect 11195 4233 11207 4236
rect 11149 4227 11207 4233
rect 11422 4224 11428 4236
rect 11480 4224 11486 4276
rect 11701 4267 11759 4273
rect 11701 4233 11713 4267
rect 11747 4264 11759 4267
rect 11885 4267 11943 4273
rect 11885 4264 11897 4267
rect 11747 4236 11897 4264
rect 11747 4233 11759 4236
rect 11701 4227 11759 4233
rect 11885 4233 11897 4236
rect 11931 4264 11943 4267
rect 13630 4264 13636 4276
rect 11931 4236 12756 4264
rect 13591 4236 13636 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 7760 4168 8064 4196
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3200 4100 6316 4128
rect 3200 4088 3206 4100
rect 1394 3952 1400 4004
rect 1452 3992 1458 4004
rect 6086 3992 6092 4004
rect 1452 3964 6092 3992
rect 1452 3952 1458 3964
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 6288 3992 6316 4100
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 7760 4128 7788 4168
rect 6420 4100 7788 4128
rect 6420 4088 6426 4100
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8036 4128 8064 4168
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 10594 4196 10600 4208
rect 8812 4168 10600 4196
rect 8812 4156 8818 4168
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 12728 4196 12756 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 15102 4196 15108 4208
rect 12728 4168 15108 4196
rect 15102 4156 15108 4168
rect 15160 4156 15166 4208
rect 8478 4128 8484 4140
rect 7892 4100 7937 4128
rect 8036 4100 8484 4128
rect 7892 4088 7898 4100
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9048 4100 9689 4128
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 6871 4032 7573 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 7852 4060 7880 4088
rect 9048 4069 9076 4100
rect 9677 4097 9689 4100
rect 9723 4128 9735 4131
rect 10686 4128 10692 4140
rect 9723 4100 10692 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 14642 4128 14648 4140
rect 13044 4100 14648 4128
rect 13044 4088 13050 4100
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 7935 4063 7993 4069
rect 7935 4060 7947 4063
rect 7852 4032 7947 4060
rect 7561 4023 7619 4029
rect 7935 4029 7947 4032
rect 7981 4029 7993 4063
rect 7935 4023 7993 4029
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4060 10195 4063
rect 10778 4060 10784 4072
rect 10183 4032 10784 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11287 4032 11713 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4060 12311 4063
rect 12434 4060 12440 4072
rect 12299 4032 12440 4060
rect 12299 4029 12311 4032
rect 12253 4023 12311 4029
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 6288 3964 8156 3992
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 8128 3933 8156 3964
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 8260 3964 12664 3992
rect 8260 3952 8266 3964
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 2372 3896 7021 3924
rect 2372 3884 2378 3896
rect 7009 3893 7021 3896
rect 7055 3893 7067 3927
rect 7009 3887 7067 3893
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3893 8171 3927
rect 8570 3924 8576 3936
rect 8531 3896 8576 3924
rect 8113 3887 8171 3893
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12636 3933 12664 3964
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3893 12679 3927
rect 12621 3887 12679 3893
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12768 3896 13093 3924
rect 12768 3884 12774 3896
rect 13081 3893 13093 3896
rect 13127 3924 13139 3927
rect 16758 3924 16764 3936
rect 13127 3896 16764 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 6270 3680 6276 3732
rect 6328 3720 6334 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 6328 3692 10425 3720
rect 6328 3680 6334 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 16298 3720 16304 3732
rect 12308 3692 16304 3720
rect 12308 3680 12314 3692
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 4798 3612 4804 3664
rect 4856 3652 4862 3664
rect 9214 3652 9220 3664
rect 4856 3624 9220 3652
rect 4856 3612 4862 3624
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 9306 3612 9312 3664
rect 9364 3652 9370 3664
rect 11054 3652 11060 3664
rect 9364 3624 11060 3652
rect 9364 3612 9370 3624
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 6822 3584 6828 3596
rect 6783 3556 6828 3584
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 8110 3584 8116 3596
rect 7616 3556 8116 3584
rect 7616 3544 7622 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 9030 3584 9036 3596
rect 8536 3556 9036 3584
rect 8536 3544 8542 3556
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 10226 3584 10232 3596
rect 10187 3556 10232 3584
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 11514 3544 11520 3596
rect 11572 3593 11578 3596
rect 11572 3584 11581 3593
rect 11572 3556 11617 3584
rect 11572 3547 11581 3556
rect 11572 3544 11578 3547
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 10318 3516 10324 3528
rect 5316 3488 10324 3516
rect 5316 3476 5322 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 15010 3516 15016 3528
rect 11296 3488 15016 3516
rect 11296 3476 11302 3488
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 8297 3451 8355 3457
rect 8297 3448 8309 3451
rect 4028 3420 8309 3448
rect 4028 3408 4034 3420
rect 8297 3417 8309 3420
rect 8343 3417 8355 3451
rect 8297 3411 8355 3417
rect 8570 3408 8576 3460
rect 8628 3448 8634 3460
rect 12066 3448 12072 3460
rect 8628 3420 12072 3448
rect 8628 3408 8634 3420
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 2682 3340 2688 3392
rect 2740 3380 2746 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 2740 3352 7021 3380
rect 2740 3340 2746 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 11701 3383 11759 3389
rect 11701 3380 11713 3383
rect 7432 3352 11713 3380
rect 7432 3340 7438 3352
rect 11701 3349 11713 3352
rect 11747 3349 11759 3383
rect 11701 3343 11759 3349
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 13170 3380 13176 3392
rect 11848 3352 13176 3380
rect 11848 3340 11854 3352
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 7650 3176 7656 3188
rect 4488 3148 7656 3176
rect 4488 3136 4494 3148
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 8110 3176 8116 3188
rect 8071 3148 8116 3176
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 9122 3176 9128 3188
rect 8720 3148 9128 3176
rect 8720 3136 8726 3148
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 11609 3179 11667 3185
rect 9824 3148 11560 3176
rect 9824 3136 9830 3148
rect 3786 3068 3792 3120
rect 3844 3108 3850 3120
rect 3844 3080 5488 3108
rect 3844 3068 3850 3080
rect 1026 3000 1032 3052
rect 1084 3040 1090 3052
rect 5350 3040 5356 3052
rect 1084 3012 5356 3040
rect 1084 3000 1090 3012
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5460 3040 5488 3080
rect 6546 3068 6552 3120
rect 6604 3108 6610 3120
rect 11422 3108 11428 3120
rect 6604 3080 11428 3108
rect 6604 3068 6610 3080
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 11532 3108 11560 3148
rect 11609 3145 11621 3179
rect 11655 3176 11667 3179
rect 11698 3176 11704 3188
rect 11655 3148 11704 3176
rect 11655 3145 11667 3148
rect 11609 3139 11667 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 13814 3176 13820 3188
rect 11808 3148 13820 3176
rect 11808 3108 11836 3148
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 11532 3080 11836 3108
rect 7282 3040 7288 3052
rect 5460 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3040 7987 3043
rect 9950 3040 9956 3052
rect 7975 3012 9956 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 14182 3040 14188 3052
rect 10100 3012 14188 3040
rect 10100 3000 10106 3012
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 566 2932 572 2984
rect 624 2972 630 2984
rect 4982 2972 4988 2984
rect 624 2944 4988 2972
rect 624 2932 630 2944
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 11330 2972 11336 2984
rect 5776 2944 11336 2972
rect 5776 2932 5782 2944
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 198 2864 204 2916
rect 256 2904 262 2916
rect 4246 2904 4252 2916
rect 256 2876 4252 2904
rect 256 2864 262 2876
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 6822 2864 6828 2916
rect 6880 2904 6886 2916
rect 7101 2907 7159 2913
rect 7101 2904 7113 2907
rect 6880 2876 7113 2904
rect 6880 2864 6886 2876
rect 7101 2873 7113 2876
rect 7147 2904 7159 2907
rect 7929 2907 7987 2913
rect 7929 2904 7941 2907
rect 7147 2876 7941 2904
rect 7147 2873 7159 2876
rect 7101 2867 7159 2873
rect 7929 2873 7941 2876
rect 7975 2873 7987 2907
rect 7929 2867 7987 2873
rect 8110 2864 8116 2916
rect 8168 2904 8174 2916
rect 13722 2904 13728 2916
rect 8168 2876 13728 2904
rect 8168 2864 8174 2876
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 1854 2796 1860 2848
rect 1912 2836 1918 2848
rect 4706 2836 4712 2848
rect 1912 2808 4712 2836
rect 1912 2796 1918 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 10134 2836 10140 2848
rect 7524 2808 10140 2836
rect 7524 2796 7530 2808
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 10226 2796 10232 2848
rect 10284 2836 10290 2848
rect 10321 2839 10379 2845
rect 10321 2836 10333 2839
rect 10284 2808 10333 2836
rect 10284 2796 10290 2808
rect 10321 2805 10333 2808
rect 10367 2836 10379 2839
rect 14550 2836 14556 2848
rect 10367 2808 14556 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 10502 2592 10508 2644
rect 10560 2632 10566 2644
rect 11238 2632 11244 2644
rect 10560 2604 11244 2632
rect 10560 2592 10566 2604
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 11606 2496 11612 2508
rect 10652 2468 11612 2496
rect 10652 2456 10658 2468
rect 11606 2456 11612 2468
rect 11664 2456 11670 2508
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 11146 1776 11152 1828
rect 11204 1816 11210 1828
rect 12526 1816 12532 1828
rect 11204 1788 12532 1816
rect 11204 1776 11210 1788
rect 12526 1776 12532 1788
rect 12584 1776 12590 1828
rect 10134 1368 10140 1420
rect 10192 1408 10198 1420
rect 10778 1408 10784 1420
rect 10192 1380 10784 1408
rect 10192 1368 10198 1380
rect 10778 1368 10784 1380
rect 10836 1368 10842 1420
<< via1 >>
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 9864 17008 9916 17060
rect 10968 17008 11020 17060
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 4896 16396 4948 16448
rect 9312 16396 9364 16448
rect 9680 16396 9732 16448
rect 11796 16396 11848 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 7932 16124 7984 16176
rect 9680 16124 9732 16176
rect 6644 16056 6696 16108
rect 8852 16056 8904 16108
rect 9588 16056 9640 16108
rect 12624 16056 12676 16108
rect 9128 15988 9180 16040
rect 12164 15988 12216 16040
rect 3700 15920 3752 15972
rect 4068 15920 4120 15972
rect 5540 15920 5592 15972
rect 8208 15920 8260 15972
rect 8668 15920 8720 15972
rect 9680 15920 9732 15972
rect 1860 15852 1912 15904
rect 5632 15852 5684 15904
rect 8852 15852 8904 15904
rect 9956 15852 10008 15904
rect 10416 15852 10468 15904
rect 11336 15852 11388 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 1400 15648 1452 15700
rect 6460 15648 6512 15700
rect 10140 15648 10192 15700
rect 10324 15648 10376 15700
rect 15476 15648 15528 15700
rect 1032 15580 1084 15632
rect 3792 15580 3844 15632
rect 4068 15580 4120 15632
rect 5080 15580 5132 15632
rect 8024 15580 8076 15632
rect 10692 15580 10744 15632
rect 13636 15580 13688 15632
rect 16764 15580 16816 15632
rect 4528 15555 4580 15564
rect 4528 15521 4537 15555
rect 4537 15521 4571 15555
rect 4571 15521 4580 15555
rect 4528 15512 4580 15521
rect 6276 15512 6328 15564
rect 9956 15512 10008 15564
rect 10140 15512 10192 15564
rect 12716 15512 12768 15564
rect 7564 15444 7616 15496
rect 9588 15444 9640 15496
rect 11704 15444 11756 15496
rect 15936 15444 15988 15496
rect 2228 15376 2280 15428
rect 5540 15376 5592 15428
rect 11428 15376 11480 15428
rect 14280 15376 14332 15428
rect 4712 15308 4764 15360
rect 6736 15308 6788 15360
rect 7196 15308 7248 15360
rect 9588 15308 9640 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 572 15104 624 15156
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 5816 14832 5868 14884
rect 4528 14764 4580 14816
rect 9680 14764 9732 14816
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 204 14560 256 14612
rect 2596 14560 2648 14612
rect 6736 14560 6788 14612
rect 9588 14560 9640 14612
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 7104 14424 7156 14433
rect 10048 14424 10100 14476
rect 5540 14220 5592 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 13728 14016 13780 14068
rect 2596 13948 2648 14000
rect 2964 13948 3016 14000
rect 9128 13880 9180 13932
rect 6276 13855 6328 13864
rect 6276 13821 6285 13855
rect 6285 13821 6319 13855
rect 6319 13821 6328 13855
rect 6276 13812 6328 13821
rect 10048 13812 10100 13864
rect 13084 13812 13136 13864
rect 7104 13676 7156 13728
rect 9220 13676 9272 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 5540 13404 5592 13456
rect 3976 13268 4028 13320
rect 6920 13132 6972 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7748 13175 7800 13184
rect 7748 13141 7757 13175
rect 7757 13141 7791 13175
rect 7791 13141 7800 13175
rect 7748 13132 7800 13141
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 3976 12928 4028 12980
rect 5540 12928 5592 12980
rect 7196 12792 7248 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 7748 12724 7800 12776
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 7104 12588 7156 12640
rect 7748 12588 7800 12640
rect 8668 12588 8720 12640
rect 9128 12588 9180 12640
rect 13728 12588 13780 12640
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 6368 12384 6420 12436
rect 6736 12384 6788 12436
rect 4528 12316 4580 12368
rect 4712 12316 4764 12368
rect 6092 12291 6144 12300
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 6276 12044 6328 12096
rect 6828 12044 6880 12096
rect 8024 12044 8076 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 5540 11840 5592 11892
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 8024 11679 8076 11688
rect 8024 11645 8058 11679
rect 8058 11645 8076 11679
rect 8024 11636 8076 11645
rect 6092 11568 6144 11620
rect 7656 11568 7708 11620
rect 8116 11568 8168 11620
rect 9864 11568 9916 11620
rect 10140 11568 10192 11620
rect 11152 11500 11204 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 6828 11296 6880 11348
rect 8668 11339 8720 11348
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 9680 11296 9732 11348
rect 10416 11296 10468 11348
rect 2964 11203 3016 11212
rect 2964 11169 2982 11203
rect 2982 11169 3016 11203
rect 2964 11160 3016 11169
rect 5540 11160 5592 11212
rect 6644 11160 6696 11212
rect 7656 11228 7708 11280
rect 5816 11092 5868 11144
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 6920 11092 6972 11144
rect 10416 11160 10468 11212
rect 8668 11092 8720 11144
rect 7196 11024 7248 11076
rect 7288 11024 7340 11076
rect 9772 11024 9824 11076
rect 3332 10956 3384 11008
rect 9864 10956 9916 11008
rect 10232 10956 10284 11008
rect 10600 10956 10652 11008
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 2964 10795 3016 10804
rect 2964 10761 2973 10795
rect 2973 10761 3007 10795
rect 3007 10761 3016 10795
rect 2964 10752 3016 10761
rect 3332 10752 3384 10804
rect 3884 10752 3936 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 9680 10795 9732 10804
rect 6184 10752 6236 10761
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 9864 10752 9916 10804
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 6828 10548 6880 10600
rect 8576 10684 8628 10736
rect 9404 10684 9456 10736
rect 7656 10548 7708 10600
rect 3884 10523 3936 10532
rect 3884 10489 3893 10523
rect 3893 10489 3927 10523
rect 3927 10489 3936 10523
rect 4804 10523 4856 10532
rect 3884 10480 3936 10489
rect 4804 10489 4813 10523
rect 4813 10489 4847 10523
rect 4847 10489 4856 10523
rect 4804 10480 4856 10489
rect 1584 10412 1636 10464
rect 2964 10412 3016 10464
rect 8668 10480 8720 10532
rect 7288 10412 7340 10464
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 10416 10616 10468 10668
rect 10600 10480 10652 10532
rect 8944 10455 8996 10464
rect 7472 10412 7524 10421
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10232 10412 10284 10421
rect 10416 10412 10468 10464
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 7288 10208 7340 10260
rect 7656 10208 7708 10260
rect 8024 10208 8076 10260
rect 8760 10208 8812 10260
rect 9128 10208 9180 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 10324 10208 10376 10260
rect 1584 10183 1636 10192
rect 1584 10149 1593 10183
rect 1593 10149 1627 10183
rect 1627 10149 1636 10183
rect 1584 10140 1636 10149
rect 2780 10140 2832 10192
rect 4804 10140 4856 10192
rect 13084 10140 13136 10192
rect 7288 10115 7340 10124
rect 1952 10004 2004 10056
rect 5816 10004 5868 10056
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 8944 10072 8996 10124
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 9128 9936 9180 9988
rect 6920 9868 6972 9920
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 10232 9868 10284 9920
rect 10600 9868 10652 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 4344 9664 4396 9716
rect 5172 9664 5224 9716
rect 6368 9664 6420 9716
rect 8024 9664 8076 9716
rect 10324 9664 10376 9716
rect 7380 9596 7432 9648
rect 7472 9596 7524 9648
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 8760 9460 8812 9512
rect 9220 9596 9272 9648
rect 12900 9596 12952 9648
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 9404 9460 9456 9512
rect 4712 9392 4764 9444
rect 9496 9392 9548 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 5816 9120 5868 9172
rect 7380 9120 7432 9172
rect 8484 9120 8536 9172
rect 9680 9120 9732 9172
rect 7012 9052 7064 9104
rect 8024 9052 8076 9104
rect 7288 8984 7340 9036
rect 7840 8916 7892 8968
rect 8944 9052 8996 9104
rect 12716 8984 12768 9036
rect 11152 8916 11204 8968
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 7840 8576 7892 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 6920 8508 6972 8560
rect 8944 8440 8996 8492
rect 9680 8372 9732 8424
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 9772 8304 9824 8356
rect 12716 8347 12768 8356
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 8852 8236 8904 8288
rect 9128 8236 9180 8288
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 5724 7488 5776 7540
rect 2964 7216 3016 7268
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 7012 6332 7064 6384
rect 9864 6400 9916 6452
rect 10048 6332 10100 6384
rect 15476 6332 15528 6384
rect 10324 6128 10376 6180
rect 6368 6060 6420 6112
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 7656 6060 7708 6069
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 3148 5856 3200 5908
rect 8208 5856 8260 5908
rect 10692 5856 10744 5908
rect 5540 5788 5592 5840
rect 4160 5720 4212 5772
rect 6644 5720 6696 5772
rect 7840 5720 7892 5772
rect 9036 5720 9088 5772
rect 9772 5720 9824 5772
rect 11244 5720 11296 5772
rect 12256 5720 12308 5772
rect 5540 5652 5592 5704
rect 10232 5652 10284 5704
rect 10692 5652 10744 5704
rect 12808 5652 12860 5704
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 4528 5516 4580 5568
rect 7748 5584 7800 5636
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 7288 5516 7340 5568
rect 9312 5516 9364 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 5540 5312 5592 5364
rect 5632 5312 5684 5364
rect 8116 5312 8168 5364
rect 2688 5244 2740 5296
rect 7840 5287 7892 5296
rect 7840 5253 7849 5287
rect 7849 5253 7883 5287
rect 7883 5253 7892 5287
rect 7840 5244 7892 5253
rect 10508 5244 10560 5296
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 9864 5176 9916 5228
rect 7472 5108 7524 5160
rect 4068 5040 4120 5092
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 9312 5108 9364 5160
rect 11796 5176 11848 5228
rect 12992 5040 13044 5092
rect 8760 4972 8812 5024
rect 9036 4972 9088 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 9772 5015 9824 5024
rect 9772 4981 9781 5015
rect 9781 4981 9815 5015
rect 9815 4981 9824 5015
rect 9772 4972 9824 4981
rect 10324 5015 10376 5024
rect 10324 4981 10333 5015
rect 10333 4981 10367 5015
rect 10367 4981 10376 5015
rect 10324 4972 10376 4981
rect 11244 4972 11296 5024
rect 11336 4972 11388 5024
rect 12256 5015 12308 5024
rect 12256 4981 12265 5015
rect 12265 4981 12299 5015
rect 12299 4981 12308 5015
rect 12256 4972 12308 4981
rect 15936 4972 15988 5024
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 3976 4768 4028 4820
rect 9956 4768 10008 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 5172 4700 5224 4752
rect 9220 4700 9272 4752
rect 10784 4700 10836 4752
rect 13820 4700 13872 4752
rect 4896 4632 4948 4684
rect 6000 4632 6052 4684
rect 6460 4632 6512 4684
rect 8668 4632 8720 4684
rect 10048 4632 10100 4684
rect 11428 4632 11480 4684
rect 12716 4632 12768 4684
rect 13636 4632 13688 4684
rect 6736 4564 6788 4616
rect 11336 4564 11388 4616
rect 5448 4496 5500 4548
rect 10324 4496 10376 4548
rect 12440 4496 12492 4548
rect 16212 4496 16264 4548
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 9956 4428 10008 4480
rect 10600 4428 10652 4480
rect 11336 4428 11388 4480
rect 13728 4471 13780 4480
rect 13728 4437 13737 4471
rect 13737 4437 13771 4471
rect 13771 4437 13780 4471
rect 13728 4428 13780 4437
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 4896 4267 4948 4276
rect 4896 4233 4905 4267
rect 4905 4233 4939 4267
rect 4939 4233 4948 4267
rect 4896 4224 4948 4233
rect 6000 4267 6052 4276
rect 6000 4233 6009 4267
rect 6009 4233 6043 4267
rect 6043 4233 6052 4267
rect 6000 4224 6052 4233
rect 10140 4224 10192 4276
rect 10784 4267 10836 4276
rect 10784 4233 10793 4267
rect 10793 4233 10827 4267
rect 10827 4233 10836 4267
rect 10784 4224 10836 4233
rect 11428 4224 11480 4276
rect 13636 4267 13688 4276
rect 3148 4088 3200 4140
rect 1400 3952 1452 4004
rect 6092 3952 6144 4004
rect 6368 4088 6420 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 8760 4156 8812 4208
rect 10600 4156 10652 4208
rect 13636 4233 13645 4267
rect 13645 4233 13679 4267
rect 13679 4233 13688 4267
rect 13636 4224 13688 4233
rect 15108 4156 15160 4208
rect 7840 4088 7892 4097
rect 8484 4088 8536 4140
rect 10692 4088 10744 4140
rect 12992 4088 13044 4140
rect 14648 4088 14700 4140
rect 10784 4020 10836 4072
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 2320 3884 2372 3936
rect 8208 3952 8260 4004
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 12716 3884 12768 3936
rect 16764 3884 16816 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 6276 3680 6328 3732
rect 12256 3680 12308 3732
rect 16304 3680 16356 3732
rect 4804 3612 4856 3664
rect 9220 3612 9272 3664
rect 9312 3612 9364 3664
rect 11060 3612 11112 3664
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 7564 3544 7616 3596
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 8484 3544 8536 3596
rect 9036 3544 9088 3596
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 11520 3587 11572 3596
rect 11520 3553 11535 3587
rect 11535 3553 11569 3587
rect 11569 3553 11572 3587
rect 11520 3544 11572 3553
rect 5264 3476 5316 3528
rect 10324 3476 10376 3528
rect 11244 3476 11296 3528
rect 15016 3476 15068 3528
rect 3976 3408 4028 3460
rect 8576 3408 8628 3460
rect 12072 3408 12124 3460
rect 2688 3340 2740 3392
rect 7380 3340 7432 3392
rect 11796 3340 11848 3392
rect 13176 3340 13228 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 4436 3136 4488 3188
rect 7656 3136 7708 3188
rect 8116 3179 8168 3188
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 8668 3136 8720 3188
rect 9128 3136 9180 3188
rect 9772 3136 9824 3188
rect 3792 3068 3844 3120
rect 1032 3000 1084 3052
rect 5356 3000 5408 3052
rect 6552 3068 6604 3120
rect 11428 3068 11480 3120
rect 11704 3136 11756 3188
rect 13820 3136 13872 3188
rect 7288 3000 7340 3052
rect 9956 3000 10008 3052
rect 10048 3000 10100 3052
rect 14188 3000 14240 3052
rect 572 2932 624 2984
rect 4988 2932 5040 2984
rect 5724 2932 5776 2984
rect 11336 2932 11388 2984
rect 204 2864 256 2916
rect 4252 2864 4304 2916
rect 6828 2864 6880 2916
rect 8116 2864 8168 2916
rect 13728 2864 13780 2916
rect 1860 2796 1912 2848
rect 4712 2796 4764 2848
rect 7472 2796 7524 2848
rect 10140 2796 10192 2848
rect 10232 2796 10284 2848
rect 14556 2796 14608 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 10508 2592 10560 2644
rect 11244 2592 11296 2644
rect 10600 2456 10652 2508
rect 11612 2456 11664 2508
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 11152 1776 11204 1828
rect 12532 1776 12584 1828
rect 10140 1368 10192 1420
rect 10784 1368 10836 1420
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1858 19200 1914 20000
rect 2226 19200 2282 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3514 19200 3570 20000
rect 3882 19200 3938 20000
rect 4342 19200 4398 20000
rect 4710 19200 4766 20000
rect 5170 19200 5226 20000
rect 5538 19200 5594 20000
rect 5998 19200 6054 20000
rect 6366 19200 6422 20000
rect 6826 19200 6882 20000
rect 7194 19200 7250 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8482 19200 8538 20000
rect 8850 19200 8906 20000
rect 9310 19200 9366 20000
rect 9678 19200 9734 20000
rect 10138 19200 10194 20000
rect 10506 19200 10562 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11794 19200 11850 20000
rect 12162 19200 12218 20000
rect 12622 19200 12678 20000
rect 12990 19200 13046 20000
rect 13450 19200 13506 20000
rect 13818 19200 13874 20000
rect 14278 19200 14334 20000
rect 14646 19200 14702 20000
rect 15106 19200 15162 20000
rect 15474 19200 15530 20000
rect 15934 19200 15990 20000
rect 16302 19200 16358 20000
rect 16762 19200 16818 20000
rect 216 14618 244 19200
rect 584 15162 612 19200
rect 1044 15638 1072 19200
rect 1412 15706 1440 19200
rect 1872 15910 1900 19200
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 1032 15632 1084 15638
rect 1032 15574 1084 15580
rect 2240 15434 2268 19200
rect 2228 15428 2280 15434
rect 2228 15370 2280 15376
rect 572 15156 624 15162
rect 572 15098 624 15104
rect 204 14612 256 14618
rect 204 14554 256 14560
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 14006 2636 14554
rect 2596 14000 2648 14006
rect 2596 13942 2648 13948
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10198 1624 10406
rect 1584 10192 1636 10198
rect 1584 10134 1636 10140
rect 1596 9382 1624 10134
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9382 1992 9998
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1596 8401 1624 9318
rect 1582 8392 1638 8401
rect 1582 8327 1638 8336
rect 1400 4004 1452 4010
rect 1400 3946 1452 3952
rect 1032 3052 1084 3058
rect 1032 2994 1084 3000
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 204 2916 256 2922
rect 204 2858 256 2864
rect 216 800 244 2858
rect 584 800 612 2926
rect 1044 800 1072 2994
rect 1412 800 1440 3946
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 800 1900 2790
rect 1964 1737 1992 9318
rect 2700 5302 2728 19200
rect 3068 19122 3096 19200
rect 3068 19094 3188 19122
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 10198 2820 14991
rect 2964 14000 3016 14006
rect 2964 13942 3016 13948
rect 2976 11218 3004 13942
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2976 10810 3004 11154
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2976 10470 3004 10746
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2976 5001 3004 7210
rect 3160 5914 3188 19094
rect 3528 17626 3556 19200
rect 3896 19122 3924 19200
rect 3896 19094 4108 19122
rect 3974 18320 4030 18329
rect 3974 18255 4030 18264
rect 3528 17598 3832 17626
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3712 15450 3740 15914
rect 3804 15638 3832 17598
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3712 15422 3832 15450
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3804 12458 3832 15422
rect 3988 13326 4016 18255
rect 4080 15978 4108 19094
rect 4068 15972 4120 15978
rect 4068 15914 4120 15920
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3988 12986 4016 13262
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3804 12430 4016 12458
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3790 11656 3846 11665
rect 3790 11591 3846 11600
rect 3804 11354 3832 11591
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10810 3372 10950
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3804 10674 3832 11290
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3896 10538 3924 10746
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 2962 4992 3018 5001
rect 2962 4927 3018 4936
rect 3988 4826 4016 12430
rect 4080 5098 4108 15574
rect 4356 9722 4384 19200
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4540 14822 4568 15506
rect 4724 15366 4752 19200
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 12374 4568 14758
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4724 9450 4752 12310
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4816 10198 4844 10474
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5370 4200 5714
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1950 1728 2006 1737
rect 1950 1663 2006 1672
rect 2332 800 2360 3878
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2700 800 2728 3334
rect 3160 800 3188 4082
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3804 1442 3832 3062
rect 3620 1414 3832 1442
rect 3620 800 3648 1414
rect 3988 800 4016 3402
rect 4264 2922 4292 5510
rect 4540 5166 4568 5510
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4448 800 4476 3130
rect 4724 2854 4752 4966
rect 4908 4690 4936 16390
rect 5184 15858 5212 19200
rect 5552 15978 5580 19200
rect 6012 17082 6040 19200
rect 6012 17054 6316 17082
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5632 15904 5684 15910
rect 5184 15830 5488 15858
rect 5632 15846 5684 15852
rect 5080 15632 5132 15638
rect 5080 15574 5132 15580
rect 5092 6458 5120 15574
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5184 4758 5212 9658
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 4282 4936 4626
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4816 800 4844 3606
rect 5000 2990 5028 4422
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5276 800 5304 3470
rect 5368 3058 5396 5510
rect 5460 4554 5488 15830
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 15162 5580 15370
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13462 5580 14214
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 12986 5580 13398
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5552 11898 5580 12922
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 5846 5580 11154
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5370 5580 5646
rect 5644 5370 5672 15846
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 6288 15570 6316 17054
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5828 11150 5856 14826
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6288 13870 6316 14418
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6104 11626 6132 12242
rect 6288 12102 6316 13806
rect 6380 12442 6408 19200
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6196 10810 6224 11086
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 7546 5764 9862
rect 5828 9382 5856 9998
rect 6380 9722 6408 9998
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9178 5856 9318
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 6012 4282 6040 4626
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 4010 6132 4422
rect 6380 4146 6408 6054
rect 6472 4690 6500 15642
rect 6656 11218 6684 16050
rect 6840 15994 6868 19200
rect 6840 15966 7052 15994
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6748 14618 6776 15302
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 5778 6684 9454
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6748 4622 6776 12378
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11354 6868 12038
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6840 10606 6868 11290
rect 6932 11150 6960 13126
rect 7024 12730 7052 15966
rect 7208 15366 7236 19200
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7116 13734 7144 14418
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12850 7512 13126
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7024 12702 7144 12730
rect 7116 12646 7144 12702
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 8566 6960 9862
rect 7024 9110 7052 12582
rect 7208 11082 7236 12786
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7300 10470 7328 11018
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7300 10130 7328 10202
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 7300 9042 7328 10066
rect 7392 9654 7420 12718
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 9654 7512 10406
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7392 8634 7420 9114
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5736 800 5764 2926
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6288 1442 6316 3674
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6104 1414 6316 1442
rect 6104 800 6132 1414
rect 6564 800 6592 3062
rect 6840 2922 6868 3538
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 7024 800 7052 6326
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 3058 7328 5510
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 5030 7512 5102
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7392 800 7420 3334
rect 7484 2854 7512 4966
rect 7576 3602 7604 15438
rect 7668 11626 7696 19200
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12782 7788 13126
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7668 10606 7696 11222
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10266 7696 10542
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7668 3194 7696 6054
rect 7760 5642 7788 12582
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 8634 7880 8910
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7852 5302 7880 5714
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7944 4162 7972 16118
rect 8036 15638 8064 19200
rect 8496 17626 8524 19200
rect 8496 17598 8708 17626
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8680 15978 8708 17598
rect 8864 16114 8892 19200
rect 9324 16454 9352 19200
rect 9692 17218 9720 19200
rect 9692 17190 9996 17218
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9692 16182 9720 16390
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9128 16040 9180 16046
rect 9048 16000 9128 16028
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11694 8064 12038
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8036 10266 8064 11630
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8036 9722 8064 10202
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8036 8634 8064 9046
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8128 5370 8156 11562
rect 8220 5914 8248 15914
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8680 11354 8708 12582
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8680 11150 8708 11290
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8588 10146 8616 10678
rect 8680 10538 8708 11086
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8680 10282 8708 10474
rect 8680 10266 8800 10282
rect 8680 10260 8812 10266
rect 8680 10254 8760 10260
rect 8760 10202 8812 10208
rect 8588 10118 8708 10146
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8680 9330 8708 10118
rect 8864 9602 8892 15846
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8956 10130 8984 10406
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8772 9574 8892 9602
rect 8772 9518 8800 9574
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8496 9178 8524 9318
rect 8680 9302 8892 9330
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8588 8090 8616 8298
rect 8864 8294 8892 9302
rect 8956 9110 8984 10066
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8956 8498 8984 9046
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 9048 5778 9076 16000
rect 9128 15982 9180 15988
rect 9600 15502 9628 16050
rect 9678 16008 9734 16017
rect 9678 15943 9680 15952
rect 9732 15943 9734 15952
rect 9680 15914 9732 15920
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9600 14618 9628 15302
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9140 12646 9168 13874
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 11898 9168 12582
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9140 9994 9168 10202
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9140 9586 9168 9930
rect 9232 9654 9260 13670
rect 9692 11506 9720 14758
rect 9876 11626 9904 17002
rect 9968 15910 9996 17190
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 10152 15706 10180 19200
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9692 11478 9904 11506
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9692 10810 9720 11290
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9416 10266 9444 10678
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9416 9518 9444 10202
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 9048 5030 9076 5714
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 7852 4146 7972 4162
rect 7840 4140 7972 4146
rect 7892 4134 7972 4140
rect 8484 4140 8536 4146
rect 7840 4082 7892 4088
rect 8484 4082 8536 4088
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 3194 8156 3538
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8220 3074 8248 3946
rect 8496 3602 8524 4082
rect 8576 3936 8628 3942
rect 8680 3924 8708 4626
rect 8772 4214 8800 4966
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8628 3896 8708 3924
rect 8576 3878 8628 3884
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8588 3466 8616 3878
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 7852 3046 8248 3074
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7852 800 7880 3046
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 8128 898 8156 2858
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8128 870 8248 898
rect 8220 800 8248 870
rect 8680 800 8708 3130
rect 9048 898 9076 3538
rect 9140 3194 9168 8230
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5166 9352 5510
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9232 4758 9260 4966
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3670 9260 3878
rect 9324 3670 9352 5102
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9048 870 9168 898
rect 9140 800 9168 870
rect 9508 800 9536 9386
rect 9692 9178 9720 9862
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9692 8430 9720 9114
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9784 8362 9812 11018
rect 9876 11014 9904 11478
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9876 6458 9904 10746
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9784 5030 9812 5714
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9784 3194 9812 4966
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 2938 9904 5170
rect 9968 4826 9996 15506
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10060 13870 10088 14418
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10060 10130 10088 13806
rect 10152 12458 10180 15506
rect 10336 12730 10364 15642
rect 10428 12866 10456 15846
rect 10520 13002 10548 19200
rect 10980 17066 11008 19200
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 11348 15910 11376 19200
rect 11808 16454 11836 19200
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 12176 16046 12204 19200
rect 12636 16114 12664 19200
rect 13004 17762 13032 19200
rect 12728 17734 13032 17762
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12622 16008 12678 16017
rect 12622 15943 12678 15952
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10520 12974 10640 13002
rect 10428 12838 10548 12866
rect 10336 12702 10456 12730
rect 10152 12430 10364 12458
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10060 9382 10088 10066
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 6390 10088 9318
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9968 3058 9996 4422
rect 10060 3942 10088 4626
rect 10152 4282 10180 11562
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10470 10272 10950
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10336 10266 10364 12430
rect 10428 11354 10456 12702
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 10674 10456 11154
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 5710 10272 9862
rect 10336 9722 10364 10202
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10336 6186 10364 9658
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10336 4554 10364 4966
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10060 3058 10088 3878
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9876 2910 9996 2938
rect 9968 800 9996 2910
rect 10244 2854 10272 3538
rect 10336 3534 10364 3878
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10152 1426 10180 2790
rect 10140 1420 10192 1426
rect 10140 1362 10192 1368
rect 10428 800 10456 10406
rect 10520 9602 10548 12838
rect 10612 11014 10640 12974
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10612 10538 10640 10950
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10612 9926 10640 10474
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10520 9574 10640 9602
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10520 2650 10548 5238
rect 10612 4486 10640 9574
rect 10704 5914 10732 15574
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 11164 8974 11192 11494
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10612 2514 10640 4150
rect 10704 4146 10732 5646
rect 11256 5030 11284 5714
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10796 4282 10824 4694
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10796 4078 10824 4218
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11072 3516 11100 3606
rect 11256 3534 11284 4966
rect 11348 4622 11376 4966
rect 11440 4690 11468 15370
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11244 3528 11296 3534
rect 11072 3488 11192 3516
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 11164 1834 11192 3488
rect 11244 3470 11296 3476
rect 11348 2990 11376 4422
rect 11440 4282 11468 4626
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3126 11468 3878
rect 11520 3596 11572 3602
rect 11716 3584 11744 15438
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11572 3556 11744 3584
rect 11520 3538 11572 3544
rect 11716 3194 11744 3556
rect 11808 3398 11836 5170
rect 12268 5030 12296 5714
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12268 3738 12296 4966
rect 12636 4826 12664 15943
rect 12728 15570 12756 17734
rect 13464 17626 13492 19200
rect 12820 17598 13492 17626
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 8362 12756 8978
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 7449 12756 8298
rect 12714 7440 12770 7449
rect 12714 7375 12770 7384
rect 12820 5710 12848 17598
rect 13726 17504 13782 17513
rect 13282 17436 13578 17456
rect 13726 17439 13782 17448
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13096 10198 13124 13806
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12452 4078 12480 4490
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12728 3942 12756 4626
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11152 1828 11204 1834
rect 11152 1770 11204 1776
rect 10784 1420 10836 1426
rect 10784 1362 10836 1368
rect 10796 800 10824 1362
rect 11256 800 11284 2586
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 11624 800 11652 2450
rect 12084 800 12112 3402
rect 12532 1828 12584 1834
rect 12532 1770 12584 1776
rect 12544 800 12572 1770
rect 12912 800 12940 9590
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 13004 4146 13032 5034
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13096 2553 13124 10134
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13648 4690 13676 15574
rect 13740 14074 13768 17439
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12481 13768 12582
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13832 4758 13860 19200
rect 14292 15434 14320 19200
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13648 4282 13676 4626
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13082 2544 13138 2553
rect 13082 2479 13138 2488
rect 13188 1986 13216 3334
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13740 2922 13768 4422
rect 14660 4298 14688 19200
rect 14568 4270 14688 4298
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13188 1958 13400 1986
rect 13372 800 13400 1958
rect 13832 800 13860 3130
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14200 800 14228 2994
rect 14568 2854 14596 4270
rect 15120 4214 15148 19200
rect 15488 15706 15516 19200
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15948 15502 15976 19200
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 16316 12458 16344 19200
rect 16776 15638 16804 19200
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16224 12430 16344 12458
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14660 800 14688 4082
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15028 800 15056 3470
rect 15488 800 15516 6326
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 800 15976 4966
rect 16224 4554 16252 12430
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16316 800 16344 3674
rect 16776 800 16804 3878
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6550 0 6606 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 12070 0 12126 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16762 0 16818 800
<< via2 >>
rect 1582 8336 1638 8392
rect 2778 15000 2834 15056
rect 3974 18264 4030 18320
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3790 11600 3846 11656
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 2962 4936 3018 4992
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 1950 1672 2006 1728
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 9678 15972 9734 16008
rect 9678 15952 9680 15972
rect 9680 15952 9732 15972
rect 9732 15952 9734 15972
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 12622 15952 12678 16008
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 12714 7384 12770 7440
rect 13726 17448 13782 17504
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13726 12416 13782 12472
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13082 2488 13138 2544
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
<< metal3 >>
rect 0 18322 800 18352
rect 3969 18322 4035 18325
rect 0 18320 4035 18322
rect 0 18264 3974 18320
rect 4030 18264 4035 18320
rect 0 18262 4035 18264
rect 0 18232 800 18262
rect 3969 18259 4035 18262
rect 13721 17506 13787 17509
rect 16200 17506 17000 17536
rect 13721 17504 17000 17506
rect 13721 17448 13726 17504
rect 13782 17448 17000 17504
rect 13721 17446 17000 17448
rect 13721 17443 13787 17446
rect 3409 17440 3729 17441
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 16200 17416 17000 17446
rect 13270 17375 13590 17376
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 9673 16010 9739 16013
rect 12617 16010 12683 16013
rect 9673 16008 12683 16010
rect 9673 15952 9678 16008
rect 9734 15952 12622 16008
rect 12678 15952 12683 16008
rect 9673 15950 12683 15952
rect 9673 15947 9739 15950
rect 12617 15947 12683 15950
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 0 15058 800 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 800 14998
rect 2773 14995 2839 14998
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 13721 12474 13787 12477
rect 16200 12474 17000 12504
rect 13721 12472 17000 12474
rect 13721 12416 13726 12472
rect 13782 12416 17000 12472
rect 13721 12414 17000 12416
rect 13721 12411 13787 12414
rect 16200 12384 17000 12414
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 0 11658 800 11688
rect 3785 11658 3851 11661
rect 0 11656 3851 11658
rect 0 11600 3790 11656
rect 3846 11600 3851 11656
rect 0 11598 3851 11600
rect 0 11568 800 11598
rect 3785 11595 3851 11598
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 0 8394 800 8424
rect 1577 8394 1643 8397
rect 0 8392 1643 8394
rect 0 8336 1582 8392
rect 1638 8336 1643 8392
rect 0 8334 1643 8336
rect 0 8304 800 8334
rect 1577 8331 1643 8334
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 12709 7442 12775 7445
rect 16200 7442 17000 7472
rect 12709 7440 17000 7442
rect 12709 7384 12714 7440
rect 12770 7384 17000 7440
rect 12709 7382 17000 7384
rect 12709 7379 12775 7382
rect 16200 7352 17000 7382
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 0 4994 800 5024
rect 2957 4994 3023 4997
rect 0 4992 3023 4994
rect 0 4936 2962 4992
rect 3018 4936 3023 4992
rect 0 4934 3023 4936
rect 0 4904 800 4934
rect 2957 4931 3023 4934
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 13077 2546 13143 2549
rect 16200 2546 17000 2576
rect 13077 2544 17000 2546
rect 13077 2488 13082 2544
rect 13138 2488 17000 2544
rect 13077 2486 17000 2488
rect 13077 2483 13143 2486
rect 16200 2456 17000 2486
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 0 1730 800 1760
rect 1945 1730 2011 1733
rect 0 1728 2011 1730
rect 0 1672 1950 1728
rect 2006 1672 2011 1728
rect 0 1670 2011 1672
rect 0 1640 800 1670
rect 1945 1667 2011 1670
<< via3 >>
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
<< metal4 >>
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 15264 3729 16288
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5874 15808 6195 16832
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 15264 8660 16288
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 16896 11125 17456
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 15808 11125 16832
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 11456 11125 12480
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2128 11125 2688
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 16352 13590 17376
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608764133
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608764133
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608764133
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608764133
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1608764133
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_149
timestamp 1608764133
transform 1 0 14812 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1608764133
transform 1 0 15456 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1608764133
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1608764133
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1608764133
transform 1 0 13708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608764133
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1608764133
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1608764133
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_106
timestamp 1608764133
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_118
timestamp 1608764133
transform 1 0 11960 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1608764133
transform 1 0 12604 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608764133
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608764133
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1608764133
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_87
timestamp 1608764133
transform 1 0 9108 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1608764133
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1608764133
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1608764133
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_63
timestamp 1608764133
transform 1 0 6900 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_75
timestamp 1608764133
transform 1 0 8004 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608764133
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1608764133
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1608764133
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1608764133
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_56
timestamp 1608764133
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608764133
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608764133
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608764133
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1608764133
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1608764133
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1608764133
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608764133
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608764133
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608764133
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1608764133
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1608764133
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1608764133
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608764133
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_147
timestamp 1608764133
transform 1 0 14628 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1608764133
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1608764133
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608764133
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1608764133
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1608764133
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1608764133
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1608764133
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1608764133
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608764133
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1608764133
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608764133
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1608764133
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1608764133
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1608764133
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608764133
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608764133
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1608764133
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608764133
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608764133
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1608764133
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1608764133
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1608764133
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1608764133
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1608764133
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608764133
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1608764133
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1608764133
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1608764133
transform 1 0 7084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_77
timestamp 1608764133
transform 1 0 8188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1608764133
transform 1 0 5980 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608764133
transform 1 0 4508 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608764133
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1608764133
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1608764133
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_36
timestamp 1608764133
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1608764133
transform 1 0 4876 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608764133
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1608764133
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1608764133
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608764133
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1608764133
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1608764133
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1608764133
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608764133
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1608764133
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1608764133
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1608764133
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1608764133
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1608764133
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1608764133
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608764133
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__03__A
timestamp 1608764133
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_45
timestamp 1608764133
transform 1 0 5244 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_50
timestamp 1608764133
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_54
timestamp 1608764133
transform 1 0 6072 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608764133
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1608764133
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608764133
transform 1 0 3772 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1608764133
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1608764133
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1608764133
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1608764133
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_37
timestamp 1608764133
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_41
timestamp 1608764133
transform 1 0 4876 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608764133
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1608764133
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1608764133
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608764133
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608764133
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1608764133
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_133
timestamp 1608764133
transform 1 0 13340 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1608764133
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1608764133
transform 1 0 11132 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1608764133
transform 1 0 12236 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1608764133
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608764133
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1608764133
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1608764133
transform 1 0 10028 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1608764133
transform 1 0 7084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_69
timestamp 1608764133
transform 1 0 7452 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_81
timestamp 1608764133
transform 1 0 8556 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764133
transform 1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_44
timestamp 1608764133
transform 1 0 5152 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1608764133
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_57
timestamp 1608764133
transform 1 0 6348 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608764133
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_28
timestamp 1608764133
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608764133
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608764133
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608764133
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608764133
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_15
timestamp 1608764133
transform 1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1608764133
transform 1 0 2944 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608764133
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1608764133
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1608764133
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1608764133
transform 1 0 15180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1608764133
transform 1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1608764133
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_143
timestamp 1608764133
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608764133
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_107
timestamp 1608764133
transform 1 0 10948 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1608764133
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608764133
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1608764133
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_91
timestamp 1608764133
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_95
timestamp 1608764133
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1608764133
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_67
timestamp 1608764133
transform 1 0 7268 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_79
timestamp 1608764133
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608764133
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1608764133
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1608764133
transform 1 0 5060 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1608764133
transform 1 0 6164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1608764133
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_62
timestamp 1608764133
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_A
timestamp 1608764133
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1608764133
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1608764133
transform 1 0 3956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1608764133
transform 1 0 2760 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608764133
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608764133
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_15
timestamp 1608764133
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608764133
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608764133
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608764133
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_147
timestamp 1608764133
transform 1 0 14628 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1608764133
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1608764133
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608764133
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1608764133
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608764133
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608764133
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1608764133
transform 1 0 11500 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1608764133
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608764133
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608764133
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608764133
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608764133
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_89
timestamp 1608764133
transform 1 0 9292 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_101
timestamp 1608764133
transform 1 0 10396 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_86
timestamp 1608764133
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608764133
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_77
timestamp 1608764133
transform 1 0 8188 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1608764133
transform 1 0 7912 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1608764133
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_73
timestamp 1608764133
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1608764133
transform 1 0 6992 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1608764133
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1608764133
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_63
timestamp 1608764133
transform 1 0 6900 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1608764133
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1608764133
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608764133
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608764133
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1608764133
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_56
timestamp 1608764133
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1608764133
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1608764133
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_51
timestamp 1608764133
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764133
transform 1 0 4324 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608764133
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608764133
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1608764133
transform 1 0 3588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_35
timestamp 1608764133
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1608764133
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608764133
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1608764133
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608764133
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608764133
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608764133
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608764133
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608764133
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608764133
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608764133
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608764133
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1608764133
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1608764133
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1608764133
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1608764133
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1608764133
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608764133
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608764133
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1608764133
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608764133
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_74
timestamp 1608764133
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_78
timestamp 1608764133
transform 1 0 8280 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764133
transform 1 0 6072 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_18_44
timestamp 1608764133
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1608764133
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608764133
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608764133
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608764133
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608764133
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608764133
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608764133
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608764133
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_147
timestamp 1608764133
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1608764133
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1608764133
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608764133
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_112
timestamp 1608764133
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608764133
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1608764133
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_88
timestamp 1608764133
transform 1 0 9200 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_100
timestamp 1608764133
transform 1 0 10304 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608764133
transform 1 0 7728 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1608764133
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608764133
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1608764133
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_51
timestamp 1608764133
transform 1 0 5796 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1608764133
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1608764133
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1608764133
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1608764133
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1608764133
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608764133
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608764133
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608764133
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608764133
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608764133
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1608764133
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1608764133
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_130
timestamp 1608764133
transform 1 0 13064 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_142
timestamp 1608764133
transform 1 0 14168 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_106
timestamp 1608764133
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_118
timestamp 1608764133
transform 1 0 11960 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1608764133
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608764133
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1608764133
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1608764133
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1608764133
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1608764133
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1608764133
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608764133
transform 1 0 7268 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1608764133
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1608764133
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_83
timestamp 1608764133
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1608764133
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1608764133
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_44
timestamp 1608764133
transform 1 0 5152 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1608764133
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608764133
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608764133
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1608764133
transform 1 0 3128 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1608764133
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608764133
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1608764133
transform 1 0 2852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608764133
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608764133
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1608764133
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608764133
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_147
timestamp 1608764133
transform 1 0 14628 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1608764133
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1608764133
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _01_
timestamp 1608764133
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608764133
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1608764133
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1608764133
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1608764133
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1608764133
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1608764133
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1608764133
transform 1 0 9752 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1608764133
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1608764133
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1608764133
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1608764133
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1608764133
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608764133
transform 1 0 7544 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1608764133
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1608764133
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1608764133
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608764133
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608764133
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1608764133
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1608764133
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_49
timestamp 1608764133
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_52
timestamp 1608764133
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_56
timestamp 1608764133
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1608764133
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608764133
transform 1 0 3680 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_TE_B
timestamp 1608764133
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1608764133
transform 1 0 3128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_41
timestamp 1608764133
transform 1 0 4876 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608764133
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR_A
timestamp 1608764133
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608764133
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1608764133
transform 1 0 2484 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_19
timestamp 1608764133
transform 1 0 2852 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608764133
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608764133
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608764133
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_147
timestamp 1608764133
transform 1 0 14628 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1608764133
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1608764133
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1608764133
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1608764133
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_130
timestamp 1608764133
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_142
timestamp 1608764133
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608764133
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1608764133
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_107
timestamp 1608764133
transform 1 0 10948 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1608764133
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1608764133
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_106
timestamp 1608764133
transform 1 0 10856 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_118
timestamp 1608764133
transform 1 0 11960 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1608764133
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1608764133
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1608764133
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1608764133
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_103
timestamp 1608764133
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1608764133
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1608764133
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608764133
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1608764133
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1608764133
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1608764133
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_89
timestamp 1608764133
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_93
timestamp 1608764133
transform 1 0 9660 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_87
timestamp 1608764133
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1608764133
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608764133
transform 1 0 7268 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1608764133
transform 1 0 8464 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1608764133
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1608764133
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_76
timestamp 1608764133
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_83
timestamp 1608764133
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1608764133
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1608764133
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_72
timestamp 1608764133
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1608764133
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_62
timestamp 1608764133
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608764133
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1608764133
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1608764133
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1608764133
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1608764133
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_56
timestamp 1608764133
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1608764133
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1608764133
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1608764133
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 1608764133
transform 1 0 5428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_44
timestamp 1608764133
transform 1 0 5152 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608764133
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_23
timestamp 1608764133
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_35
timestamp 1608764133
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1608764133
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608764133
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608764133
transform 1 0 1380 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608764133
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608764133
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_TE_B
timestamp 1608764133
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608764133
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1608764133
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1608764133
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_11
timestamp 1608764133
transform 1 0 2116 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_16
timestamp 1608764133
transform 1 0 2576 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608764133
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608764133
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1608764133
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_133
timestamp 1608764133
transform 1 0 13340 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1608764133
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608764133
transform 1 0 12236 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1608764133
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1608764133
transform 1 0 11868 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608764133
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1608764133
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1608764133
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1608764133
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1608764133
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1608764133
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1608764133
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1608764133
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1608764133
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_80
timestamp 1608764133
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608764133
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_56
timestamp 1608764133
transform 1 0 6256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608764133
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608764133
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608764133
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608764133
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608764133
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608764133
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608764133
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_151
timestamp 1608764133
transform 1 0 14996 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1608764133
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1608764133
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608764133
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608764133
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1608764133
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1608764133
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1608764133
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_86
timestamp 1608764133
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_90
timestamp 1608764133
transform 1 0 9384 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_102
timestamp 1608764133
transform 1 0 10488 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1608764133
transform 1 0 8188 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1608764133
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1608764133
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1608764133
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_66
timestamp 1608764133
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1608764133
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_73
timestamp 1608764133
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608764133
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608764133
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608764133
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1608764133
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608764133
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608764133
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608764133
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608764133
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608764133
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608764133
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608764133
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1608764133
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1608764133
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1608764133
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1608764133
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1608764133
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608764133
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1608764133
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1608764133
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1608764133
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1608764133
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_80
timestamp 1608764133
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_83
timestamp 1608764133
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608764133
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608764133
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608764133
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608764133
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608764133
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608764133
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608764133
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608764133
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608764133
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_147
timestamp 1608764133
transform 1 0 14628 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1608764133
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1608764133
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608764133
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1608764133
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608764133
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1608764133
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1608764133
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1608764133
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608764133
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_46
timestamp 1608764133
transform 1 0 5336 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1608764133
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608764133
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608764133
transform 1 0 3312 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608764133
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_23
timestamp 1608764133
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_30
timestamp 1608764133
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_34
timestamp 1608764133
transform 1 0 4232 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608764133
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608764133
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1608764133
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608764133
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608764133
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1608764133
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1608764133
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1608764133
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1608764133
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1608764133
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608764133
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1608764133
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1608764133
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1608764133
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608764133
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608764133
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608764133
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608764133
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608764133
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608764133
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608764133
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608764133
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608764133
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608764133
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608764133
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_146
timestamp 1608764133
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1608764133
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1608764133
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_147
timestamp 1608764133
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1608764133
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_134
timestamp 1608764133
transform 1 0 13432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1608764133
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1608764133
transform 1 0 10764 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1608764133
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608764133
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 1608764133
transform 1 0 11132 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_117
timestamp 1608764133
transform 1 0 11868 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_122
timestamp 1608764133
transform 1 0 12328 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_107
timestamp 1608764133
transform 1 0 10948 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1608764133
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1608764133
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_95
timestamp 1608764133
transform 1 0 9844 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1608764133
transform 1 0 10028 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1608764133
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608764133
transform 1 0 9108 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608764133
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__08__A
timestamp 1608764133
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1608764133
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1608764133
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1608764133
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1608764133
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1608764133
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1608764133
transform 1 0 8096 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1608764133
transform 1 0 7452 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1608764133
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_68
timestamp 1608764133
transform 1 0 7360 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_80
timestamp 1608764133
transform 1 0 8464 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1608764133
transform 1 0 7360 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_73
timestamp 1608764133
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_77
timestamp 1608764133
transform 1 0 8188 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1608764133
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608764133
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1608764133
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_48
timestamp 1608764133
transform 1 0 5520 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1608764133
transform 1 0 6624 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1608764133
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_49
timestamp 1608764133
transform 1 0 5612 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1608764133
transform 1 0 6808 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1608764133
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608764133
transform 1 0 4876 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608764133
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1608764133
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608764133
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_36
timestamp 1608764133
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_40
timestamp 1608764133
transform 1 0 4784 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608764133
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1608764133
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608764133
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608764133
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608764133
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608764133
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608764133
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608764133
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608764133
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1608764133
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1608764133
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1608764133
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_131
timestamp 1608764133
transform 1 0 13156 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_143
timestamp 1608764133
transform 1 0 14260 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1608764133
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1608764133
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608764133
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1608764133
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1608764133
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1608764133
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_106
timestamp 1608764133
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1608764133
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1608764133
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1608764133
transform 1 0 9016 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1608764133
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__10__A
timestamp 1608764133
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__11__A
timestamp 1608764133
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1608764133
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_90
timestamp 1608764133
transform 1 0 9384 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_95
timestamp 1608764133
transform 1 0 9844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1608764133
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1608764133
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__04__A
timestamp 1608764133
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__05__A
timestamp 1608764133
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__06__A
timestamp 1608764133
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1608764133
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1608764133
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1608764133
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1608764133
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _02_
timestamp 1608764133
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1608764133
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608764133
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__02__A
timestamp 1608764133
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1608764133
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_46
timestamp 1608764133
transform 1 0 5336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1608764133
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 1608764133
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1608764133
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1608764133
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1608764133
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1608764133
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_34
timestamp 1608764133
transform 1 0 4232 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_41
timestamp 1608764133
transform 1 0 4876 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608764133
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608764133
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608764133
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608764133
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608764133
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608764133
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1608764133
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608764133
transform 1 0 13524 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_127
timestamp 1608764133
transform 1 0 12788 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_139
timestamp 1608764133
transform 1 0 13892 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1608764133
transform 1 0 12420 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608764133
transform 1 0 11040 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_112
timestamp 1608764133
transform 1 0 11408 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_120
timestamp 1608764133
transform 1 0 12144 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1608764133
transform 1 0 9936 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608764133
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1608764133
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1608764133
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_100
timestamp 1608764133
transform 1 0 10304 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1608764133
transform 1 0 7820 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1608764133
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_72
timestamp 1608764133
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_77
timestamp 1608764133
transform 1 0 8188 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1608764133
transform 1 0 5888 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_44
timestamp 1608764133
transform 1 0 5152 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608764133
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1608764133
transform 1 0 4784 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608764133
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608764133
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1608764133
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608764133
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608764133
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608764133
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608764133
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149
timestamp 1608764133
transform 1 0 14812 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1608764133
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1608764133
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1608764133
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1608764133
transform 1 0 13156 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1608764133
transform 1 0 13708 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608764133
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608764133
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608764133
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1608764133
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1608764133
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1608764133
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1608764133
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1608764133
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1608764133
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1608764133
transform 1 0 9016 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608764133
transform 1 0 10120 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1608764133
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1608764133
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1608764133
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1608764133
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1608764133
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1608764133
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1608764133
transform 1 0 7912 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__07__A
timestamp 1608764133
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1608764133
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1608764133
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1608764133
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1608764133
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1608764133
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_82
timestamp 1608764133
transform 1 0 8648 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1608764133
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608764133
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1608764133
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_42
timestamp 1608764133
transform 1 0 4968 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1608764133
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_54
timestamp 1608764133
transform 1 0 6072 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608764133
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1608764133
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608764133
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_39
timestamp 1608764133
transform 1 0 4692 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608764133
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608764133
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608764133
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608764133
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608764133
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1608764133
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608764133
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608764133
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608764133
transform 1 0 11500 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1608764133
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1608764133
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608764133
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608764133
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_93
timestamp 1608764133
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_103
timestamp 1608764133
transform 1 0 10580 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1608764133
transform 1 0 8096 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_66
timestamp 1608764133
transform 1 0 7176 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1608764133
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608764133
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1608764133
transform 1 0 6808 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608764133
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_56
timestamp 1608764133
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608764133
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608764133
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608764133
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608764133
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608764133
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608764133
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608764133
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608764133
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608764133
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608764133
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1608764133
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1608764133
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1608764133
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608764133
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1608764133
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608764133
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608764133
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1608764133
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608764133
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608764133
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608764133
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115
timestamp 1608764133
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608764133
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1608764133
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608764133
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1608764133
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608764133
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608764133
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_90
timestamp 1608764133
transform 1 0 9384 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_98
timestamp 1608764133
transform 1 0 10120 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_101
timestamp 1608764133
transform 1 0 10396 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1608764133
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1608764133
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608764133
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608764133
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_66
timestamp 1608764133
transform 1 0 7176 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1608764133
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_78
timestamp 1608764133
transform 1 0 8280 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608764133
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608764133
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608764133
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608764133
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51
timestamp 1608764133
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608764133
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1608764133
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608764133
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608764133
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608764133
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608764133
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608764133
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608764133
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608764133
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608764133
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608764133
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608764133
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1608764133
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 4 IO_ISOL_N
port 1 nsew
rlabel metal3 s 0 18232 800 18352 4 ccff_head
port 2 nsew
rlabel metal3 s 16200 12384 17000 12504 4 ccff_tail
port 3 nsew
rlabel metal2 s 8666 0 8722 800 4 chany_bottom_in[0]
port 4 nsew
rlabel metal2 s 12898 0 12954 800 4 chany_bottom_in[10]
port 5 nsew
rlabel metal2 s 13358 0 13414 800 4 chany_bottom_in[11]
port 6 nsew
rlabel metal2 s 13818 0 13874 800 4 chany_bottom_in[12]
port 7 nsew
rlabel metal2 s 14186 0 14242 800 4 chany_bottom_in[13]
port 8 nsew
rlabel metal2 s 14646 0 14702 800 4 chany_bottom_in[14]
port 9 nsew
rlabel metal2 s 15014 0 15070 800 4 chany_bottom_in[15]
port 10 nsew
rlabel metal2 s 15474 0 15530 800 4 chany_bottom_in[16]
port 11 nsew
rlabel metal2 s 15934 0 15990 800 4 chany_bottom_in[17]
port 12 nsew
rlabel metal2 s 16302 0 16358 800 4 chany_bottom_in[18]
port 13 nsew
rlabel metal2 s 16762 0 16818 800 4 chany_bottom_in[19]
port 14 nsew
rlabel metal2 s 9126 0 9182 800 4 chany_bottom_in[1]
port 15 nsew
rlabel metal2 s 9494 0 9550 800 4 chany_bottom_in[2]
port 16 nsew
rlabel metal2 s 9954 0 10010 800 4 chany_bottom_in[3]
port 17 nsew
rlabel metal2 s 10414 0 10470 800 4 chany_bottom_in[4]
port 18 nsew
rlabel metal2 s 10782 0 10838 800 4 chany_bottom_in[5]
port 19 nsew
rlabel metal2 s 11242 0 11298 800 4 chany_bottom_in[6]
port 20 nsew
rlabel metal2 s 11610 0 11666 800 4 chany_bottom_in[7]
port 21 nsew
rlabel metal2 s 12070 0 12126 800 4 chany_bottom_in[8]
port 22 nsew
rlabel metal2 s 12530 0 12586 800 4 chany_bottom_in[9]
port 23 nsew
rlabel metal2 s 202 0 258 800 4 chany_bottom_out[0]
port 24 nsew
rlabel metal2 s 4434 0 4490 800 4 chany_bottom_out[10]
port 25 nsew
rlabel metal2 s 4802 0 4858 800 4 chany_bottom_out[11]
port 26 nsew
rlabel metal2 s 5262 0 5318 800 4 chany_bottom_out[12]
port 27 nsew
rlabel metal2 s 5722 0 5778 800 4 chany_bottom_out[13]
port 28 nsew
rlabel metal2 s 6090 0 6146 800 4 chany_bottom_out[14]
port 29 nsew
rlabel metal2 s 6550 0 6606 800 4 chany_bottom_out[15]
port 30 nsew
rlabel metal2 s 7010 0 7066 800 4 chany_bottom_out[16]
port 31 nsew
rlabel metal2 s 7378 0 7434 800 4 chany_bottom_out[17]
port 32 nsew
rlabel metal2 s 7838 0 7894 800 4 chany_bottom_out[18]
port 33 nsew
rlabel metal2 s 8206 0 8262 800 4 chany_bottom_out[19]
port 34 nsew
rlabel metal2 s 570 0 626 800 4 chany_bottom_out[1]
port 35 nsew
rlabel metal2 s 1030 0 1086 800 4 chany_bottom_out[2]
port 36 nsew
rlabel metal2 s 1398 0 1454 800 4 chany_bottom_out[3]
port 37 nsew
rlabel metal2 s 1858 0 1914 800 4 chany_bottom_out[4]
port 38 nsew
rlabel metal2 s 2318 0 2374 800 4 chany_bottom_out[5]
port 39 nsew
rlabel metal2 s 2686 0 2742 800 4 chany_bottom_out[6]
port 40 nsew
rlabel metal2 s 3146 0 3202 800 4 chany_bottom_out[7]
port 41 nsew
rlabel metal2 s 3606 0 3662 800 4 chany_bottom_out[8]
port 42 nsew
rlabel metal2 s 3974 0 4030 800 4 chany_bottom_out[9]
port 43 nsew
rlabel metal2 s 8850 19200 8906 20000 4 chany_top_in[0]
port 44 nsew
rlabel metal2 s 12990 19200 13046 20000 4 chany_top_in[10]
port 45 nsew
rlabel metal2 s 13450 19200 13506 20000 4 chany_top_in[11]
port 46 nsew
rlabel metal2 s 13818 19200 13874 20000 4 chany_top_in[12]
port 47 nsew
rlabel metal2 s 14278 19200 14334 20000 4 chany_top_in[13]
port 48 nsew
rlabel metal2 s 14646 19200 14702 20000 4 chany_top_in[14]
port 49 nsew
rlabel metal2 s 15106 19200 15162 20000 4 chany_top_in[15]
port 50 nsew
rlabel metal2 s 15474 19200 15530 20000 4 chany_top_in[16]
port 51 nsew
rlabel metal2 s 15934 19200 15990 20000 4 chany_top_in[17]
port 52 nsew
rlabel metal2 s 16302 19200 16358 20000 4 chany_top_in[18]
port 53 nsew
rlabel metal2 s 16762 19200 16818 20000 4 chany_top_in[19]
port 54 nsew
rlabel metal2 s 9310 19200 9366 20000 4 chany_top_in[1]
port 55 nsew
rlabel metal2 s 9678 19200 9734 20000 4 chany_top_in[2]
port 56 nsew
rlabel metal2 s 10138 19200 10194 20000 4 chany_top_in[3]
port 57 nsew
rlabel metal2 s 10506 19200 10562 20000 4 chany_top_in[4]
port 58 nsew
rlabel metal2 s 10966 19200 11022 20000 4 chany_top_in[5]
port 59 nsew
rlabel metal2 s 11334 19200 11390 20000 4 chany_top_in[6]
port 60 nsew
rlabel metal2 s 11794 19200 11850 20000 4 chany_top_in[7]
port 61 nsew
rlabel metal2 s 12162 19200 12218 20000 4 chany_top_in[8]
port 62 nsew
rlabel metal2 s 12622 19200 12678 20000 4 chany_top_in[9]
port 63 nsew
rlabel metal2 s 570 19200 626 20000 4 chany_top_out[0]
port 64 nsew
rlabel metal2 s 4710 19200 4766 20000 4 chany_top_out[10]
port 65 nsew
rlabel metal2 s 5170 19200 5226 20000 4 chany_top_out[11]
port 66 nsew
rlabel metal2 s 5538 19200 5594 20000 4 chany_top_out[12]
port 67 nsew
rlabel metal2 s 5998 19200 6054 20000 4 chany_top_out[13]
port 68 nsew
rlabel metal2 s 6366 19200 6422 20000 4 chany_top_out[14]
port 69 nsew
rlabel metal2 s 6826 19200 6882 20000 4 chany_top_out[15]
port 70 nsew
rlabel metal2 s 7194 19200 7250 20000 4 chany_top_out[16]
port 71 nsew
rlabel metal2 s 7654 19200 7710 20000 4 chany_top_out[17]
port 72 nsew
rlabel metal2 s 8022 19200 8078 20000 4 chany_top_out[18]
port 73 nsew
rlabel metal2 s 8482 19200 8538 20000 4 chany_top_out[19]
port 74 nsew
rlabel metal2 s 1030 19200 1086 20000 4 chany_top_out[1]
port 75 nsew
rlabel metal2 s 1398 19200 1454 20000 4 chany_top_out[2]
port 76 nsew
rlabel metal2 s 1858 19200 1914 20000 4 chany_top_out[3]
port 77 nsew
rlabel metal2 s 2226 19200 2282 20000 4 chany_top_out[4]
port 78 nsew
rlabel metal2 s 2686 19200 2742 20000 4 chany_top_out[5]
port 79 nsew
rlabel metal2 s 3054 19200 3110 20000 4 chany_top_out[6]
port 80 nsew
rlabel metal2 s 3514 19200 3570 20000 4 chany_top_out[7]
port 81 nsew
rlabel metal2 s 3882 19200 3938 20000 4 chany_top_out[8]
port 82 nsew
rlabel metal2 s 4342 19200 4398 20000 4 chany_top_out[9]
port 83 nsew
rlabel metal3 s 0 8304 800 8424 4 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 84 nsew
rlabel metal3 s 0 11568 800 11688 4 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 85 nsew
rlabel metal3 s 0 14968 800 15088 4 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 86 nsew
rlabel metal3 s 0 4904 800 5024 4 left_grid_pin_0_
port 87 nsew
rlabel metal3 s 16200 7352 17000 7472 4 prog_clk_0_E_in
port 88 nsew
rlabel metal3 s 0 1640 800 1760 4 right_width_0_height_0__pin_0_
port 89 nsew
rlabel metal3 s 16200 2456 17000 2576 4 right_width_0_height_0__pin_1_lower
port 90 nsew
rlabel metal3 s 16200 17416 17000 17536 4 right_width_0_height_0__pin_1_upper
port 91 nsew
rlabel metal4 s 3409 2128 3729 17456 4 VPWR
port 92 nsew
rlabel metal4 s 5875 2128 6195 17456 4 VGND
port 93 nsew
<< properties >>
string FIXED_BBOX 0 0 17000 20000
string GDS_FILE /ef/openfpga/openlane/runs/cby_0__1_/results/magic/cby_0__1_.gds
string GDS_END 456698
string GDS_START 101802
<< end >>
