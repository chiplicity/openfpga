magic
tech EFS8A
magscale 1 2
timestamp 1604431007
<< viali >>
rect 23949 19231 23983 19265
rect 24593 19231 24627 19265
rect 24133 19095 24167 19129
rect 16773 18891 16807 18925
rect 20821 18891 20855 18925
rect 8852 18823 8886 18857
rect 8585 18755 8619 18789
rect 15660 18755 15694 18789
rect 20637 18755 20671 18789
rect 23949 18755 23983 18789
rect 25053 18755 25087 18789
rect 15393 18687 15427 18721
rect 9965 18551 9999 18585
rect 24133 18551 24167 18585
rect 25237 18551 25271 18585
rect 8677 18347 8711 18381
rect 23857 18347 23891 18381
rect 25053 18347 25087 18381
rect 8953 18279 8987 18313
rect 15485 18143 15519 18177
rect 23949 18143 23983 18177
rect 24501 18143 24535 18177
rect 15853 18075 15887 18109
rect 20637 18007 20671 18041
rect 24133 18007 24167 18041
rect 23949 17667 23983 17701
rect 24133 17463 24167 17497
rect 18061 17259 18095 17293
rect 23949 17259 23983 17293
rect 17969 17123 18003 17157
rect 18705 17123 18739 17157
rect 18521 16987 18555 17021
rect 17509 16919 17543 16953
rect 18429 16919 18463 16953
rect 14473 16715 14507 16749
rect 18337 16715 18371 16749
rect 13093 16579 13127 16613
rect 13360 16579 13394 16613
rect 7021 16171 7055 16205
rect 13093 16171 13127 16205
rect 24501 16171 24535 16205
rect 7113 16035 7147 16069
rect 23949 15967 23983 16001
rect 7358 15899 7392 15933
rect 8493 15831 8527 15865
rect 13461 15831 13495 15865
rect 24133 15831 24167 15865
rect 7205 15627 7239 15661
rect 19073 15287 19107 15321
rect 18981 15083 19015 15117
rect 18797 14947 18831 14981
rect 19533 14947 19567 14981
rect 19349 14879 19383 14913
rect 19441 14743 19475 14777
rect 19073 14539 19107 14573
rect 19441 14539 19475 14573
rect 19809 14539 19843 14573
rect 23949 14403 23983 14437
rect 19901 14335 19935 14369
rect 19993 14335 20027 14369
rect 24133 14199 24167 14233
rect 19533 13995 19567 14029
rect 20177 13995 20211 14029
rect 24041 13995 24075 14029
rect 19809 13791 19843 13825
rect 13553 13451 13587 13485
rect 19165 13451 19199 13485
rect 1409 13315 1443 13349
rect 13921 13315 13955 13349
rect 19533 13315 19567 13349
rect 14013 13247 14047 13281
rect 14105 13247 14139 13281
rect 19625 13247 19659 13281
rect 19809 13247 19843 13281
rect 1593 13111 1627 13145
rect 13645 12907 13679 12941
rect 19993 12907 20027 12941
rect 19625 12771 19659 12805
rect 20913 12771 20947 12805
rect 1409 12703 1443 12737
rect 1961 12703 1995 12737
rect 19165 12703 19199 12737
rect 14289 12635 14323 12669
rect 1593 12567 1627 12601
rect 13921 12567 13955 12601
rect 1593 12363 1627 12397
rect 8401 12363 8435 12397
rect 13093 12363 13127 12397
rect 8309 12227 8343 12261
rect 13461 12227 13495 12261
rect 8493 12159 8527 12193
rect 13553 12159 13587 12193
rect 13645 12159 13679 12193
rect 7941 12091 7975 12125
rect 12173 12023 12207 12057
rect 8033 11819 8067 11853
rect 11989 11819 12023 11853
rect 12173 11819 12207 11853
rect 13921 11819 13955 11853
rect 24501 11819 24535 11853
rect 13185 11751 13219 11785
rect 12725 11683 12759 11717
rect 13553 11683 13587 11717
rect 1409 11615 1443 11649
rect 1961 11615 1995 11649
rect 12633 11615 12667 11649
rect 23949 11615 23983 11649
rect 1593 11479 1627 11513
rect 8309 11479 8343 11513
rect 8677 11479 8711 11513
rect 12541 11479 12575 11513
rect 24133 11479 24167 11513
rect 7757 11275 7791 11309
rect 12173 11275 12207 11309
rect 8125 11207 8159 11241
rect 1409 11139 1443 11173
rect 23949 11139 23983 11173
rect 8217 11071 8251 11105
rect 8309 11071 8343 11105
rect 1593 11003 1627 11037
rect 24133 11003 24167 11037
rect 2053 10731 2087 10765
rect 2421 10731 2455 10765
rect 7113 10731 7147 10765
rect 7941 10731 7975 10765
rect 8953 10731 8987 10765
rect 23949 10731 23983 10765
rect 8585 10595 8619 10629
rect 1409 10527 1443 10561
rect 8309 10459 8343 10493
rect 1593 10391 1627 10425
rect 7389 10391 7423 10425
rect 7849 10391 7883 10425
rect 8401 10391 8435 10425
rect 8033 10187 8067 10221
rect 8401 10187 8435 10221
rect 1409 10051 1443 10085
rect 1593 9847 1627 9881
rect 2053 9643 2087 9677
rect 2421 9575 2455 9609
rect 1409 9439 1443 9473
rect 23949 9439 23983 9473
rect 24501 9439 24535 9473
rect 1593 9303 1627 9337
rect 24133 9303 24167 9337
rect 1409 8963 1443 8997
rect 23949 8963 23983 8997
rect 1593 8759 1627 8793
rect 24133 8759 24167 8793
rect 1593 8555 1627 8589
rect 23765 8555 23799 8589
rect 24501 8555 24535 8589
rect 24133 8487 24167 8521
rect 23949 8351 23983 8385
rect 24133 8011 24167 8045
rect 23949 7875 23983 7909
rect 22477 7467 22511 7501
rect 22937 7467 22971 7501
rect 23949 7467 23983 7501
rect 18613 7399 18647 7433
rect 13093 7263 13127 7297
rect 13645 7263 13679 7297
rect 18429 7263 18463 7297
rect 18981 7263 19015 7297
rect 22293 7263 22327 7297
rect 13277 7127 13311 7161
rect 14749 6787 14783 6821
rect 23949 6787 23983 6821
rect 14933 6651 14967 6685
rect 24133 6651 24167 6685
rect 14749 6379 14783 6413
rect 24041 6379 24075 6413
rect 13093 5835 13127 5869
rect 4169 5699 4203 5733
rect 12909 5699 12943 5733
rect 4353 5563 4387 5597
rect 4261 5291 4295 5325
rect 13645 5291 13679 5325
rect 24593 5291 24627 5325
rect 12633 5087 12667 5121
rect 13185 5087 13219 5121
rect 23949 5087 23983 5121
rect 12817 4951 12851 4985
rect 24133 4951 24167 4985
rect 15577 4611 15611 4645
rect 20453 4611 20487 4645
rect 15761 4475 15795 4509
rect 20637 4475 20671 4509
rect 15577 4203 15611 4237
rect 20453 4203 20487 4237
rect 21465 4067 21499 4101
rect 20913 3999 20947 4033
rect 23949 3999 23983 4033
rect 24501 3999 24535 4033
rect 21097 3863 21131 3897
rect 24133 3863 24167 3897
rect 23949 3523 23983 3557
rect 24133 3387 24167 3421
rect 1961 3115 1995 3149
rect 23857 3115 23891 3149
rect 1409 2911 1443 2945
rect 23949 2911 23983 2945
rect 24501 2911 24535 2945
rect 1593 2775 1627 2809
rect 24133 2775 24167 2809
rect 24225 2571 24259 2605
rect 1409 2435 1443 2469
rect 24041 2435 24075 2469
rect 24593 2435 24627 2469
rect 25145 2435 25179 2469
rect 25697 2435 25731 2469
rect 2053 2367 2087 2401
rect 1593 2231 1627 2265
rect 25329 2231 25363 2265
<< metal1 >>
rect 1104 21756 28888 21778
rect 1104 21704 5982 21756
rect 6034 21704 6046 21756
rect 6098 21704 6110 21756
rect 6162 21704 6174 21756
rect 6226 21704 15982 21756
rect 16034 21704 16046 21756
rect 16098 21704 16110 21756
rect 16162 21704 16174 21756
rect 16226 21704 25982 21756
rect 26034 21704 26046 21756
rect 26098 21704 26110 21756
rect 26162 21704 26174 21756
rect 26226 21704 28888 21756
rect 1104 21682 28888 21704
rect 1104 21212 28888 21234
rect 1104 21160 10982 21212
rect 11034 21160 11046 21212
rect 11098 21160 11110 21212
rect 11162 21160 11174 21212
rect 11226 21160 20982 21212
rect 21034 21160 21046 21212
rect 21098 21160 21110 21212
rect 21162 21160 21174 21212
rect 21226 21160 28888 21212
rect 1104 21138 28888 21160
rect 3418 20718 3424 20770
rect 3476 20758 3482 20770
rect 19426 20758 19432 20770
rect 3476 20730 19432 20758
rect 3476 20718 3482 20730
rect 19426 20718 19432 20730
rect 19484 20718 19490 20770
rect 19610 20718 19616 20770
rect 19668 20758 19674 20770
rect 24854 20758 24860 20770
rect 19668 20730 24860 20758
rect 19668 20718 19674 20730
rect 24854 20718 24860 20730
rect 24912 20718 24918 20770
rect 1104 20668 28888 20690
rect 1104 20616 5982 20668
rect 6034 20616 6046 20668
rect 6098 20616 6110 20668
rect 6162 20616 6174 20668
rect 6226 20616 15982 20668
rect 16034 20616 16046 20668
rect 16098 20616 16110 20668
rect 16162 20616 16174 20668
rect 16226 20616 25982 20668
rect 26034 20616 26046 20668
rect 26098 20616 26110 20668
rect 26162 20616 26174 20668
rect 26226 20616 28888 20668
rect 1104 20594 28888 20616
rect 1104 20124 28888 20146
rect 1104 20072 10982 20124
rect 11034 20072 11046 20124
rect 11098 20072 11110 20124
rect 11162 20072 11174 20124
rect 11226 20072 20982 20124
rect 21034 20072 21046 20124
rect 21098 20072 21110 20124
rect 21162 20072 21174 20124
rect 21226 20072 28888 20124
rect 1104 20050 28888 20072
rect 1104 19580 28888 19602
rect 1104 19528 5982 19580
rect 6034 19528 6046 19580
rect 6098 19528 6110 19580
rect 6162 19528 6174 19580
rect 6226 19528 15982 19580
rect 16034 19528 16046 19580
rect 16098 19528 16110 19580
rect 16162 19528 16174 19580
rect 16226 19528 25982 19580
rect 26034 19528 26046 19580
rect 26098 19528 26110 19580
rect 26162 19528 26174 19580
rect 26226 19528 28888 19580
rect 1104 19506 28888 19528
rect 23937 19265 23995 19271
rect 23937 19231 23949 19265
rect 23983 19262 23995 19265
rect 24581 19265 24639 19271
rect 24581 19262 24593 19265
rect 23983 19234 24593 19262
rect 23983 19231 23995 19234
rect 23937 19225 23995 19231
rect 24581 19231 24593 19234
rect 24627 19262 24639 19265
rect 24762 19262 24768 19274
rect 24627 19234 24768 19262
rect 24627 19231 24639 19234
rect 24581 19225 24639 19231
rect 24762 19222 24768 19234
rect 24820 19222 24826 19274
rect 23474 19086 23480 19138
rect 23532 19126 23538 19138
rect 24121 19129 24179 19135
rect 24121 19126 24133 19129
rect 23532 19098 24133 19126
rect 23532 19086 23538 19098
rect 24121 19095 24133 19098
rect 24167 19095 24179 19129
rect 24121 19089 24179 19095
rect 1104 19036 28888 19058
rect 1104 18984 10982 19036
rect 11034 18984 11046 19036
rect 11098 18984 11110 19036
rect 11162 18984 11174 19036
rect 11226 18984 20982 19036
rect 21034 18984 21046 19036
rect 21098 18984 21110 19036
rect 21162 18984 21174 19036
rect 21226 18984 28888 19036
rect 1104 18962 28888 18984
rect 16758 18922 16764 18934
rect 16719 18894 16764 18922
rect 16758 18882 16764 18894
rect 16816 18882 16822 18934
rect 20806 18922 20812 18934
rect 20767 18894 20812 18922
rect 20806 18882 20812 18894
rect 20864 18882 20870 18934
rect 3142 18814 3148 18866
rect 3200 18854 3206 18866
rect 3694 18854 3700 18866
rect 3200 18826 3700 18854
rect 3200 18814 3206 18826
rect 3694 18814 3700 18826
rect 3752 18814 3758 18866
rect 8846 18863 8852 18866
rect 8840 18854 8852 18863
rect 8807 18826 8852 18854
rect 8840 18817 8852 18826
rect 8846 18814 8852 18817
rect 8904 18814 8910 18866
rect 8570 18786 8576 18798
rect 8531 18758 8576 18786
rect 8570 18746 8576 18758
rect 8628 18746 8634 18798
rect 15654 18795 15660 18798
rect 15648 18786 15660 18795
rect 15615 18758 15660 18786
rect 15648 18749 15660 18758
rect 15654 18746 15660 18749
rect 15712 18746 15718 18798
rect 20622 18786 20628 18798
rect 20583 18758 20628 18786
rect 20622 18746 20628 18758
rect 20680 18746 20686 18798
rect 23934 18786 23940 18798
rect 23895 18758 23940 18786
rect 23934 18746 23940 18758
rect 23992 18746 23998 18798
rect 25038 18786 25044 18798
rect 24999 18758 25044 18786
rect 25038 18746 25044 18758
rect 25096 18746 25102 18798
rect 15378 18718 15384 18730
rect 15339 18690 15384 18718
rect 15378 18678 15384 18690
rect 15436 18678 15442 18730
rect 9950 18582 9956 18594
rect 9911 18554 9956 18582
rect 9950 18542 9956 18554
rect 10008 18542 10014 18594
rect 24118 18582 24124 18594
rect 24079 18554 24124 18582
rect 24118 18542 24124 18554
rect 24176 18542 24182 18594
rect 25222 18582 25228 18594
rect 25183 18554 25228 18582
rect 25222 18542 25228 18554
rect 25280 18542 25286 18594
rect 1104 18492 28888 18514
rect 1104 18440 5982 18492
rect 6034 18440 6046 18492
rect 6098 18440 6110 18492
rect 6162 18440 6174 18492
rect 6226 18440 15982 18492
rect 16034 18440 16046 18492
rect 16098 18440 16110 18492
rect 16162 18440 16174 18492
rect 16226 18440 25982 18492
rect 26034 18440 26046 18492
rect 26098 18440 26110 18492
rect 26162 18440 26174 18492
rect 26226 18440 28888 18492
rect 1104 18418 28888 18440
rect 8665 18381 8723 18387
rect 8665 18347 8677 18381
rect 8711 18378 8723 18381
rect 8846 18378 8852 18390
rect 8711 18350 8852 18378
rect 8711 18347 8723 18350
rect 8665 18341 8723 18347
rect 8846 18338 8852 18350
rect 8904 18338 8910 18390
rect 23845 18381 23903 18387
rect 23845 18347 23857 18381
rect 23891 18378 23903 18381
rect 23934 18378 23940 18390
rect 23891 18350 23940 18378
rect 23891 18347 23903 18350
rect 23845 18341 23903 18347
rect 23934 18338 23940 18350
rect 23992 18338 23998 18390
rect 25038 18378 25044 18390
rect 24999 18350 25044 18378
rect 25038 18338 25044 18350
rect 25096 18338 25102 18390
rect 8570 18270 8576 18322
rect 8628 18310 8634 18322
rect 8941 18313 8999 18319
rect 8941 18310 8953 18313
rect 8628 18282 8953 18310
rect 8628 18270 8634 18282
rect 8941 18279 8953 18282
rect 8987 18279 8999 18313
rect 8941 18273 8999 18279
rect 15378 18134 15384 18186
rect 15436 18174 15442 18186
rect 15473 18177 15531 18183
rect 15473 18174 15485 18177
rect 15436 18146 15485 18174
rect 15436 18134 15442 18146
rect 15473 18143 15485 18146
rect 15519 18143 15531 18177
rect 23934 18174 23940 18186
rect 23895 18146 23940 18174
rect 15473 18137 15531 18143
rect 23934 18134 23940 18146
rect 23992 18174 23998 18186
rect 24489 18177 24547 18183
rect 24489 18174 24501 18177
rect 23992 18146 24501 18174
rect 23992 18134 23998 18146
rect 24489 18143 24501 18146
rect 24535 18143 24547 18177
rect 24489 18137 24547 18143
rect 15194 18066 15200 18118
rect 15252 18106 15258 18118
rect 15654 18106 15660 18118
rect 15252 18078 15660 18106
rect 15252 18066 15258 18078
rect 15654 18066 15660 18078
rect 15712 18106 15718 18118
rect 15841 18109 15899 18115
rect 15841 18106 15853 18109
rect 15712 18078 15853 18106
rect 15712 18066 15718 18078
rect 15841 18075 15853 18078
rect 15887 18075 15899 18109
rect 15841 18069 15899 18075
rect 19334 17998 19340 18050
rect 19392 18038 19398 18050
rect 20622 18038 20628 18050
rect 19392 18010 20628 18038
rect 19392 17998 19398 18010
rect 20622 17998 20628 18010
rect 20680 17998 20686 18050
rect 24121 18041 24179 18047
rect 24121 18007 24133 18041
rect 24167 18038 24179 18041
rect 24302 18038 24308 18050
rect 24167 18010 24308 18038
rect 24167 18007 24179 18010
rect 24121 18001 24179 18007
rect 24302 17998 24308 18010
rect 24360 17998 24366 18050
rect 1104 17948 28888 17970
rect 1104 17896 10982 17948
rect 11034 17896 11046 17948
rect 11098 17896 11110 17948
rect 11162 17896 11174 17948
rect 11226 17896 20982 17948
rect 21034 17896 21046 17948
rect 21098 17896 21110 17948
rect 21162 17896 21174 17948
rect 21226 17896 28888 17948
rect 1104 17874 28888 17896
rect 23934 17698 23940 17710
rect 23895 17670 23940 17698
rect 23934 17658 23940 17670
rect 23992 17658 23998 17710
rect 24121 17497 24179 17503
rect 24121 17463 24133 17497
rect 24167 17494 24179 17497
rect 24210 17494 24216 17506
rect 24167 17466 24216 17494
rect 24167 17463 24179 17466
rect 24121 17457 24179 17463
rect 24210 17454 24216 17466
rect 24268 17454 24274 17506
rect 1104 17404 28888 17426
rect 1104 17352 5982 17404
rect 6034 17352 6046 17404
rect 6098 17352 6110 17404
rect 6162 17352 6174 17404
rect 6226 17352 15982 17404
rect 16034 17352 16046 17404
rect 16098 17352 16110 17404
rect 16162 17352 16174 17404
rect 16226 17352 25982 17404
rect 26034 17352 26046 17404
rect 26098 17352 26110 17404
rect 26162 17352 26174 17404
rect 26226 17352 28888 17404
rect 1104 17330 28888 17352
rect 18049 17293 18107 17299
rect 18049 17259 18061 17293
rect 18095 17290 18107 17293
rect 19242 17290 19248 17302
rect 18095 17262 19248 17290
rect 18095 17259 18107 17262
rect 18049 17253 18107 17259
rect 19242 17250 19248 17262
rect 19300 17250 19306 17302
rect 23934 17290 23940 17302
rect 23895 17262 23940 17290
rect 23934 17250 23940 17262
rect 23992 17250 23998 17302
rect 17957 17157 18015 17163
rect 17957 17123 17969 17157
rect 18003 17154 18015 17157
rect 18690 17154 18696 17166
rect 18003 17126 18696 17154
rect 18003 17123 18015 17126
rect 17957 17117 18015 17123
rect 18690 17114 18696 17126
rect 18748 17114 18754 17166
rect 18509 17021 18567 17027
rect 18509 17018 18521 17021
rect 17512 16990 18521 17018
rect 17512 16962 17540 16990
rect 18509 16987 18521 16990
rect 18555 16987 18567 17021
rect 18509 16981 18567 16987
rect 17494 16950 17500 16962
rect 17455 16922 17500 16950
rect 17494 16910 17500 16922
rect 17552 16910 17558 16962
rect 18322 16910 18328 16962
rect 18380 16950 18386 16962
rect 18417 16953 18475 16959
rect 18417 16950 18429 16953
rect 18380 16922 18429 16950
rect 18380 16910 18386 16922
rect 18417 16919 18429 16922
rect 18463 16919 18475 16953
rect 18417 16913 18475 16919
rect 1104 16860 28888 16882
rect 1104 16808 10982 16860
rect 11034 16808 11046 16860
rect 11098 16808 11110 16860
rect 11162 16808 11174 16860
rect 11226 16808 20982 16860
rect 21034 16808 21046 16860
rect 21098 16808 21110 16860
rect 21162 16808 21174 16860
rect 21226 16808 28888 16860
rect 1104 16786 28888 16808
rect 14090 16706 14096 16758
rect 14148 16746 14154 16758
rect 14461 16749 14519 16755
rect 14461 16746 14473 16749
rect 14148 16718 14473 16746
rect 14148 16706 14154 16718
rect 14461 16715 14473 16718
rect 14507 16746 14519 16749
rect 15194 16746 15200 16758
rect 14507 16718 15200 16746
rect 14507 16715 14519 16718
rect 14461 16709 14519 16715
rect 15194 16706 15200 16718
rect 15252 16706 15258 16758
rect 18322 16746 18328 16758
rect 18283 16718 18328 16746
rect 18322 16706 18328 16718
rect 18380 16706 18386 16758
rect 13078 16610 13084 16622
rect 13039 16582 13084 16610
rect 13078 16570 13084 16582
rect 13136 16570 13142 16622
rect 13348 16613 13406 16619
rect 13348 16579 13360 16613
rect 13394 16610 13406 16613
rect 13630 16610 13636 16622
rect 13394 16582 13636 16610
rect 13394 16579 13406 16582
rect 13348 16573 13406 16579
rect 13630 16570 13636 16582
rect 13688 16570 13694 16622
rect 1104 16316 28888 16338
rect 1104 16264 5982 16316
rect 6034 16264 6046 16316
rect 6098 16264 6110 16316
rect 6162 16264 6174 16316
rect 6226 16264 15982 16316
rect 16034 16264 16046 16316
rect 16098 16264 16110 16316
rect 16162 16264 16174 16316
rect 16226 16264 25982 16316
rect 26034 16264 26046 16316
rect 26098 16264 26110 16316
rect 26162 16264 26174 16316
rect 26226 16264 28888 16316
rect 1104 16242 28888 16264
rect 7006 16202 7012 16214
rect 6967 16174 7012 16202
rect 7006 16162 7012 16174
rect 7064 16162 7070 16214
rect 13078 16202 13084 16214
rect 13039 16174 13084 16202
rect 13078 16162 13084 16174
rect 13136 16162 13142 16214
rect 24486 16202 24492 16214
rect 24447 16174 24492 16202
rect 24486 16162 24492 16174
rect 24544 16162 24550 16214
rect 7024 16066 7052 16162
rect 7101 16069 7159 16075
rect 7101 16066 7113 16069
rect 7024 16038 7113 16066
rect 7101 16035 7113 16038
rect 7147 16035 7159 16069
rect 7101 16029 7159 16035
rect 23937 16001 23995 16007
rect 23937 15967 23949 16001
rect 23983 15998 23995 16001
rect 24486 15998 24492 16010
rect 23983 15970 24492 15998
rect 23983 15967 23995 15970
rect 23937 15961 23995 15967
rect 24486 15958 24492 15970
rect 24544 15958 24550 16010
rect 7190 15890 7196 15942
rect 7248 15930 7254 15942
rect 7346 15933 7404 15939
rect 7346 15930 7358 15933
rect 7248 15902 7358 15930
rect 7248 15890 7254 15902
rect 7346 15899 7358 15902
rect 7392 15899 7404 15933
rect 7346 15893 7404 15899
rect 8478 15862 8484 15874
rect 8439 15834 8484 15862
rect 8478 15822 8484 15834
rect 8536 15822 8542 15874
rect 13446 15862 13452 15874
rect 13407 15834 13452 15862
rect 13446 15822 13452 15834
rect 13504 15862 13510 15874
rect 13630 15862 13636 15874
rect 13504 15834 13636 15862
rect 13504 15822 13510 15834
rect 13630 15822 13636 15834
rect 13688 15822 13694 15874
rect 23658 15822 23664 15874
rect 23716 15862 23722 15874
rect 24121 15865 24179 15871
rect 24121 15862 24133 15865
rect 23716 15834 24133 15862
rect 23716 15822 23722 15834
rect 24121 15831 24133 15834
rect 24167 15831 24179 15865
rect 24121 15825 24179 15831
rect 1104 15772 28888 15794
rect 1104 15720 10982 15772
rect 11034 15720 11046 15772
rect 11098 15720 11110 15772
rect 11162 15720 11174 15772
rect 11226 15720 20982 15772
rect 21034 15720 21046 15772
rect 21098 15720 21110 15772
rect 21162 15720 21174 15772
rect 21226 15720 28888 15772
rect 1104 15698 28888 15720
rect 7190 15658 7196 15670
rect 7151 15630 7196 15658
rect 7190 15618 7196 15630
rect 7248 15618 7254 15670
rect 19061 15321 19119 15327
rect 19061 15287 19073 15321
rect 19107 15318 19119 15321
rect 19242 15318 19248 15330
rect 19107 15290 19248 15318
rect 19107 15287 19119 15290
rect 19061 15281 19119 15287
rect 19242 15278 19248 15290
rect 19300 15278 19306 15330
rect 1104 15228 28888 15250
rect 1104 15176 5982 15228
rect 6034 15176 6046 15228
rect 6098 15176 6110 15228
rect 6162 15176 6174 15228
rect 6226 15176 15982 15228
rect 16034 15176 16046 15228
rect 16098 15176 16110 15228
rect 16162 15176 16174 15228
rect 16226 15176 25982 15228
rect 26034 15176 26046 15228
rect 26098 15176 26110 15228
rect 26162 15176 26174 15228
rect 26226 15176 28888 15228
rect 1104 15154 28888 15176
rect 18322 15074 18328 15126
rect 18380 15114 18386 15126
rect 18969 15117 19027 15123
rect 18969 15114 18981 15117
rect 18380 15086 18981 15114
rect 18380 15074 18386 15086
rect 18969 15083 18981 15086
rect 19015 15083 19027 15117
rect 18969 15077 19027 15083
rect 18782 14978 18788 14990
rect 18743 14950 18788 14978
rect 18782 14938 18788 14950
rect 18840 14978 18846 14990
rect 19521 14981 19579 14987
rect 19521 14978 19533 14981
rect 18840 14950 19533 14978
rect 18840 14938 18846 14950
rect 19521 14947 19533 14950
rect 19567 14947 19579 14981
rect 19521 14941 19579 14947
rect 19334 14910 19340 14922
rect 19295 14882 19340 14910
rect 19334 14870 19340 14882
rect 19392 14870 19398 14922
rect 19426 14734 19432 14786
rect 19484 14774 19490 14786
rect 19484 14746 19529 14774
rect 19484 14734 19490 14746
rect 1104 14684 28888 14706
rect 1104 14632 10982 14684
rect 11034 14632 11046 14684
rect 11098 14632 11110 14684
rect 11162 14632 11174 14684
rect 11226 14632 20982 14684
rect 21034 14632 21046 14684
rect 21098 14632 21110 14684
rect 21162 14632 21174 14684
rect 21226 14632 28888 14684
rect 1104 14610 28888 14632
rect 19061 14573 19119 14579
rect 19061 14539 19073 14573
rect 19107 14570 19119 14573
rect 19426 14570 19432 14582
rect 19107 14542 19432 14570
rect 19107 14539 19119 14542
rect 19061 14533 19119 14539
rect 19426 14530 19432 14542
rect 19484 14530 19490 14582
rect 19518 14530 19524 14582
rect 19576 14570 19582 14582
rect 19797 14573 19855 14579
rect 19797 14570 19809 14573
rect 19576 14542 19809 14570
rect 19576 14530 19582 14542
rect 19797 14539 19809 14542
rect 19843 14539 19855 14573
rect 19797 14533 19855 14539
rect 23937 14437 23995 14443
rect 23937 14403 23949 14437
rect 23983 14434 23995 14437
rect 24026 14434 24032 14446
rect 23983 14406 24032 14434
rect 23983 14403 23995 14406
rect 23937 14397 23995 14403
rect 24026 14394 24032 14406
rect 24084 14394 24090 14446
rect 19702 14326 19708 14378
rect 19760 14366 19766 14378
rect 19886 14366 19892 14378
rect 19760 14338 19892 14366
rect 19760 14326 19766 14338
rect 19886 14326 19892 14338
rect 19944 14326 19950 14378
rect 19978 14326 19984 14378
rect 20036 14366 20042 14378
rect 20036 14338 20081 14366
rect 20036 14326 20042 14338
rect 23566 14190 23572 14242
rect 23624 14230 23630 14242
rect 24121 14233 24179 14239
rect 24121 14230 24133 14233
rect 23624 14202 24133 14230
rect 23624 14190 23630 14202
rect 24121 14199 24133 14202
rect 24167 14199 24179 14233
rect 24121 14193 24179 14199
rect 1104 14140 28888 14162
rect 1104 14088 5982 14140
rect 6034 14088 6046 14140
rect 6098 14088 6110 14140
rect 6162 14088 6174 14140
rect 6226 14088 15982 14140
rect 16034 14088 16046 14140
rect 16098 14088 16110 14140
rect 16162 14088 16174 14140
rect 16226 14088 25982 14140
rect 26034 14088 26046 14140
rect 26098 14088 26110 14140
rect 26162 14088 26174 14140
rect 26226 14088 28888 14140
rect 1104 14066 28888 14088
rect 19518 14026 19524 14038
rect 19479 13998 19524 14026
rect 19518 13986 19524 13998
rect 19576 13986 19582 14038
rect 19978 13986 19984 14038
rect 20036 14026 20042 14038
rect 20165 14029 20223 14035
rect 20165 14026 20177 14029
rect 20036 13998 20177 14026
rect 20036 13986 20042 13998
rect 20165 13995 20177 13998
rect 20211 13995 20223 14029
rect 24026 14026 24032 14038
rect 23987 13998 24032 14026
rect 20165 13989 20223 13995
rect 24026 13986 24032 13998
rect 24084 13986 24090 14038
rect 19702 13782 19708 13834
rect 19760 13822 19766 13834
rect 19797 13825 19855 13831
rect 19797 13822 19809 13825
rect 19760 13794 19809 13822
rect 19760 13782 19766 13794
rect 19797 13791 19809 13794
rect 19843 13791 19855 13825
rect 19797 13785 19855 13791
rect 1104 13596 28888 13618
rect 1104 13544 10982 13596
rect 11034 13544 11046 13596
rect 11098 13544 11110 13596
rect 11162 13544 11174 13596
rect 11226 13544 20982 13596
rect 21034 13544 21046 13596
rect 21098 13544 21110 13596
rect 21162 13544 21174 13596
rect 21226 13544 28888 13596
rect 1104 13522 28888 13544
rect 13538 13482 13544 13494
rect 13499 13454 13544 13482
rect 13538 13442 13544 13454
rect 13596 13442 13602 13494
rect 19153 13485 19211 13491
rect 19153 13451 19165 13485
rect 19199 13482 19211 13485
rect 19242 13482 19248 13494
rect 19199 13454 19248 13482
rect 19199 13451 19211 13454
rect 19153 13445 19211 13451
rect 19242 13442 19248 13454
rect 19300 13442 19306 13494
rect 1397 13349 1455 13355
rect 1397 13315 1409 13349
rect 1443 13346 1455 13349
rect 1486 13346 1492 13358
rect 1443 13318 1492 13346
rect 1443 13315 1455 13318
rect 1397 13309 1455 13315
rect 1486 13306 1492 13318
rect 1544 13306 1550 13358
rect 3234 13306 3240 13358
rect 3292 13346 3298 13358
rect 3878 13346 3884 13358
rect 3292 13318 3884 13346
rect 3292 13306 3298 13318
rect 3878 13306 3884 13318
rect 3936 13306 3942 13358
rect 13814 13306 13820 13358
rect 13872 13346 13878 13358
rect 13909 13349 13967 13355
rect 13909 13346 13921 13349
rect 13872 13318 13921 13346
rect 13872 13306 13878 13318
rect 13909 13315 13921 13318
rect 13955 13315 13967 13349
rect 19518 13346 19524 13358
rect 19479 13318 19524 13346
rect 13909 13309 13967 13315
rect 19518 13306 19524 13318
rect 19576 13306 19582 13358
rect 14001 13281 14059 13287
rect 14001 13247 14013 13281
rect 14047 13247 14059 13281
rect 14001 13241 14059 13247
rect 13906 13170 13912 13222
rect 13964 13210 13970 13222
rect 14016 13210 14044 13241
rect 14090 13238 14096 13290
rect 14148 13278 14154 13290
rect 14148 13250 14193 13278
rect 14148 13238 14154 13250
rect 19150 13238 19156 13290
rect 19208 13278 19214 13290
rect 19610 13278 19616 13290
rect 19208 13250 19616 13278
rect 19208 13238 19214 13250
rect 19610 13238 19616 13250
rect 19668 13238 19674 13290
rect 19797 13281 19855 13287
rect 19797 13247 19809 13281
rect 19843 13278 19855 13281
rect 19978 13278 19984 13290
rect 19843 13250 19984 13278
rect 19843 13247 19855 13250
rect 19797 13241 19855 13247
rect 19978 13238 19984 13250
rect 20036 13238 20042 13290
rect 13964 13182 14044 13210
rect 13964 13170 13970 13182
rect 1581 13145 1639 13151
rect 1581 13111 1593 13145
rect 1627 13142 1639 13145
rect 1854 13142 1860 13154
rect 1627 13114 1860 13142
rect 1627 13111 1639 13114
rect 1581 13105 1639 13111
rect 1854 13102 1860 13114
rect 1912 13102 1918 13154
rect 1104 13052 28888 13074
rect 1104 13000 5982 13052
rect 6034 13000 6046 13052
rect 6098 13000 6110 13052
rect 6162 13000 6174 13052
rect 6226 13000 15982 13052
rect 16034 13000 16046 13052
rect 16098 13000 16110 13052
rect 16162 13000 16174 13052
rect 16226 13000 25982 13052
rect 26034 13000 26046 13052
rect 26098 13000 26110 13052
rect 26162 13000 26174 13052
rect 26226 13000 28888 13052
rect 1104 12978 28888 13000
rect 13633 12941 13691 12947
rect 13633 12907 13645 12941
rect 13679 12938 13691 12941
rect 14090 12938 14096 12950
rect 13679 12910 14096 12938
rect 13679 12907 13691 12910
rect 13633 12901 13691 12907
rect 14090 12898 14096 12910
rect 14148 12898 14154 12950
rect 19978 12938 19984 12950
rect 19939 12910 19984 12938
rect 19978 12898 19984 12910
rect 20036 12898 20042 12950
rect 19518 12762 19524 12814
rect 19576 12802 19582 12814
rect 19613 12805 19671 12811
rect 19613 12802 19625 12805
rect 19576 12774 19625 12802
rect 19576 12762 19582 12774
rect 19613 12771 19625 12774
rect 19659 12802 19671 12805
rect 20901 12805 20959 12811
rect 20901 12802 20913 12805
rect 19659 12774 20913 12802
rect 19659 12771 19671 12774
rect 19613 12765 19671 12771
rect 20901 12771 20913 12774
rect 20947 12771 20959 12805
rect 20901 12765 20959 12771
rect 1394 12734 1400 12746
rect 1355 12706 1400 12734
rect 1394 12694 1400 12706
rect 1452 12734 1458 12746
rect 1949 12737 2007 12743
rect 1949 12734 1961 12737
rect 1452 12706 1961 12734
rect 1452 12694 1458 12706
rect 1949 12703 1961 12706
rect 1995 12703 2007 12737
rect 19150 12734 19156 12746
rect 19111 12706 19156 12734
rect 1949 12697 2007 12703
rect 19150 12694 19156 12706
rect 19208 12694 19214 12746
rect 13814 12626 13820 12678
rect 13872 12666 13878 12678
rect 14277 12669 14335 12675
rect 14277 12666 14289 12669
rect 13872 12638 14289 12666
rect 13872 12626 13878 12638
rect 14277 12635 14289 12638
rect 14323 12635 14335 12669
rect 14277 12629 14335 12635
rect 1581 12601 1639 12607
rect 1581 12567 1593 12601
rect 1627 12598 1639 12601
rect 1670 12598 1676 12610
rect 1627 12570 1676 12598
rect 1627 12567 1639 12570
rect 1581 12561 1639 12567
rect 1670 12558 1676 12570
rect 1728 12558 1734 12610
rect 13906 12598 13912 12610
rect 13867 12570 13912 12598
rect 13906 12558 13912 12570
rect 13964 12558 13970 12610
rect 1104 12508 28888 12530
rect 1104 12456 10982 12508
rect 11034 12456 11046 12508
rect 11098 12456 11110 12508
rect 11162 12456 11174 12508
rect 11226 12456 20982 12508
rect 21034 12456 21046 12508
rect 21098 12456 21110 12508
rect 21162 12456 21174 12508
rect 21226 12456 28888 12508
rect 1104 12434 28888 12456
rect 1486 12354 1492 12406
rect 1544 12394 1550 12406
rect 1581 12397 1639 12403
rect 1581 12394 1593 12397
rect 1544 12366 1593 12394
rect 1544 12354 1550 12366
rect 1581 12363 1593 12366
rect 1627 12363 1639 12397
rect 1581 12357 1639 12363
rect 8294 12354 8300 12406
rect 8352 12394 8358 12406
rect 8389 12397 8447 12403
rect 8389 12394 8401 12397
rect 8352 12366 8401 12394
rect 8352 12354 8358 12366
rect 8389 12363 8401 12366
rect 8435 12363 8447 12397
rect 8389 12357 8447 12363
rect 13081 12397 13139 12403
rect 13081 12363 13093 12397
rect 13127 12394 13139 12397
rect 13722 12394 13728 12406
rect 13127 12366 13728 12394
rect 13127 12363 13139 12366
rect 13081 12357 13139 12363
rect 13722 12354 13728 12366
rect 13780 12354 13786 12406
rect 8297 12261 8355 12267
rect 8297 12227 8309 12261
rect 8343 12258 8355 12261
rect 8662 12258 8668 12270
rect 8343 12230 8668 12258
rect 8343 12227 8355 12230
rect 8297 12221 8355 12227
rect 8662 12218 8668 12230
rect 8720 12218 8726 12270
rect 13078 12218 13084 12270
rect 13136 12258 13142 12270
rect 13449 12261 13507 12267
rect 13449 12258 13461 12261
rect 13136 12230 13461 12258
rect 13136 12218 13142 12230
rect 13449 12227 13461 12230
rect 13495 12227 13507 12261
rect 13449 12221 13507 12227
rect 8478 12190 8484 12202
rect 8439 12162 8484 12190
rect 8478 12150 8484 12162
rect 8536 12150 8542 12202
rect 13538 12190 13544 12202
rect 13499 12162 13544 12190
rect 13538 12150 13544 12162
rect 13596 12150 13602 12202
rect 13633 12193 13691 12199
rect 13633 12159 13645 12193
rect 13679 12159 13691 12193
rect 13633 12153 13691 12159
rect 7926 12122 7932 12134
rect 7887 12094 7932 12122
rect 7926 12082 7932 12094
rect 7984 12082 7990 12134
rect 13446 12082 13452 12134
rect 13504 12122 13510 12134
rect 13648 12122 13676 12153
rect 13504 12094 13676 12122
rect 13504 12082 13510 12094
rect 12066 12014 12072 12066
rect 12124 12054 12130 12066
rect 12161 12057 12219 12063
rect 12161 12054 12173 12057
rect 12124 12026 12173 12054
rect 12124 12014 12130 12026
rect 12161 12023 12173 12026
rect 12207 12023 12219 12057
rect 12161 12017 12219 12023
rect 1104 11964 28888 11986
rect 1104 11912 5982 11964
rect 6034 11912 6046 11964
rect 6098 11912 6110 11964
rect 6162 11912 6174 11964
rect 6226 11912 15982 11964
rect 16034 11912 16046 11964
rect 16098 11912 16110 11964
rect 16162 11912 16174 11964
rect 16226 11912 25982 11964
rect 26034 11912 26046 11964
rect 26098 11912 26110 11964
rect 26162 11912 26174 11964
rect 26226 11912 28888 11964
rect 1104 11890 28888 11912
rect 8021 11853 8079 11859
rect 8021 11819 8033 11853
rect 8067 11850 8079 11853
rect 8478 11850 8484 11862
rect 8067 11822 8484 11850
rect 8067 11819 8079 11822
rect 8021 11813 8079 11819
rect 8478 11810 8484 11822
rect 8536 11810 8542 11862
rect 11974 11850 11980 11862
rect 11935 11822 11980 11850
rect 11974 11810 11980 11822
rect 12032 11810 12038 11862
rect 12161 11853 12219 11859
rect 12161 11819 12173 11853
rect 12207 11850 12219 11853
rect 13538 11850 13544 11862
rect 12207 11822 13544 11850
rect 12207 11819 12219 11822
rect 12161 11813 12219 11819
rect 13538 11810 13544 11822
rect 13596 11850 13602 11862
rect 13909 11853 13967 11859
rect 13909 11850 13921 11853
rect 13596 11822 13921 11850
rect 13596 11810 13602 11822
rect 13909 11819 13921 11822
rect 13955 11819 13967 11853
rect 13909 11813 13967 11819
rect 24394 11810 24400 11862
rect 24452 11850 24458 11862
rect 24489 11853 24547 11859
rect 24489 11850 24501 11853
rect 24452 11822 24501 11850
rect 24452 11810 24458 11822
rect 24489 11819 24501 11822
rect 24535 11819 24547 11853
rect 24489 11813 24547 11819
rect 13078 11742 13084 11794
rect 13136 11782 13142 11794
rect 13173 11785 13231 11791
rect 13173 11782 13185 11785
rect 13136 11754 13185 11782
rect 13136 11742 13142 11754
rect 13173 11751 13185 11754
rect 13219 11751 13231 11785
rect 13173 11745 13231 11751
rect 12066 11674 12072 11726
rect 12124 11714 12130 11726
rect 12713 11717 12771 11723
rect 12713 11714 12725 11717
rect 12124 11686 12725 11714
rect 12124 11674 12130 11686
rect 12713 11683 12725 11686
rect 12759 11683 12771 11717
rect 12713 11677 12771 11683
rect 13446 11674 13452 11726
rect 13504 11714 13510 11726
rect 13541 11717 13599 11723
rect 13541 11714 13553 11717
rect 13504 11686 13553 11714
rect 13504 11674 13510 11686
rect 13541 11683 13553 11686
rect 13587 11683 13599 11717
rect 13541 11677 13599 11683
rect 1397 11649 1455 11655
rect 1397 11615 1409 11649
rect 1443 11646 1455 11649
rect 1578 11646 1584 11658
rect 1443 11618 1584 11646
rect 1443 11615 1455 11618
rect 1397 11609 1455 11615
rect 1578 11606 1584 11618
rect 1636 11646 1642 11658
rect 1949 11649 2007 11655
rect 1949 11646 1961 11649
rect 1636 11618 1961 11646
rect 1636 11606 1642 11618
rect 1949 11615 1961 11618
rect 1995 11615 2007 11649
rect 1949 11609 2007 11615
rect 11974 11606 11980 11658
rect 12032 11646 12038 11658
rect 12618 11646 12624 11658
rect 12032 11618 12624 11646
rect 12032 11606 12038 11618
rect 12618 11606 12624 11618
rect 12676 11606 12682 11658
rect 23937 11649 23995 11655
rect 23937 11615 23949 11649
rect 23983 11646 23995 11649
rect 24394 11646 24400 11658
rect 23983 11618 24400 11646
rect 23983 11615 23995 11618
rect 23937 11609 23995 11615
rect 24394 11606 24400 11618
rect 24452 11606 24458 11658
rect 1581 11513 1639 11519
rect 1581 11479 1593 11513
rect 1627 11510 1639 11513
rect 2130 11510 2136 11522
rect 1627 11482 2136 11510
rect 1627 11479 1639 11482
rect 1581 11473 1639 11479
rect 2130 11470 2136 11482
rect 2188 11470 2194 11522
rect 8294 11510 8300 11522
rect 8255 11482 8300 11510
rect 8294 11470 8300 11482
rect 8352 11470 8358 11522
rect 8662 11510 8668 11522
rect 8623 11482 8668 11510
rect 8662 11470 8668 11482
rect 8720 11470 8726 11522
rect 12158 11470 12164 11522
rect 12216 11510 12222 11522
rect 12529 11513 12587 11519
rect 12529 11510 12541 11513
rect 12216 11482 12541 11510
rect 12216 11470 12222 11482
rect 12529 11479 12541 11482
rect 12575 11479 12587 11513
rect 24118 11510 24124 11522
rect 24079 11482 24124 11510
rect 12529 11473 12587 11479
rect 24118 11470 24124 11482
rect 24176 11470 24182 11522
rect 1104 11420 28888 11442
rect 1104 11368 10982 11420
rect 11034 11368 11046 11420
rect 11098 11368 11110 11420
rect 11162 11368 11174 11420
rect 11226 11368 20982 11420
rect 21034 11368 21046 11420
rect 21098 11368 21110 11420
rect 21162 11368 21174 11420
rect 21226 11368 28888 11420
rect 1104 11346 28888 11368
rect 7745 11309 7803 11315
rect 7745 11275 7757 11309
rect 7791 11306 7803 11309
rect 8662 11306 8668 11318
rect 7791 11278 8668 11306
rect 7791 11275 7803 11278
rect 7745 11269 7803 11275
rect 8662 11266 8668 11278
rect 8720 11266 8726 11318
rect 12158 11306 12164 11318
rect 12119 11278 12164 11306
rect 12158 11266 12164 11278
rect 12216 11266 12222 11318
rect 8110 11238 8116 11250
rect 8071 11210 8116 11238
rect 8110 11198 8116 11210
rect 8168 11198 8174 11250
rect 1397 11173 1455 11179
rect 1397 11139 1409 11173
rect 1443 11170 1455 11173
rect 2038 11170 2044 11182
rect 1443 11142 2044 11170
rect 1443 11139 1455 11142
rect 1397 11133 1455 11139
rect 2038 11130 2044 11142
rect 2096 11130 2102 11182
rect 7190 11130 7196 11182
rect 7248 11170 7254 11182
rect 23934 11170 23940 11182
rect 7248 11142 8340 11170
rect 23895 11142 23940 11170
rect 7248 11130 7254 11142
rect 8312 11114 8340 11142
rect 23934 11130 23940 11142
rect 23992 11130 23998 11182
rect 7374 11062 7380 11114
rect 7432 11102 7438 11114
rect 8205 11105 8263 11111
rect 8205 11102 8217 11105
rect 7432 11074 8217 11102
rect 7432 11062 7438 11074
rect 8205 11071 8217 11074
rect 8251 11071 8263 11105
rect 8205 11065 8263 11071
rect 8294 11062 8300 11114
rect 8352 11102 8358 11114
rect 8352 11074 8445 11102
rect 8352 11062 8358 11074
rect 1581 11037 1639 11043
rect 1581 11003 1593 11037
rect 1627 11034 1639 11037
rect 1946 11034 1952 11046
rect 1627 11006 1952 11034
rect 1627 11003 1639 11006
rect 1581 10997 1639 11003
rect 1946 10994 1952 11006
rect 2004 10994 2010 11046
rect 24121 11037 24179 11043
rect 24121 11003 24133 11037
rect 24167 11034 24179 11037
rect 24854 11034 24860 11046
rect 24167 11006 24860 11034
rect 24167 11003 24179 11006
rect 24121 10997 24179 11003
rect 24854 10994 24860 11006
rect 24912 10994 24918 11046
rect 1104 10876 28888 10898
rect 1104 10824 5982 10876
rect 6034 10824 6046 10876
rect 6098 10824 6110 10876
rect 6162 10824 6174 10876
rect 6226 10824 15982 10876
rect 16034 10824 16046 10876
rect 16098 10824 16110 10876
rect 16162 10824 16174 10876
rect 16226 10824 25982 10876
rect 26034 10824 26046 10876
rect 26098 10824 26110 10876
rect 26162 10824 26174 10876
rect 26226 10824 28888 10876
rect 1104 10802 28888 10824
rect 2038 10762 2044 10774
rect 1999 10734 2044 10762
rect 2038 10722 2044 10734
rect 2096 10722 2102 10774
rect 2406 10762 2412 10774
rect 2367 10734 2412 10762
rect 2406 10722 2412 10734
rect 2464 10722 2470 10774
rect 7098 10762 7104 10774
rect 7059 10734 7104 10762
rect 7098 10722 7104 10734
rect 7156 10722 7162 10774
rect 7929 10765 7987 10771
rect 7929 10731 7941 10765
rect 7975 10762 7987 10765
rect 8202 10762 8208 10774
rect 7975 10734 8208 10762
rect 7975 10731 7987 10734
rect 7929 10725 7987 10731
rect 8202 10722 8208 10734
rect 8260 10722 8266 10774
rect 8294 10722 8300 10774
rect 8352 10762 8358 10774
rect 8941 10765 8999 10771
rect 8941 10762 8953 10765
rect 8352 10734 8953 10762
rect 8352 10722 8358 10734
rect 8588 10638 8616 10734
rect 8941 10731 8953 10734
rect 8987 10731 8999 10765
rect 23934 10762 23940 10774
rect 23895 10734 23940 10762
rect 8941 10725 8999 10731
rect 23934 10722 23940 10734
rect 23992 10722 23998 10774
rect 8570 10626 8576 10638
rect 8483 10598 8576 10626
rect 8570 10586 8576 10598
rect 8628 10586 8634 10638
rect 1397 10561 1455 10567
rect 1397 10527 1409 10561
rect 1443 10558 1455 10561
rect 2406 10558 2412 10570
rect 1443 10530 2412 10558
rect 1443 10527 1455 10530
rect 1397 10521 1455 10527
rect 2406 10518 2412 10530
rect 2464 10518 2470 10570
rect 8294 10490 8300 10502
rect 8255 10462 8300 10490
rect 8294 10450 8300 10462
rect 8352 10450 8358 10502
rect 1581 10425 1639 10431
rect 1581 10391 1593 10425
rect 1627 10422 1639 10425
rect 1762 10422 1768 10434
rect 1627 10394 1768 10422
rect 1627 10391 1639 10394
rect 1581 10385 1639 10391
rect 1762 10382 1768 10394
rect 1820 10382 1826 10434
rect 7374 10422 7380 10434
rect 7335 10394 7380 10422
rect 7374 10382 7380 10394
rect 7432 10382 7438 10434
rect 7834 10422 7840 10434
rect 7747 10394 7840 10422
rect 7834 10382 7840 10394
rect 7892 10422 7898 10434
rect 8386 10422 8392 10434
rect 7892 10394 8392 10422
rect 7892 10382 7898 10394
rect 8386 10382 8392 10394
rect 8444 10382 8450 10434
rect 1104 10332 28888 10354
rect 1104 10280 10982 10332
rect 11034 10280 11046 10332
rect 11098 10280 11110 10332
rect 11162 10280 11174 10332
rect 11226 10280 20982 10332
rect 21034 10280 21046 10332
rect 21098 10280 21110 10332
rect 21162 10280 21174 10332
rect 21226 10280 28888 10332
rect 1104 10258 28888 10280
rect 8021 10221 8079 10227
rect 8021 10187 8033 10221
rect 8067 10218 8079 10221
rect 8294 10218 8300 10230
rect 8067 10190 8300 10218
rect 8067 10187 8079 10190
rect 8021 10181 8079 10187
rect 8294 10178 8300 10190
rect 8352 10178 8358 10230
rect 8389 10221 8447 10227
rect 8389 10187 8401 10221
rect 8435 10218 8447 10221
rect 8570 10218 8576 10230
rect 8435 10190 8576 10218
rect 8435 10187 8447 10190
rect 8389 10181 8447 10187
rect 8570 10178 8576 10190
rect 8628 10178 8634 10230
rect 1397 10085 1455 10091
rect 1397 10051 1409 10085
rect 1443 10082 1455 10085
rect 2222 10082 2228 10094
rect 1443 10054 2228 10082
rect 1443 10051 1455 10054
rect 1397 10045 1455 10051
rect 2222 10042 2228 10054
rect 2280 10042 2286 10094
rect 1578 9878 1584 9890
rect 1539 9850 1584 9878
rect 1578 9838 1584 9850
rect 1636 9838 1642 9890
rect 1104 9788 28888 9810
rect 1104 9736 5982 9788
rect 6034 9736 6046 9788
rect 6098 9736 6110 9788
rect 6162 9736 6174 9788
rect 6226 9736 15982 9788
rect 16034 9736 16046 9788
rect 16098 9736 16110 9788
rect 16162 9736 16174 9788
rect 16226 9736 25982 9788
rect 26034 9736 26046 9788
rect 26098 9736 26110 9788
rect 26162 9736 26174 9788
rect 26226 9736 28888 9788
rect 1104 9714 28888 9736
rect 2041 9677 2099 9683
rect 2041 9643 2053 9677
rect 2087 9674 2099 9677
rect 2222 9674 2228 9686
rect 2087 9646 2228 9674
rect 2087 9643 2099 9646
rect 2041 9637 2099 9643
rect 2222 9634 2228 9646
rect 2280 9634 2286 9686
rect 2409 9609 2467 9615
rect 2409 9575 2421 9609
rect 2455 9606 2467 9609
rect 2498 9606 2504 9618
rect 2455 9578 2504 9606
rect 2455 9575 2467 9578
rect 2409 9569 2467 9575
rect 1397 9473 1455 9479
rect 1397 9439 1409 9473
rect 1443 9470 1455 9473
rect 2424 9470 2452 9569
rect 2498 9566 2504 9578
rect 2556 9566 2562 9618
rect 23934 9470 23940 9482
rect 1443 9442 2452 9470
rect 23895 9442 23940 9470
rect 1443 9439 1455 9442
rect 1397 9433 1455 9439
rect 23934 9430 23940 9442
rect 23992 9470 23998 9482
rect 24489 9473 24547 9479
rect 24489 9470 24501 9473
rect 23992 9442 24501 9470
rect 23992 9430 23998 9442
rect 24489 9439 24501 9442
rect 24535 9439 24547 9473
rect 24489 9433 24547 9439
rect 1578 9334 1584 9346
rect 1539 9306 1584 9334
rect 1578 9294 1584 9306
rect 1636 9294 1642 9346
rect 24118 9334 24124 9346
rect 24079 9306 24124 9334
rect 24118 9294 24124 9306
rect 24176 9294 24182 9346
rect 1104 9244 28888 9266
rect 1104 9192 10982 9244
rect 11034 9192 11046 9244
rect 11098 9192 11110 9244
rect 11162 9192 11174 9244
rect 11226 9192 20982 9244
rect 21034 9192 21046 9244
rect 21098 9192 21110 9244
rect 21162 9192 21174 9244
rect 21226 9192 28888 9244
rect 1104 9170 28888 9192
rect 1394 8994 1400 9006
rect 1355 8966 1400 8994
rect 1394 8954 1400 8966
rect 1452 8954 1458 9006
rect 23934 8994 23940 9006
rect 23895 8966 23940 8994
rect 23934 8954 23940 8966
rect 23992 8954 23998 9006
rect 1394 8750 1400 8802
rect 1452 8790 1458 8802
rect 1581 8793 1639 8799
rect 1581 8790 1593 8793
rect 1452 8762 1593 8790
rect 1452 8750 1458 8762
rect 1581 8759 1593 8762
rect 1627 8759 1639 8793
rect 1581 8753 1639 8759
rect 1946 8750 1952 8802
rect 2004 8790 2010 8802
rect 2682 8790 2688 8802
rect 2004 8762 2688 8790
rect 2004 8750 2010 8762
rect 2682 8750 2688 8762
rect 2740 8750 2746 8802
rect 24118 8790 24124 8802
rect 24079 8762 24124 8790
rect 24118 8750 24124 8762
rect 24176 8750 24182 8802
rect 1104 8700 28888 8722
rect 1104 8648 5982 8700
rect 6034 8648 6046 8700
rect 6098 8648 6110 8700
rect 6162 8648 6174 8700
rect 6226 8648 15982 8700
rect 16034 8648 16046 8700
rect 16098 8648 16110 8700
rect 16162 8648 16174 8700
rect 16226 8648 25982 8700
rect 26034 8648 26046 8700
rect 26098 8648 26110 8700
rect 26162 8648 26174 8700
rect 26226 8648 28888 8700
rect 1104 8626 28888 8648
rect 1486 8546 1492 8598
rect 1544 8586 1550 8598
rect 1581 8589 1639 8595
rect 1581 8586 1593 8589
rect 1544 8558 1593 8586
rect 1544 8546 1550 8558
rect 1581 8555 1593 8558
rect 1627 8555 1639 8589
rect 23750 8586 23756 8598
rect 23711 8558 23756 8586
rect 1581 8549 1639 8555
rect 23750 8546 23756 8558
rect 23808 8546 23814 8598
rect 23934 8546 23940 8598
rect 23992 8586 23998 8598
rect 24489 8589 24547 8595
rect 24489 8586 24501 8589
rect 23992 8558 24501 8586
rect 23992 8546 23998 8558
rect 24489 8555 24501 8558
rect 24535 8555 24547 8589
rect 24489 8549 24547 8555
rect 23474 8478 23480 8530
rect 23532 8518 23538 8530
rect 24121 8521 24179 8527
rect 24121 8518 24133 8521
rect 23532 8490 24133 8518
rect 23532 8478 23538 8490
rect 24121 8487 24133 8490
rect 24167 8487 24179 8521
rect 24121 8481 24179 8487
rect 23750 8342 23756 8394
rect 23808 8382 23814 8394
rect 23937 8385 23995 8391
rect 23937 8382 23949 8385
rect 23808 8354 23949 8382
rect 23808 8342 23814 8354
rect 23937 8351 23949 8354
rect 23983 8351 23995 8385
rect 23937 8345 23995 8351
rect 1104 8156 28888 8178
rect 1104 8104 10982 8156
rect 11034 8104 11046 8156
rect 11098 8104 11110 8156
rect 11162 8104 11174 8156
rect 11226 8104 20982 8156
rect 21034 8104 21046 8156
rect 21098 8104 21110 8156
rect 21162 8104 21174 8156
rect 21226 8104 28888 8156
rect 1104 8082 28888 8104
rect 24118 8042 24124 8054
rect 24079 8014 24124 8042
rect 24118 8002 24124 8014
rect 24176 8002 24182 8054
rect 23934 7906 23940 7918
rect 23895 7878 23940 7906
rect 23934 7866 23940 7878
rect 23992 7866 23998 7918
rect 1104 7612 28888 7634
rect 1104 7560 5982 7612
rect 6034 7560 6046 7612
rect 6098 7560 6110 7612
rect 6162 7560 6174 7612
rect 6226 7560 15982 7612
rect 16034 7560 16046 7612
rect 16098 7560 16110 7612
rect 16162 7560 16174 7612
rect 16226 7560 25982 7612
rect 26034 7560 26046 7612
rect 26098 7560 26110 7612
rect 26162 7560 26174 7612
rect 26226 7560 28888 7612
rect 1104 7538 28888 7560
rect 22462 7498 22468 7510
rect 22423 7470 22468 7498
rect 22462 7458 22468 7470
rect 22520 7458 22526 7510
rect 22922 7498 22928 7510
rect 22883 7470 22928 7498
rect 22922 7458 22928 7470
rect 22980 7458 22986 7510
rect 23934 7498 23940 7510
rect 23895 7470 23940 7498
rect 23934 7458 23940 7470
rect 23992 7458 23998 7510
rect 18598 7430 18604 7442
rect 18559 7402 18604 7430
rect 18598 7390 18604 7402
rect 18656 7390 18662 7442
rect 13078 7294 13084 7306
rect 13039 7266 13084 7294
rect 13078 7254 13084 7266
rect 13136 7294 13142 7306
rect 13633 7297 13691 7303
rect 13633 7294 13645 7297
rect 13136 7266 13645 7294
rect 13136 7254 13142 7266
rect 13633 7263 13645 7266
rect 13679 7263 13691 7297
rect 18414 7294 18420 7306
rect 18375 7266 18420 7294
rect 13633 7257 13691 7263
rect 18414 7254 18420 7266
rect 18472 7294 18478 7306
rect 18969 7297 19027 7303
rect 18969 7294 18981 7297
rect 18472 7266 18981 7294
rect 18472 7254 18478 7266
rect 18969 7263 18981 7266
rect 19015 7263 19027 7297
rect 18969 7257 19027 7263
rect 22281 7297 22339 7303
rect 22281 7263 22293 7297
rect 22327 7294 22339 7297
rect 22922 7294 22928 7306
rect 22327 7266 22928 7294
rect 22327 7263 22339 7266
rect 22281 7257 22339 7263
rect 22922 7254 22928 7266
rect 22980 7254 22986 7306
rect 13262 7158 13268 7170
rect 13223 7130 13268 7158
rect 13262 7118 13268 7130
rect 13320 7118 13326 7170
rect 1104 7068 28888 7090
rect 1104 7016 10982 7068
rect 11034 7016 11046 7068
rect 11098 7016 11110 7068
rect 11162 7016 11174 7068
rect 11226 7016 20982 7068
rect 21034 7016 21046 7068
rect 21098 7016 21110 7068
rect 21162 7016 21174 7068
rect 21226 7016 28888 7068
rect 1104 6994 28888 7016
rect 1302 6846 1308 6898
rect 1360 6886 1366 6898
rect 1854 6886 1860 6898
rect 1360 6858 1860 6886
rect 1360 6846 1366 6858
rect 1854 6846 1860 6858
rect 1912 6846 1918 6898
rect 14734 6818 14740 6830
rect 14695 6790 14740 6818
rect 14734 6778 14740 6790
rect 14792 6778 14798 6830
rect 23937 6821 23995 6827
rect 23937 6787 23949 6821
rect 23983 6818 23995 6821
rect 24026 6818 24032 6830
rect 23983 6790 24032 6818
rect 23983 6787 23995 6790
rect 23937 6781 23995 6787
rect 24026 6778 24032 6790
rect 24084 6778 24090 6830
rect 14918 6682 14924 6694
rect 14879 6654 14924 6682
rect 14918 6642 14924 6654
rect 14976 6642 14982 6694
rect 24118 6682 24124 6694
rect 24079 6654 24124 6682
rect 24118 6642 24124 6654
rect 24176 6642 24182 6694
rect 1104 6524 28888 6546
rect 1104 6472 5982 6524
rect 6034 6472 6046 6524
rect 6098 6472 6110 6524
rect 6162 6472 6174 6524
rect 6226 6472 15982 6524
rect 16034 6472 16046 6524
rect 16098 6472 16110 6524
rect 16162 6472 16174 6524
rect 16226 6472 25982 6524
rect 26034 6472 26046 6524
rect 26098 6472 26110 6524
rect 26162 6472 26174 6524
rect 26226 6472 28888 6524
rect 1104 6450 28888 6472
rect 14734 6410 14740 6422
rect 14695 6382 14740 6410
rect 14734 6370 14740 6382
rect 14792 6370 14798 6422
rect 24026 6410 24032 6422
rect 23987 6382 24032 6410
rect 24026 6370 24032 6382
rect 24084 6370 24090 6422
rect 1104 5980 28888 6002
rect 1104 5928 10982 5980
rect 11034 5928 11046 5980
rect 11098 5928 11110 5980
rect 11162 5928 11174 5980
rect 11226 5928 20982 5980
rect 21034 5928 21046 5980
rect 21098 5928 21110 5980
rect 21162 5928 21174 5980
rect 21226 5928 28888 5980
rect 1104 5906 28888 5928
rect 13078 5866 13084 5878
rect 13039 5838 13084 5866
rect 13078 5826 13084 5838
rect 13136 5826 13142 5878
rect 4154 5730 4160 5742
rect 4115 5702 4160 5730
rect 4154 5690 4160 5702
rect 4212 5690 4218 5742
rect 12897 5733 12955 5739
rect 12897 5699 12909 5733
rect 12943 5730 12955 5733
rect 13630 5730 13636 5742
rect 12943 5702 13636 5730
rect 12943 5699 12955 5702
rect 12897 5693 12955 5699
rect 13630 5690 13636 5702
rect 13688 5690 13694 5742
rect 4338 5594 4344 5606
rect 4299 5566 4344 5594
rect 4338 5554 4344 5566
rect 4396 5554 4402 5606
rect 1104 5436 28888 5458
rect 1104 5384 5982 5436
rect 6034 5384 6046 5436
rect 6098 5384 6110 5436
rect 6162 5384 6174 5436
rect 6226 5384 15982 5436
rect 16034 5384 16046 5436
rect 16098 5384 16110 5436
rect 16162 5384 16174 5436
rect 16226 5384 25982 5436
rect 26034 5384 26046 5436
rect 26098 5384 26110 5436
rect 26162 5384 26174 5436
rect 26226 5384 28888 5436
rect 1104 5362 28888 5384
rect 4154 5282 4160 5334
rect 4212 5322 4218 5334
rect 4249 5325 4307 5331
rect 4249 5322 4261 5325
rect 4212 5294 4261 5322
rect 4212 5282 4218 5294
rect 4249 5291 4261 5294
rect 4295 5291 4307 5325
rect 13630 5322 13636 5334
rect 13591 5294 13636 5322
rect 4249 5285 4307 5291
rect 13630 5282 13636 5294
rect 13688 5282 13694 5334
rect 24581 5325 24639 5331
rect 24581 5291 24593 5325
rect 24627 5322 24639 5325
rect 24762 5322 24768 5334
rect 24627 5294 24768 5322
rect 24627 5291 24639 5294
rect 24581 5285 24639 5291
rect 12618 5118 12624 5130
rect 12579 5090 12624 5118
rect 12618 5078 12624 5090
rect 12676 5118 12682 5130
rect 13173 5121 13231 5127
rect 13173 5118 13185 5121
rect 12676 5090 13185 5118
rect 12676 5078 12682 5090
rect 13173 5087 13185 5090
rect 13219 5087 13231 5121
rect 13173 5081 13231 5087
rect 23937 5121 23995 5127
rect 23937 5087 23949 5121
rect 23983 5118 23995 5121
rect 24596 5118 24624 5285
rect 24762 5282 24768 5294
rect 24820 5282 24826 5334
rect 23983 5090 24624 5118
rect 23983 5087 23995 5090
rect 23937 5081 23995 5087
rect 12802 4982 12808 4994
rect 12763 4954 12808 4982
rect 12802 4942 12808 4954
rect 12860 4942 12866 4994
rect 24118 4982 24124 4994
rect 24079 4954 24124 4982
rect 24118 4942 24124 4954
rect 24176 4942 24182 4994
rect 1104 4892 28888 4914
rect 1104 4840 10982 4892
rect 11034 4840 11046 4892
rect 11098 4840 11110 4892
rect 11162 4840 11174 4892
rect 11226 4840 20982 4892
rect 21034 4840 21046 4892
rect 21098 4840 21110 4892
rect 21162 4840 21174 4892
rect 21226 4840 28888 4892
rect 1104 4818 28888 4840
rect 15562 4642 15568 4654
rect 15523 4614 15568 4642
rect 15562 4602 15568 4614
rect 15620 4602 15626 4654
rect 20438 4642 20444 4654
rect 20399 4614 20444 4642
rect 20438 4602 20444 4614
rect 20496 4602 20502 4654
rect 15746 4506 15752 4518
rect 15707 4478 15752 4506
rect 15746 4466 15752 4478
rect 15804 4466 15810 4518
rect 20622 4506 20628 4518
rect 20583 4478 20628 4506
rect 20622 4466 20628 4478
rect 20680 4466 20686 4518
rect 1104 4348 28888 4370
rect 1104 4296 5982 4348
rect 6034 4296 6046 4348
rect 6098 4296 6110 4348
rect 6162 4296 6174 4348
rect 6226 4296 15982 4348
rect 16034 4296 16046 4348
rect 16098 4296 16110 4348
rect 16162 4296 16174 4348
rect 16226 4296 25982 4348
rect 26034 4296 26046 4348
rect 26098 4296 26110 4348
rect 26162 4296 26174 4348
rect 26226 4296 28888 4348
rect 1104 4274 28888 4296
rect 15562 4234 15568 4246
rect 15523 4206 15568 4234
rect 15562 4194 15568 4206
rect 15620 4194 15626 4246
rect 20438 4234 20444 4246
rect 20399 4206 20444 4234
rect 20438 4194 20444 4206
rect 20496 4194 20502 4246
rect 21450 4098 21456 4110
rect 20916 4070 21456 4098
rect 20916 4039 20944 4070
rect 21450 4058 21456 4070
rect 21508 4058 21514 4110
rect 20901 4033 20959 4039
rect 20901 3999 20913 4033
rect 20947 3999 20959 4033
rect 23934 4030 23940 4042
rect 23895 4002 23940 4030
rect 20901 3993 20959 3999
rect 23934 3990 23940 4002
rect 23992 4030 23998 4042
rect 24489 4033 24547 4039
rect 24489 4030 24501 4033
rect 23992 4002 24501 4030
rect 23992 3990 23998 4002
rect 24489 3999 24501 4002
rect 24535 3999 24547 4033
rect 24489 3993 24547 3999
rect 20714 3854 20720 3906
rect 20772 3894 20778 3906
rect 21085 3897 21143 3903
rect 21085 3894 21097 3897
rect 20772 3866 21097 3894
rect 20772 3854 20778 3866
rect 21085 3863 21097 3866
rect 21131 3863 21143 3897
rect 24118 3894 24124 3906
rect 24079 3866 24124 3894
rect 21085 3857 21143 3863
rect 24118 3854 24124 3866
rect 24176 3854 24182 3906
rect 1104 3804 28888 3826
rect 1104 3752 10982 3804
rect 11034 3752 11046 3804
rect 11098 3752 11110 3804
rect 11162 3752 11174 3804
rect 11226 3752 20982 3804
rect 21034 3752 21046 3804
rect 21098 3752 21110 3804
rect 21162 3752 21174 3804
rect 21226 3752 28888 3804
rect 1104 3730 28888 3752
rect 23842 3514 23848 3566
rect 23900 3554 23906 3566
rect 23937 3557 23995 3563
rect 23937 3554 23949 3557
rect 23900 3526 23949 3554
rect 23900 3514 23906 3526
rect 23937 3523 23949 3526
rect 23983 3554 23995 3557
rect 24670 3554 24676 3566
rect 23983 3526 24676 3554
rect 23983 3523 23995 3526
rect 23937 3517 23995 3523
rect 24670 3514 24676 3526
rect 24728 3514 24734 3566
rect 24118 3418 24124 3430
rect 24079 3390 24124 3418
rect 24118 3378 24124 3390
rect 24176 3378 24182 3430
rect 1104 3260 28888 3282
rect 1104 3208 5982 3260
rect 6034 3208 6046 3260
rect 6098 3208 6110 3260
rect 6162 3208 6174 3260
rect 6226 3208 15982 3260
rect 16034 3208 16046 3260
rect 16098 3208 16110 3260
rect 16162 3208 16174 3260
rect 16226 3208 25982 3260
rect 26034 3208 26046 3260
rect 26098 3208 26110 3260
rect 26162 3208 26174 3260
rect 26226 3208 28888 3260
rect 1104 3186 28888 3208
rect 1946 3146 1952 3158
rect 1907 3118 1952 3146
rect 1946 3106 1952 3118
rect 2004 3106 2010 3158
rect 23842 3146 23848 3158
rect 23803 3118 23848 3146
rect 23842 3106 23848 3118
rect 23900 3106 23906 3158
rect 1397 2945 1455 2951
rect 1397 2911 1409 2945
rect 1443 2942 1455 2945
rect 1946 2942 1952 2954
rect 1443 2914 1952 2942
rect 1443 2911 1455 2914
rect 1397 2905 1455 2911
rect 1946 2902 1952 2914
rect 2004 2902 2010 2954
rect 23934 2942 23940 2954
rect 23895 2914 23940 2942
rect 23934 2902 23940 2914
rect 23992 2942 23998 2954
rect 24489 2945 24547 2951
rect 24489 2942 24501 2945
rect 23992 2914 24501 2942
rect 23992 2902 23998 2914
rect 24489 2911 24501 2914
rect 24535 2911 24547 2945
rect 24489 2905 24547 2911
rect 1581 2809 1639 2815
rect 1581 2775 1593 2809
rect 1627 2806 1639 2809
rect 9490 2806 9496 2818
rect 1627 2778 9496 2806
rect 1627 2775 1639 2778
rect 1581 2769 1639 2775
rect 9490 2766 9496 2778
rect 9548 2766 9554 2818
rect 24121 2809 24179 2815
rect 24121 2775 24133 2809
rect 24167 2806 24179 2809
rect 24854 2806 24860 2818
rect 24167 2778 24860 2806
rect 24167 2775 24179 2778
rect 24121 2769 24179 2775
rect 24854 2766 24860 2778
rect 24912 2766 24918 2818
rect 1104 2716 28888 2738
rect 1104 2664 10982 2716
rect 11034 2664 11046 2716
rect 11098 2664 11110 2716
rect 11162 2664 11174 2716
rect 11226 2664 20982 2716
rect 21034 2664 21046 2716
rect 21098 2664 21110 2716
rect 21162 2664 21174 2716
rect 21226 2664 28888 2716
rect 1104 2642 28888 2664
rect 24210 2602 24216 2614
rect 24171 2574 24216 2602
rect 24210 2562 24216 2574
rect 24268 2562 24274 2614
rect 1397 2469 1455 2475
rect 1397 2435 1409 2469
rect 1443 2435 1455 2469
rect 24026 2466 24032 2478
rect 23987 2438 24032 2466
rect 1397 2429 1455 2435
rect 1412 2398 1440 2429
rect 24026 2426 24032 2438
rect 24084 2466 24090 2478
rect 24581 2469 24639 2475
rect 24581 2466 24593 2469
rect 24084 2438 24593 2466
rect 24084 2426 24090 2438
rect 24581 2435 24593 2438
rect 24627 2435 24639 2469
rect 25130 2466 25136 2478
rect 25091 2438 25136 2466
rect 24581 2429 24639 2435
rect 25130 2426 25136 2438
rect 25188 2466 25194 2478
rect 25685 2469 25743 2475
rect 25685 2466 25697 2469
rect 25188 2438 25697 2466
rect 25188 2426 25194 2438
rect 25685 2435 25697 2438
rect 25731 2435 25743 2469
rect 25685 2429 25743 2435
rect 2038 2398 2044 2410
rect 1412 2370 2044 2398
rect 2038 2358 2044 2370
rect 2096 2358 2102 2410
rect 1578 2262 1584 2274
rect 1539 2234 1584 2262
rect 1578 2222 1584 2234
rect 1636 2222 1642 2274
rect 25314 2262 25320 2274
rect 25275 2234 25320 2262
rect 25314 2222 25320 2234
rect 25372 2222 25378 2274
rect 1104 2172 28888 2194
rect 1104 2120 5982 2172
rect 6034 2120 6046 2172
rect 6098 2120 6110 2172
rect 6162 2120 6174 2172
rect 6226 2120 15982 2172
rect 16034 2120 16046 2172
rect 16098 2120 16110 2172
rect 16162 2120 16174 2172
rect 16226 2120 25982 2172
rect 26034 2120 26046 2172
rect 26098 2120 26110 2172
rect 26162 2120 26174 2172
rect 26226 2120 28888 2172
rect 1104 2098 28888 2120
<< via1 >>
rect 5982 21704 6034 21756
rect 6046 21704 6098 21756
rect 6110 21704 6162 21756
rect 6174 21704 6226 21756
rect 15982 21704 16034 21756
rect 16046 21704 16098 21756
rect 16110 21704 16162 21756
rect 16174 21704 16226 21756
rect 25982 21704 26034 21756
rect 26046 21704 26098 21756
rect 26110 21704 26162 21756
rect 26174 21704 26226 21756
rect 10982 21160 11034 21212
rect 11046 21160 11098 21212
rect 11110 21160 11162 21212
rect 11174 21160 11226 21212
rect 20982 21160 21034 21212
rect 21046 21160 21098 21212
rect 21110 21160 21162 21212
rect 21174 21160 21226 21212
rect 3424 20718 3476 20770
rect 19432 20718 19484 20770
rect 19616 20718 19668 20770
rect 24860 20718 24912 20770
rect 5982 20616 6034 20668
rect 6046 20616 6098 20668
rect 6110 20616 6162 20668
rect 6174 20616 6226 20668
rect 15982 20616 16034 20668
rect 16046 20616 16098 20668
rect 16110 20616 16162 20668
rect 16174 20616 16226 20668
rect 25982 20616 26034 20668
rect 26046 20616 26098 20668
rect 26110 20616 26162 20668
rect 26174 20616 26226 20668
rect 10982 20072 11034 20124
rect 11046 20072 11098 20124
rect 11110 20072 11162 20124
rect 11174 20072 11226 20124
rect 20982 20072 21034 20124
rect 21046 20072 21098 20124
rect 21110 20072 21162 20124
rect 21174 20072 21226 20124
rect 5982 19528 6034 19580
rect 6046 19528 6098 19580
rect 6110 19528 6162 19580
rect 6174 19528 6226 19580
rect 15982 19528 16034 19580
rect 16046 19528 16098 19580
rect 16110 19528 16162 19580
rect 16174 19528 16226 19580
rect 25982 19528 26034 19580
rect 26046 19528 26098 19580
rect 26110 19528 26162 19580
rect 26174 19528 26226 19580
rect 24768 19222 24820 19274
rect 23480 19086 23532 19138
rect 10982 18984 11034 19036
rect 11046 18984 11098 19036
rect 11110 18984 11162 19036
rect 11174 18984 11226 19036
rect 20982 18984 21034 19036
rect 21046 18984 21098 19036
rect 21110 18984 21162 19036
rect 21174 18984 21226 19036
rect 16764 18925 16816 18934
rect 16764 18891 16773 18925
rect 16773 18891 16807 18925
rect 16807 18891 16816 18925
rect 16764 18882 16816 18891
rect 20812 18925 20864 18934
rect 20812 18891 20821 18925
rect 20821 18891 20855 18925
rect 20855 18891 20864 18925
rect 20812 18882 20864 18891
rect 3148 18814 3200 18866
rect 3700 18814 3752 18866
rect 8852 18857 8904 18866
rect 8852 18823 8886 18857
rect 8886 18823 8904 18857
rect 8852 18814 8904 18823
rect 8576 18789 8628 18798
rect 8576 18755 8585 18789
rect 8585 18755 8619 18789
rect 8619 18755 8628 18789
rect 8576 18746 8628 18755
rect 15660 18789 15712 18798
rect 15660 18755 15694 18789
rect 15694 18755 15712 18789
rect 15660 18746 15712 18755
rect 20628 18789 20680 18798
rect 20628 18755 20637 18789
rect 20637 18755 20671 18789
rect 20671 18755 20680 18789
rect 20628 18746 20680 18755
rect 23940 18789 23992 18798
rect 23940 18755 23949 18789
rect 23949 18755 23983 18789
rect 23983 18755 23992 18789
rect 23940 18746 23992 18755
rect 25044 18789 25096 18798
rect 25044 18755 25053 18789
rect 25053 18755 25087 18789
rect 25087 18755 25096 18789
rect 25044 18746 25096 18755
rect 15384 18721 15436 18730
rect 15384 18687 15393 18721
rect 15393 18687 15427 18721
rect 15427 18687 15436 18721
rect 15384 18678 15436 18687
rect 9956 18585 10008 18594
rect 9956 18551 9965 18585
rect 9965 18551 9999 18585
rect 9999 18551 10008 18585
rect 9956 18542 10008 18551
rect 24124 18585 24176 18594
rect 24124 18551 24133 18585
rect 24133 18551 24167 18585
rect 24167 18551 24176 18585
rect 24124 18542 24176 18551
rect 25228 18585 25280 18594
rect 25228 18551 25237 18585
rect 25237 18551 25271 18585
rect 25271 18551 25280 18585
rect 25228 18542 25280 18551
rect 5982 18440 6034 18492
rect 6046 18440 6098 18492
rect 6110 18440 6162 18492
rect 6174 18440 6226 18492
rect 15982 18440 16034 18492
rect 16046 18440 16098 18492
rect 16110 18440 16162 18492
rect 16174 18440 16226 18492
rect 25982 18440 26034 18492
rect 26046 18440 26098 18492
rect 26110 18440 26162 18492
rect 26174 18440 26226 18492
rect 8852 18338 8904 18390
rect 23940 18338 23992 18390
rect 25044 18381 25096 18390
rect 25044 18347 25053 18381
rect 25053 18347 25087 18381
rect 25087 18347 25096 18381
rect 25044 18338 25096 18347
rect 8576 18270 8628 18322
rect 15384 18134 15436 18186
rect 23940 18177 23992 18186
rect 23940 18143 23949 18177
rect 23949 18143 23983 18177
rect 23983 18143 23992 18177
rect 23940 18134 23992 18143
rect 15200 18066 15252 18118
rect 15660 18066 15712 18118
rect 19340 17998 19392 18050
rect 20628 18041 20680 18050
rect 20628 18007 20637 18041
rect 20637 18007 20671 18041
rect 20671 18007 20680 18041
rect 20628 17998 20680 18007
rect 24308 17998 24360 18050
rect 10982 17896 11034 17948
rect 11046 17896 11098 17948
rect 11110 17896 11162 17948
rect 11174 17896 11226 17948
rect 20982 17896 21034 17948
rect 21046 17896 21098 17948
rect 21110 17896 21162 17948
rect 21174 17896 21226 17948
rect 23940 17701 23992 17710
rect 23940 17667 23949 17701
rect 23949 17667 23983 17701
rect 23983 17667 23992 17701
rect 23940 17658 23992 17667
rect 24216 17454 24268 17506
rect 5982 17352 6034 17404
rect 6046 17352 6098 17404
rect 6110 17352 6162 17404
rect 6174 17352 6226 17404
rect 15982 17352 16034 17404
rect 16046 17352 16098 17404
rect 16110 17352 16162 17404
rect 16174 17352 16226 17404
rect 25982 17352 26034 17404
rect 26046 17352 26098 17404
rect 26110 17352 26162 17404
rect 26174 17352 26226 17404
rect 19248 17250 19300 17302
rect 23940 17293 23992 17302
rect 23940 17259 23949 17293
rect 23949 17259 23983 17293
rect 23983 17259 23992 17293
rect 23940 17250 23992 17259
rect 18696 17157 18748 17166
rect 18696 17123 18705 17157
rect 18705 17123 18739 17157
rect 18739 17123 18748 17157
rect 18696 17114 18748 17123
rect 17500 16953 17552 16962
rect 17500 16919 17509 16953
rect 17509 16919 17543 16953
rect 17543 16919 17552 16953
rect 17500 16910 17552 16919
rect 18328 16910 18380 16962
rect 10982 16808 11034 16860
rect 11046 16808 11098 16860
rect 11110 16808 11162 16860
rect 11174 16808 11226 16860
rect 20982 16808 21034 16860
rect 21046 16808 21098 16860
rect 21110 16808 21162 16860
rect 21174 16808 21226 16860
rect 14096 16706 14148 16758
rect 15200 16706 15252 16758
rect 18328 16749 18380 16758
rect 18328 16715 18337 16749
rect 18337 16715 18371 16749
rect 18371 16715 18380 16749
rect 18328 16706 18380 16715
rect 13084 16613 13136 16622
rect 13084 16579 13093 16613
rect 13093 16579 13127 16613
rect 13127 16579 13136 16613
rect 13084 16570 13136 16579
rect 13636 16570 13688 16622
rect 5982 16264 6034 16316
rect 6046 16264 6098 16316
rect 6110 16264 6162 16316
rect 6174 16264 6226 16316
rect 15982 16264 16034 16316
rect 16046 16264 16098 16316
rect 16110 16264 16162 16316
rect 16174 16264 16226 16316
rect 25982 16264 26034 16316
rect 26046 16264 26098 16316
rect 26110 16264 26162 16316
rect 26174 16264 26226 16316
rect 7012 16205 7064 16214
rect 7012 16171 7021 16205
rect 7021 16171 7055 16205
rect 7055 16171 7064 16205
rect 7012 16162 7064 16171
rect 13084 16205 13136 16214
rect 13084 16171 13093 16205
rect 13093 16171 13127 16205
rect 13127 16171 13136 16205
rect 13084 16162 13136 16171
rect 24492 16205 24544 16214
rect 24492 16171 24501 16205
rect 24501 16171 24535 16205
rect 24535 16171 24544 16205
rect 24492 16162 24544 16171
rect 24492 15958 24544 16010
rect 7196 15890 7248 15942
rect 8484 15865 8536 15874
rect 8484 15831 8493 15865
rect 8493 15831 8527 15865
rect 8527 15831 8536 15865
rect 8484 15822 8536 15831
rect 13452 15865 13504 15874
rect 13452 15831 13461 15865
rect 13461 15831 13495 15865
rect 13495 15831 13504 15865
rect 13452 15822 13504 15831
rect 13636 15822 13688 15874
rect 23664 15822 23716 15874
rect 10982 15720 11034 15772
rect 11046 15720 11098 15772
rect 11110 15720 11162 15772
rect 11174 15720 11226 15772
rect 20982 15720 21034 15772
rect 21046 15720 21098 15772
rect 21110 15720 21162 15772
rect 21174 15720 21226 15772
rect 7196 15661 7248 15670
rect 7196 15627 7205 15661
rect 7205 15627 7239 15661
rect 7239 15627 7248 15661
rect 7196 15618 7248 15627
rect 19248 15278 19300 15330
rect 5982 15176 6034 15228
rect 6046 15176 6098 15228
rect 6110 15176 6162 15228
rect 6174 15176 6226 15228
rect 15982 15176 16034 15228
rect 16046 15176 16098 15228
rect 16110 15176 16162 15228
rect 16174 15176 16226 15228
rect 25982 15176 26034 15228
rect 26046 15176 26098 15228
rect 26110 15176 26162 15228
rect 26174 15176 26226 15228
rect 18328 15074 18380 15126
rect 18788 14981 18840 14990
rect 18788 14947 18797 14981
rect 18797 14947 18831 14981
rect 18831 14947 18840 14981
rect 18788 14938 18840 14947
rect 19340 14913 19392 14922
rect 19340 14879 19349 14913
rect 19349 14879 19383 14913
rect 19383 14879 19392 14913
rect 19340 14870 19392 14879
rect 19432 14777 19484 14786
rect 19432 14743 19441 14777
rect 19441 14743 19475 14777
rect 19475 14743 19484 14777
rect 19432 14734 19484 14743
rect 10982 14632 11034 14684
rect 11046 14632 11098 14684
rect 11110 14632 11162 14684
rect 11174 14632 11226 14684
rect 20982 14632 21034 14684
rect 21046 14632 21098 14684
rect 21110 14632 21162 14684
rect 21174 14632 21226 14684
rect 19432 14573 19484 14582
rect 19432 14539 19441 14573
rect 19441 14539 19475 14573
rect 19475 14539 19484 14573
rect 19432 14530 19484 14539
rect 19524 14530 19576 14582
rect 24032 14394 24084 14446
rect 19708 14326 19760 14378
rect 19892 14369 19944 14378
rect 19892 14335 19901 14369
rect 19901 14335 19935 14369
rect 19935 14335 19944 14369
rect 19892 14326 19944 14335
rect 19984 14369 20036 14378
rect 19984 14335 19993 14369
rect 19993 14335 20027 14369
rect 20027 14335 20036 14369
rect 19984 14326 20036 14335
rect 23572 14190 23624 14242
rect 5982 14088 6034 14140
rect 6046 14088 6098 14140
rect 6110 14088 6162 14140
rect 6174 14088 6226 14140
rect 15982 14088 16034 14140
rect 16046 14088 16098 14140
rect 16110 14088 16162 14140
rect 16174 14088 16226 14140
rect 25982 14088 26034 14140
rect 26046 14088 26098 14140
rect 26110 14088 26162 14140
rect 26174 14088 26226 14140
rect 19524 14029 19576 14038
rect 19524 13995 19533 14029
rect 19533 13995 19567 14029
rect 19567 13995 19576 14029
rect 19524 13986 19576 13995
rect 19984 13986 20036 14038
rect 24032 14029 24084 14038
rect 24032 13995 24041 14029
rect 24041 13995 24075 14029
rect 24075 13995 24084 14029
rect 24032 13986 24084 13995
rect 19708 13782 19760 13834
rect 10982 13544 11034 13596
rect 11046 13544 11098 13596
rect 11110 13544 11162 13596
rect 11174 13544 11226 13596
rect 20982 13544 21034 13596
rect 21046 13544 21098 13596
rect 21110 13544 21162 13596
rect 21174 13544 21226 13596
rect 13544 13485 13596 13494
rect 13544 13451 13553 13485
rect 13553 13451 13587 13485
rect 13587 13451 13596 13485
rect 13544 13442 13596 13451
rect 19248 13442 19300 13494
rect 1492 13306 1544 13358
rect 3240 13306 3292 13358
rect 3884 13306 3936 13358
rect 13820 13306 13872 13358
rect 19524 13349 19576 13358
rect 19524 13315 19533 13349
rect 19533 13315 19567 13349
rect 19567 13315 19576 13349
rect 19524 13306 19576 13315
rect 13912 13170 13964 13222
rect 14096 13281 14148 13290
rect 14096 13247 14105 13281
rect 14105 13247 14139 13281
rect 14139 13247 14148 13281
rect 14096 13238 14148 13247
rect 19156 13238 19208 13290
rect 19616 13281 19668 13290
rect 19616 13247 19625 13281
rect 19625 13247 19659 13281
rect 19659 13247 19668 13281
rect 19616 13238 19668 13247
rect 19984 13238 20036 13290
rect 1860 13102 1912 13154
rect 5982 13000 6034 13052
rect 6046 13000 6098 13052
rect 6110 13000 6162 13052
rect 6174 13000 6226 13052
rect 15982 13000 16034 13052
rect 16046 13000 16098 13052
rect 16110 13000 16162 13052
rect 16174 13000 16226 13052
rect 25982 13000 26034 13052
rect 26046 13000 26098 13052
rect 26110 13000 26162 13052
rect 26174 13000 26226 13052
rect 14096 12898 14148 12950
rect 19984 12941 20036 12950
rect 19984 12907 19993 12941
rect 19993 12907 20027 12941
rect 20027 12907 20036 12941
rect 19984 12898 20036 12907
rect 19524 12762 19576 12814
rect 1400 12737 1452 12746
rect 1400 12703 1409 12737
rect 1409 12703 1443 12737
rect 1443 12703 1452 12737
rect 1400 12694 1452 12703
rect 19156 12737 19208 12746
rect 19156 12703 19165 12737
rect 19165 12703 19199 12737
rect 19199 12703 19208 12737
rect 19156 12694 19208 12703
rect 13820 12626 13872 12678
rect 1676 12558 1728 12610
rect 13912 12601 13964 12610
rect 13912 12567 13921 12601
rect 13921 12567 13955 12601
rect 13955 12567 13964 12601
rect 13912 12558 13964 12567
rect 10982 12456 11034 12508
rect 11046 12456 11098 12508
rect 11110 12456 11162 12508
rect 11174 12456 11226 12508
rect 20982 12456 21034 12508
rect 21046 12456 21098 12508
rect 21110 12456 21162 12508
rect 21174 12456 21226 12508
rect 1492 12354 1544 12406
rect 8300 12354 8352 12406
rect 13728 12354 13780 12406
rect 8668 12218 8720 12270
rect 13084 12218 13136 12270
rect 8484 12193 8536 12202
rect 8484 12159 8493 12193
rect 8493 12159 8527 12193
rect 8527 12159 8536 12193
rect 8484 12150 8536 12159
rect 13544 12193 13596 12202
rect 13544 12159 13553 12193
rect 13553 12159 13587 12193
rect 13587 12159 13596 12193
rect 13544 12150 13596 12159
rect 7932 12125 7984 12134
rect 7932 12091 7941 12125
rect 7941 12091 7975 12125
rect 7975 12091 7984 12125
rect 7932 12082 7984 12091
rect 13452 12082 13504 12134
rect 12072 12014 12124 12066
rect 5982 11912 6034 11964
rect 6046 11912 6098 11964
rect 6110 11912 6162 11964
rect 6174 11912 6226 11964
rect 15982 11912 16034 11964
rect 16046 11912 16098 11964
rect 16110 11912 16162 11964
rect 16174 11912 16226 11964
rect 25982 11912 26034 11964
rect 26046 11912 26098 11964
rect 26110 11912 26162 11964
rect 26174 11912 26226 11964
rect 8484 11810 8536 11862
rect 11980 11853 12032 11862
rect 11980 11819 11989 11853
rect 11989 11819 12023 11853
rect 12023 11819 12032 11853
rect 11980 11810 12032 11819
rect 13544 11810 13596 11862
rect 24400 11810 24452 11862
rect 13084 11742 13136 11794
rect 12072 11674 12124 11726
rect 13452 11674 13504 11726
rect 1584 11606 1636 11658
rect 11980 11606 12032 11658
rect 12624 11649 12676 11658
rect 12624 11615 12633 11649
rect 12633 11615 12667 11649
rect 12667 11615 12676 11649
rect 12624 11606 12676 11615
rect 24400 11606 24452 11658
rect 2136 11470 2188 11522
rect 8300 11513 8352 11522
rect 8300 11479 8309 11513
rect 8309 11479 8343 11513
rect 8343 11479 8352 11513
rect 8300 11470 8352 11479
rect 8668 11513 8720 11522
rect 8668 11479 8677 11513
rect 8677 11479 8711 11513
rect 8711 11479 8720 11513
rect 8668 11470 8720 11479
rect 12164 11470 12216 11522
rect 24124 11513 24176 11522
rect 24124 11479 24133 11513
rect 24133 11479 24167 11513
rect 24167 11479 24176 11513
rect 24124 11470 24176 11479
rect 10982 11368 11034 11420
rect 11046 11368 11098 11420
rect 11110 11368 11162 11420
rect 11174 11368 11226 11420
rect 20982 11368 21034 11420
rect 21046 11368 21098 11420
rect 21110 11368 21162 11420
rect 21174 11368 21226 11420
rect 8668 11266 8720 11318
rect 12164 11309 12216 11318
rect 12164 11275 12173 11309
rect 12173 11275 12207 11309
rect 12207 11275 12216 11309
rect 12164 11266 12216 11275
rect 8116 11241 8168 11250
rect 8116 11207 8125 11241
rect 8125 11207 8159 11241
rect 8159 11207 8168 11241
rect 8116 11198 8168 11207
rect 2044 11130 2096 11182
rect 7196 11130 7248 11182
rect 23940 11173 23992 11182
rect 23940 11139 23949 11173
rect 23949 11139 23983 11173
rect 23983 11139 23992 11173
rect 23940 11130 23992 11139
rect 7380 11062 7432 11114
rect 8300 11105 8352 11114
rect 8300 11071 8309 11105
rect 8309 11071 8343 11105
rect 8343 11071 8352 11105
rect 8300 11062 8352 11071
rect 1952 10994 2004 11046
rect 24860 10994 24912 11046
rect 5982 10824 6034 10876
rect 6046 10824 6098 10876
rect 6110 10824 6162 10876
rect 6174 10824 6226 10876
rect 15982 10824 16034 10876
rect 16046 10824 16098 10876
rect 16110 10824 16162 10876
rect 16174 10824 16226 10876
rect 25982 10824 26034 10876
rect 26046 10824 26098 10876
rect 26110 10824 26162 10876
rect 26174 10824 26226 10876
rect 2044 10765 2096 10774
rect 2044 10731 2053 10765
rect 2053 10731 2087 10765
rect 2087 10731 2096 10765
rect 2044 10722 2096 10731
rect 2412 10765 2464 10774
rect 2412 10731 2421 10765
rect 2421 10731 2455 10765
rect 2455 10731 2464 10765
rect 2412 10722 2464 10731
rect 7104 10765 7156 10774
rect 7104 10731 7113 10765
rect 7113 10731 7147 10765
rect 7147 10731 7156 10765
rect 7104 10722 7156 10731
rect 8208 10722 8260 10774
rect 8300 10722 8352 10774
rect 23940 10765 23992 10774
rect 23940 10731 23949 10765
rect 23949 10731 23983 10765
rect 23983 10731 23992 10765
rect 23940 10722 23992 10731
rect 8576 10629 8628 10638
rect 8576 10595 8585 10629
rect 8585 10595 8619 10629
rect 8619 10595 8628 10629
rect 8576 10586 8628 10595
rect 2412 10518 2464 10570
rect 8300 10493 8352 10502
rect 8300 10459 8309 10493
rect 8309 10459 8343 10493
rect 8343 10459 8352 10493
rect 8300 10450 8352 10459
rect 1768 10382 1820 10434
rect 7380 10425 7432 10434
rect 7380 10391 7389 10425
rect 7389 10391 7423 10425
rect 7423 10391 7432 10425
rect 7380 10382 7432 10391
rect 7840 10425 7892 10434
rect 7840 10391 7849 10425
rect 7849 10391 7883 10425
rect 7883 10391 7892 10425
rect 8392 10425 8444 10434
rect 7840 10382 7892 10391
rect 8392 10391 8401 10425
rect 8401 10391 8435 10425
rect 8435 10391 8444 10425
rect 8392 10382 8444 10391
rect 10982 10280 11034 10332
rect 11046 10280 11098 10332
rect 11110 10280 11162 10332
rect 11174 10280 11226 10332
rect 20982 10280 21034 10332
rect 21046 10280 21098 10332
rect 21110 10280 21162 10332
rect 21174 10280 21226 10332
rect 8300 10178 8352 10230
rect 8576 10178 8628 10230
rect 2228 10042 2280 10094
rect 1584 9881 1636 9890
rect 1584 9847 1593 9881
rect 1593 9847 1627 9881
rect 1627 9847 1636 9881
rect 1584 9838 1636 9847
rect 5982 9736 6034 9788
rect 6046 9736 6098 9788
rect 6110 9736 6162 9788
rect 6174 9736 6226 9788
rect 15982 9736 16034 9788
rect 16046 9736 16098 9788
rect 16110 9736 16162 9788
rect 16174 9736 16226 9788
rect 25982 9736 26034 9788
rect 26046 9736 26098 9788
rect 26110 9736 26162 9788
rect 26174 9736 26226 9788
rect 2228 9634 2280 9686
rect 2504 9566 2556 9618
rect 23940 9473 23992 9482
rect 23940 9439 23949 9473
rect 23949 9439 23983 9473
rect 23983 9439 23992 9473
rect 23940 9430 23992 9439
rect 1584 9337 1636 9346
rect 1584 9303 1593 9337
rect 1593 9303 1627 9337
rect 1627 9303 1636 9337
rect 1584 9294 1636 9303
rect 24124 9337 24176 9346
rect 24124 9303 24133 9337
rect 24133 9303 24167 9337
rect 24167 9303 24176 9337
rect 24124 9294 24176 9303
rect 10982 9192 11034 9244
rect 11046 9192 11098 9244
rect 11110 9192 11162 9244
rect 11174 9192 11226 9244
rect 20982 9192 21034 9244
rect 21046 9192 21098 9244
rect 21110 9192 21162 9244
rect 21174 9192 21226 9244
rect 1400 8997 1452 9006
rect 1400 8963 1409 8997
rect 1409 8963 1443 8997
rect 1443 8963 1452 8997
rect 1400 8954 1452 8963
rect 23940 8997 23992 9006
rect 23940 8963 23949 8997
rect 23949 8963 23983 8997
rect 23983 8963 23992 8997
rect 23940 8954 23992 8963
rect 1400 8750 1452 8802
rect 1952 8750 2004 8802
rect 2688 8750 2740 8802
rect 24124 8793 24176 8802
rect 24124 8759 24133 8793
rect 24133 8759 24167 8793
rect 24167 8759 24176 8793
rect 24124 8750 24176 8759
rect 5982 8648 6034 8700
rect 6046 8648 6098 8700
rect 6110 8648 6162 8700
rect 6174 8648 6226 8700
rect 15982 8648 16034 8700
rect 16046 8648 16098 8700
rect 16110 8648 16162 8700
rect 16174 8648 16226 8700
rect 25982 8648 26034 8700
rect 26046 8648 26098 8700
rect 26110 8648 26162 8700
rect 26174 8648 26226 8700
rect 1492 8546 1544 8598
rect 23756 8589 23808 8598
rect 23756 8555 23765 8589
rect 23765 8555 23799 8589
rect 23799 8555 23808 8589
rect 23756 8546 23808 8555
rect 23940 8546 23992 8598
rect 23480 8478 23532 8530
rect 23756 8342 23808 8394
rect 10982 8104 11034 8156
rect 11046 8104 11098 8156
rect 11110 8104 11162 8156
rect 11174 8104 11226 8156
rect 20982 8104 21034 8156
rect 21046 8104 21098 8156
rect 21110 8104 21162 8156
rect 21174 8104 21226 8156
rect 24124 8045 24176 8054
rect 24124 8011 24133 8045
rect 24133 8011 24167 8045
rect 24167 8011 24176 8045
rect 24124 8002 24176 8011
rect 23940 7909 23992 7918
rect 23940 7875 23949 7909
rect 23949 7875 23983 7909
rect 23983 7875 23992 7909
rect 23940 7866 23992 7875
rect 5982 7560 6034 7612
rect 6046 7560 6098 7612
rect 6110 7560 6162 7612
rect 6174 7560 6226 7612
rect 15982 7560 16034 7612
rect 16046 7560 16098 7612
rect 16110 7560 16162 7612
rect 16174 7560 16226 7612
rect 25982 7560 26034 7612
rect 26046 7560 26098 7612
rect 26110 7560 26162 7612
rect 26174 7560 26226 7612
rect 22468 7501 22520 7510
rect 22468 7467 22477 7501
rect 22477 7467 22511 7501
rect 22511 7467 22520 7501
rect 22468 7458 22520 7467
rect 22928 7501 22980 7510
rect 22928 7467 22937 7501
rect 22937 7467 22971 7501
rect 22971 7467 22980 7501
rect 22928 7458 22980 7467
rect 23940 7501 23992 7510
rect 23940 7467 23949 7501
rect 23949 7467 23983 7501
rect 23983 7467 23992 7501
rect 23940 7458 23992 7467
rect 18604 7433 18656 7442
rect 18604 7399 18613 7433
rect 18613 7399 18647 7433
rect 18647 7399 18656 7433
rect 18604 7390 18656 7399
rect 13084 7297 13136 7306
rect 13084 7263 13093 7297
rect 13093 7263 13127 7297
rect 13127 7263 13136 7297
rect 13084 7254 13136 7263
rect 18420 7297 18472 7306
rect 18420 7263 18429 7297
rect 18429 7263 18463 7297
rect 18463 7263 18472 7297
rect 18420 7254 18472 7263
rect 22928 7254 22980 7306
rect 13268 7161 13320 7170
rect 13268 7127 13277 7161
rect 13277 7127 13311 7161
rect 13311 7127 13320 7161
rect 13268 7118 13320 7127
rect 10982 7016 11034 7068
rect 11046 7016 11098 7068
rect 11110 7016 11162 7068
rect 11174 7016 11226 7068
rect 20982 7016 21034 7068
rect 21046 7016 21098 7068
rect 21110 7016 21162 7068
rect 21174 7016 21226 7068
rect 1308 6846 1360 6898
rect 1860 6846 1912 6898
rect 14740 6821 14792 6830
rect 14740 6787 14749 6821
rect 14749 6787 14783 6821
rect 14783 6787 14792 6821
rect 14740 6778 14792 6787
rect 24032 6778 24084 6830
rect 14924 6685 14976 6694
rect 14924 6651 14933 6685
rect 14933 6651 14967 6685
rect 14967 6651 14976 6685
rect 14924 6642 14976 6651
rect 24124 6685 24176 6694
rect 24124 6651 24133 6685
rect 24133 6651 24167 6685
rect 24167 6651 24176 6685
rect 24124 6642 24176 6651
rect 5982 6472 6034 6524
rect 6046 6472 6098 6524
rect 6110 6472 6162 6524
rect 6174 6472 6226 6524
rect 15982 6472 16034 6524
rect 16046 6472 16098 6524
rect 16110 6472 16162 6524
rect 16174 6472 16226 6524
rect 25982 6472 26034 6524
rect 26046 6472 26098 6524
rect 26110 6472 26162 6524
rect 26174 6472 26226 6524
rect 14740 6413 14792 6422
rect 14740 6379 14749 6413
rect 14749 6379 14783 6413
rect 14783 6379 14792 6413
rect 14740 6370 14792 6379
rect 24032 6413 24084 6422
rect 24032 6379 24041 6413
rect 24041 6379 24075 6413
rect 24075 6379 24084 6413
rect 24032 6370 24084 6379
rect 10982 5928 11034 5980
rect 11046 5928 11098 5980
rect 11110 5928 11162 5980
rect 11174 5928 11226 5980
rect 20982 5928 21034 5980
rect 21046 5928 21098 5980
rect 21110 5928 21162 5980
rect 21174 5928 21226 5980
rect 13084 5869 13136 5878
rect 13084 5835 13093 5869
rect 13093 5835 13127 5869
rect 13127 5835 13136 5869
rect 13084 5826 13136 5835
rect 4160 5733 4212 5742
rect 4160 5699 4169 5733
rect 4169 5699 4203 5733
rect 4203 5699 4212 5733
rect 4160 5690 4212 5699
rect 13636 5690 13688 5742
rect 4344 5597 4396 5606
rect 4344 5563 4353 5597
rect 4353 5563 4387 5597
rect 4387 5563 4396 5597
rect 4344 5554 4396 5563
rect 5982 5384 6034 5436
rect 6046 5384 6098 5436
rect 6110 5384 6162 5436
rect 6174 5384 6226 5436
rect 15982 5384 16034 5436
rect 16046 5384 16098 5436
rect 16110 5384 16162 5436
rect 16174 5384 16226 5436
rect 25982 5384 26034 5436
rect 26046 5384 26098 5436
rect 26110 5384 26162 5436
rect 26174 5384 26226 5436
rect 4160 5282 4212 5334
rect 13636 5325 13688 5334
rect 13636 5291 13645 5325
rect 13645 5291 13679 5325
rect 13679 5291 13688 5325
rect 13636 5282 13688 5291
rect 12624 5121 12676 5130
rect 12624 5087 12633 5121
rect 12633 5087 12667 5121
rect 12667 5087 12676 5121
rect 12624 5078 12676 5087
rect 24768 5282 24820 5334
rect 12808 4985 12860 4994
rect 12808 4951 12817 4985
rect 12817 4951 12851 4985
rect 12851 4951 12860 4985
rect 12808 4942 12860 4951
rect 24124 4985 24176 4994
rect 24124 4951 24133 4985
rect 24133 4951 24167 4985
rect 24167 4951 24176 4985
rect 24124 4942 24176 4951
rect 10982 4840 11034 4892
rect 11046 4840 11098 4892
rect 11110 4840 11162 4892
rect 11174 4840 11226 4892
rect 20982 4840 21034 4892
rect 21046 4840 21098 4892
rect 21110 4840 21162 4892
rect 21174 4840 21226 4892
rect 15568 4645 15620 4654
rect 15568 4611 15577 4645
rect 15577 4611 15611 4645
rect 15611 4611 15620 4645
rect 15568 4602 15620 4611
rect 20444 4645 20496 4654
rect 20444 4611 20453 4645
rect 20453 4611 20487 4645
rect 20487 4611 20496 4645
rect 20444 4602 20496 4611
rect 15752 4509 15804 4518
rect 15752 4475 15761 4509
rect 15761 4475 15795 4509
rect 15795 4475 15804 4509
rect 15752 4466 15804 4475
rect 20628 4509 20680 4518
rect 20628 4475 20637 4509
rect 20637 4475 20671 4509
rect 20671 4475 20680 4509
rect 20628 4466 20680 4475
rect 5982 4296 6034 4348
rect 6046 4296 6098 4348
rect 6110 4296 6162 4348
rect 6174 4296 6226 4348
rect 15982 4296 16034 4348
rect 16046 4296 16098 4348
rect 16110 4296 16162 4348
rect 16174 4296 16226 4348
rect 25982 4296 26034 4348
rect 26046 4296 26098 4348
rect 26110 4296 26162 4348
rect 26174 4296 26226 4348
rect 15568 4237 15620 4246
rect 15568 4203 15577 4237
rect 15577 4203 15611 4237
rect 15611 4203 15620 4237
rect 15568 4194 15620 4203
rect 20444 4237 20496 4246
rect 20444 4203 20453 4237
rect 20453 4203 20487 4237
rect 20487 4203 20496 4237
rect 20444 4194 20496 4203
rect 21456 4101 21508 4110
rect 21456 4067 21465 4101
rect 21465 4067 21499 4101
rect 21499 4067 21508 4101
rect 21456 4058 21508 4067
rect 23940 4033 23992 4042
rect 23940 3999 23949 4033
rect 23949 3999 23983 4033
rect 23983 3999 23992 4033
rect 23940 3990 23992 3999
rect 20720 3854 20772 3906
rect 24124 3897 24176 3906
rect 24124 3863 24133 3897
rect 24133 3863 24167 3897
rect 24167 3863 24176 3897
rect 24124 3854 24176 3863
rect 10982 3752 11034 3804
rect 11046 3752 11098 3804
rect 11110 3752 11162 3804
rect 11174 3752 11226 3804
rect 20982 3752 21034 3804
rect 21046 3752 21098 3804
rect 21110 3752 21162 3804
rect 21174 3752 21226 3804
rect 23848 3514 23900 3566
rect 24676 3514 24728 3566
rect 24124 3421 24176 3430
rect 24124 3387 24133 3421
rect 24133 3387 24167 3421
rect 24167 3387 24176 3421
rect 24124 3378 24176 3387
rect 5982 3208 6034 3260
rect 6046 3208 6098 3260
rect 6110 3208 6162 3260
rect 6174 3208 6226 3260
rect 15982 3208 16034 3260
rect 16046 3208 16098 3260
rect 16110 3208 16162 3260
rect 16174 3208 16226 3260
rect 25982 3208 26034 3260
rect 26046 3208 26098 3260
rect 26110 3208 26162 3260
rect 26174 3208 26226 3260
rect 1952 3149 2004 3158
rect 1952 3115 1961 3149
rect 1961 3115 1995 3149
rect 1995 3115 2004 3149
rect 1952 3106 2004 3115
rect 23848 3149 23900 3158
rect 23848 3115 23857 3149
rect 23857 3115 23891 3149
rect 23891 3115 23900 3149
rect 23848 3106 23900 3115
rect 1952 2902 2004 2954
rect 23940 2945 23992 2954
rect 23940 2911 23949 2945
rect 23949 2911 23983 2945
rect 23983 2911 23992 2945
rect 23940 2902 23992 2911
rect 9496 2766 9548 2818
rect 24860 2766 24912 2818
rect 10982 2664 11034 2716
rect 11046 2664 11098 2716
rect 11110 2664 11162 2716
rect 11174 2664 11226 2716
rect 20982 2664 21034 2716
rect 21046 2664 21098 2716
rect 21110 2664 21162 2716
rect 21174 2664 21226 2716
rect 24216 2605 24268 2614
rect 24216 2571 24225 2605
rect 24225 2571 24259 2605
rect 24259 2571 24268 2605
rect 24216 2562 24268 2571
rect 24032 2469 24084 2478
rect 24032 2435 24041 2469
rect 24041 2435 24075 2469
rect 24075 2435 24084 2469
rect 24032 2426 24084 2435
rect 25136 2469 25188 2478
rect 25136 2435 25145 2469
rect 25145 2435 25179 2469
rect 25179 2435 25188 2469
rect 25136 2426 25188 2435
rect 2044 2401 2096 2410
rect 2044 2367 2053 2401
rect 2053 2367 2087 2401
rect 2087 2367 2096 2401
rect 2044 2358 2096 2367
rect 1584 2265 1636 2274
rect 1584 2231 1593 2265
rect 1593 2231 1627 2265
rect 1627 2231 1636 2265
rect 1584 2222 1636 2231
rect 25320 2265 25372 2274
rect 25320 2231 25329 2265
rect 25329 2231 25363 2265
rect 25363 2231 25372 2265
rect 25320 2222 25372 2231
rect 5982 2120 6034 2172
rect 6046 2120 6098 2172
rect 6110 2120 6162 2172
rect 6174 2120 6226 2172
rect 15982 2120 16034 2172
rect 16046 2120 16098 2172
rect 16110 2120 16162 2172
rect 16174 2120 16226 2172
rect 25982 2120 26034 2172
rect 26046 2120 26098 2172
rect 26110 2120 26162 2172
rect 26174 2120 26226 2172
<< metal2 >>
rect 3698 23490 3754 23970
rect 3882 23594 3938 23603
rect 3882 23529 3938 23538
rect 3330 23050 3386 23059
rect 3330 22985 3386 22994
rect 3146 21282 3202 21291
rect 3146 21217 3202 21226
rect 3160 18872 3188 21217
rect 3148 18866 3200 18872
rect 3148 18808 3200 18814
rect 3238 18834 3294 18843
rect 3238 18769 3294 18778
rect 2870 18290 2926 18299
rect 2870 18225 2926 18234
rect 1398 15298 1454 15307
rect 1398 15233 1454 15242
rect 1412 12752 1440 15233
rect 1582 14074 1638 14083
rect 1582 14009 1638 14018
rect 1490 13394 1546 13403
rect 1490 13329 1492 13338
rect 1544 13329 1546 13338
rect 1492 13300 1544 13306
rect 1400 12746 1452 12752
rect 1400 12688 1452 12694
rect 1504 12412 1532 13300
rect 1492 12406 1544 12412
rect 1492 12348 1544 12354
rect 1596 11664 1624 14009
rect 1860 13154 1912 13160
rect 1860 13096 1912 13102
rect 1676 12610 1728 12616
rect 1676 12552 1728 12558
rect 1584 11658 1636 11664
rect 1584 11600 1636 11606
rect 1398 9994 1454 10003
rect 1398 9929 1454 9938
rect 1412 9012 1440 9929
rect 1584 9890 1636 9896
rect 1582 9858 1584 9867
rect 1636 9858 1638 9867
rect 1582 9793 1638 9802
rect 1584 9346 1636 9352
rect 1584 9288 1636 9294
rect 1400 9006 1452 9012
rect 1400 8948 1452 8954
rect 1412 8892 1440 8948
rect 1412 8864 1532 8892
rect 1400 8802 1452 8808
rect 1400 8744 1452 8750
rect 1308 6898 1360 6904
rect 1308 6840 1360 6846
rect 1320 6331 1348 6840
rect 1306 6322 1362 6331
rect 1306 6257 1362 6266
rect 1412 347 1440 8744
rect 1504 8604 1532 8864
rect 1492 8598 1544 8604
rect 1492 8540 1544 8546
rect 1596 2364 1624 9288
rect 1688 2931 1716 12552
rect 1768 10434 1820 10440
rect 1768 10376 1820 10382
rect 1674 2922 1730 2931
rect 1674 2857 1730 2866
rect 1780 2659 1808 10376
rect 1872 6904 1900 13096
rect 2778 12850 2834 12859
rect 2778 12785 2834 12794
rect 2226 12714 2282 12723
rect 2226 12649 2282 12658
rect 2136 11522 2188 11528
rect 2136 11464 2188 11470
rect 2042 11218 2098 11227
rect 2042 11153 2044 11162
rect 2096 11153 2098 11162
rect 2044 11124 2096 11130
rect 1952 11046 2004 11052
rect 1952 10988 2004 10994
rect 1964 8892 1992 10988
rect 2056 10780 2084 11124
rect 2044 10774 2096 10780
rect 2044 10716 2096 10722
rect 1964 8864 2084 8892
rect 1952 8802 2004 8808
rect 1952 8744 2004 8750
rect 1860 6898 1912 6904
rect 1860 6840 1912 6846
rect 1964 3164 1992 8744
rect 1952 3158 2004 3164
rect 1952 3100 2004 3106
rect 1964 2960 1992 3100
rect 1952 2954 2004 2960
rect 1952 2896 2004 2902
rect 1766 2650 1822 2659
rect 1766 2585 1822 2594
rect 2056 2523 2084 8864
rect 2042 2514 2098 2523
rect 2042 2449 2098 2458
rect 2044 2410 2096 2416
rect 1504 2336 1624 2364
rect 2042 2378 2044 2387
rect 2096 2378 2098 2387
rect 1504 1435 1532 2336
rect 2042 2313 2098 2322
rect 1584 2274 1636 2280
rect 1584 2216 1636 2222
rect 1490 1426 1546 1435
rect 1490 1361 1546 1370
rect 1596 891 1624 2216
rect 2148 1435 2176 11464
rect 2240 10100 2268 12649
rect 2410 11490 2466 11499
rect 2410 11425 2466 11434
rect 2424 10780 2452 11425
rect 2502 11354 2558 11363
rect 2502 11289 2558 11298
rect 2412 10774 2464 10780
rect 2412 10716 2464 10722
rect 2424 10576 2452 10716
rect 2412 10570 2464 10576
rect 2412 10512 2464 10518
rect 2228 10094 2280 10100
rect 2228 10036 2280 10042
rect 2240 9692 2268 10036
rect 2228 9686 2280 9692
rect 2228 9628 2280 9634
rect 2516 9624 2544 11289
rect 2792 9708 2820 12785
rect 2884 11771 2912 18225
rect 3054 15842 3110 15851
rect 3054 15777 3110 15786
rect 2870 11762 2926 11771
rect 2870 11697 2926 11706
rect 2700 9680 2820 9708
rect 2504 9618 2556 9624
rect 2504 9560 2556 9566
rect 2700 8808 2728 9680
rect 3068 9436 3096 15777
rect 3252 13364 3280 18769
rect 3344 18299 3372 22985
rect 3514 22370 3570 22379
rect 3514 22305 3570 22314
rect 3422 21826 3478 21835
rect 3422 21761 3478 21770
rect 3436 20776 3464 21761
rect 3424 20770 3476 20776
rect 3424 20712 3476 20718
rect 3330 18290 3386 18299
rect 3330 18225 3386 18234
rect 3528 17755 3556 22305
rect 3606 20058 3662 20067
rect 3606 19993 3662 20002
rect 3514 17746 3570 17755
rect 3514 17681 3570 17690
rect 3330 17610 3386 17619
rect 3330 17545 3386 17554
rect 3240 13358 3292 13364
rect 3240 13300 3292 13306
rect 3238 13258 3294 13267
rect 3238 13193 3294 13202
rect 3146 12306 3202 12315
rect 3146 12241 3202 12250
rect 3160 10275 3188 12241
rect 3252 12179 3280 13193
rect 3344 12428 3372 17545
rect 3514 17066 3570 17075
rect 3514 17001 3570 17010
rect 3422 14618 3478 14627
rect 3422 14553 3478 14562
rect 3436 13267 3464 14553
rect 3422 13258 3478 13267
rect 3422 13193 3478 13202
rect 3344 12400 3464 12428
rect 3330 12306 3386 12315
rect 3330 12241 3386 12250
rect 3238 12170 3294 12179
rect 3238 12105 3294 12114
rect 3344 11635 3372 12241
rect 3330 11626 3386 11635
rect 3330 11561 3386 11570
rect 3146 10266 3202 10275
rect 3146 10201 3202 10210
rect 3436 9595 3464 12400
rect 3422 9586 3478 9595
rect 3422 9521 3478 9530
rect 3068 9408 3464 9436
rect 2688 8802 2740 8808
rect 2688 8744 2740 8750
rect 3436 4019 3464 9408
rect 3528 5243 3556 17001
rect 3620 7283 3648 19993
rect 3712 18979 3740 23490
rect 3790 19378 3846 19387
rect 3790 19313 3846 19322
rect 3698 18970 3754 18979
rect 3698 18905 3754 18914
rect 3700 18866 3752 18872
rect 3700 18808 3752 18814
rect 3712 9459 3740 18808
rect 3698 9450 3754 9459
rect 3698 9385 3754 9394
rect 3804 7419 3832 19313
rect 3896 18843 3924 23529
rect 11150 23490 11206 23970
rect 18694 23490 18750 23970
rect 24766 23594 24822 23603
rect 24766 23529 24822 23538
rect 5956 21758 6252 21778
rect 6012 21756 6036 21758
rect 6092 21756 6116 21758
rect 6172 21756 6196 21758
rect 6034 21704 6036 21756
rect 6098 21704 6110 21756
rect 6172 21704 6174 21756
rect 6012 21702 6036 21704
rect 6092 21702 6116 21704
rect 6172 21702 6196 21704
rect 5956 21682 6252 21702
rect 11164 21404 11192 23490
rect 15956 21758 16252 21778
rect 16012 21756 16036 21758
rect 16092 21756 16116 21758
rect 16172 21756 16196 21758
rect 16034 21704 16036 21756
rect 16098 21704 16110 21756
rect 16172 21704 16174 21756
rect 16012 21702 16036 21704
rect 16092 21702 16116 21704
rect 16172 21702 16196 21704
rect 15956 21682 16252 21702
rect 11164 21376 11376 21404
rect 10956 21214 11252 21234
rect 11012 21212 11036 21214
rect 11092 21212 11116 21214
rect 11172 21212 11196 21214
rect 11034 21160 11036 21212
rect 11098 21160 11110 21212
rect 11172 21160 11174 21212
rect 11012 21158 11036 21160
rect 11092 21158 11116 21160
rect 11172 21158 11196 21160
rect 10956 21138 11252 21158
rect 5956 20670 6252 20690
rect 6012 20668 6036 20670
rect 6092 20668 6116 20670
rect 6172 20668 6196 20670
rect 6034 20616 6036 20668
rect 6098 20616 6110 20668
rect 6172 20616 6174 20668
rect 6012 20614 6036 20616
rect 6092 20614 6116 20616
rect 6172 20614 6196 20616
rect 3974 20602 4030 20611
rect 5956 20594 6252 20614
rect 3974 20537 4030 20546
rect 3882 18834 3938 18843
rect 3882 18769 3938 18778
rect 3884 13358 3936 13364
rect 3884 13300 3936 13306
rect 3896 7827 3924 13300
rect 3988 9051 4016 20537
rect 10956 20126 11252 20146
rect 11012 20124 11036 20126
rect 11092 20124 11116 20126
rect 11172 20124 11196 20126
rect 11034 20072 11036 20124
rect 11098 20072 11110 20124
rect 11172 20072 11174 20124
rect 11012 20070 11036 20072
rect 11092 20070 11116 20072
rect 11172 20070 11196 20072
rect 10956 20050 11252 20070
rect 5956 19582 6252 19602
rect 6012 19580 6036 19582
rect 6092 19580 6116 19582
rect 6172 19580 6196 19582
rect 6034 19528 6036 19580
rect 6098 19528 6110 19580
rect 6172 19528 6174 19580
rect 6012 19526 6036 19528
rect 6092 19526 6116 19528
rect 6172 19526 6196 19528
rect 5956 19506 6252 19526
rect 11348 19387 11376 21376
rect 15956 20670 16252 20690
rect 16012 20668 16036 20670
rect 16092 20668 16116 20670
rect 16172 20668 16196 20670
rect 16034 20616 16036 20668
rect 16098 20616 16110 20668
rect 16172 20616 16174 20668
rect 16012 20614 16036 20616
rect 16092 20614 16116 20616
rect 16172 20614 16196 20616
rect 15956 20594 16252 20614
rect 15956 19582 16252 19602
rect 16012 19580 16036 19582
rect 16092 19580 16116 19582
rect 16172 19580 16196 19582
rect 16034 19528 16036 19580
rect 16098 19528 16110 19580
rect 16172 19528 16174 19580
rect 16012 19526 16036 19528
rect 16092 19526 16116 19528
rect 16172 19526 16196 19528
rect 15956 19506 16252 19526
rect 8850 19378 8906 19387
rect 8850 19313 8906 19322
rect 11334 19378 11390 19387
rect 11334 19313 11390 19322
rect 7010 18970 7066 18979
rect 7010 18905 7066 18914
rect 8574 18970 8630 18979
rect 8574 18905 8630 18914
rect 5956 18494 6252 18514
rect 6012 18492 6036 18494
rect 6092 18492 6116 18494
rect 6172 18492 6196 18494
rect 6034 18440 6036 18492
rect 6098 18440 6110 18492
rect 6172 18440 6174 18492
rect 6012 18438 6036 18440
rect 6092 18438 6116 18440
rect 6172 18438 6196 18440
rect 5956 18418 6252 18438
rect 5956 17406 6252 17426
rect 6012 17404 6036 17406
rect 6092 17404 6116 17406
rect 6172 17404 6196 17406
rect 6034 17352 6036 17404
rect 6098 17352 6110 17404
rect 6172 17352 6174 17404
rect 6012 17350 6036 17352
rect 6092 17350 6116 17352
rect 6172 17350 6196 17352
rect 5956 17330 6252 17350
rect 4066 16386 4122 16395
rect 4066 16321 4122 16330
rect 3974 9042 4030 9051
rect 3974 8977 4030 8986
rect 3882 7818 3938 7827
rect 3882 7753 3938 7762
rect 4080 7668 4108 16321
rect 5956 16318 6252 16338
rect 6012 16316 6036 16318
rect 6092 16316 6116 16318
rect 6172 16316 6196 16318
rect 6034 16264 6036 16316
rect 6098 16264 6110 16316
rect 6172 16264 6174 16316
rect 6012 16262 6036 16264
rect 6092 16262 6116 16264
rect 6172 16262 6196 16264
rect 5956 16242 6252 16262
rect 7024 16220 7052 18905
rect 8588 18804 8616 18905
rect 8864 18872 8892 19313
rect 10956 19038 11252 19058
rect 11012 19036 11036 19038
rect 11092 19036 11116 19038
rect 11172 19036 11196 19038
rect 11034 18984 11036 19036
rect 11098 18984 11110 19036
rect 11172 18984 11174 19036
rect 11012 18982 11036 18984
rect 11092 18982 11116 18984
rect 11172 18982 11196 18984
rect 10956 18962 11252 18982
rect 18708 18979 18736 23490
rect 24398 22370 24454 22379
rect 24398 22305 24454 22314
rect 20956 21214 21252 21234
rect 21012 21212 21036 21214
rect 21092 21212 21116 21214
rect 21172 21212 21196 21214
rect 21034 21160 21036 21212
rect 21098 21160 21110 21212
rect 21172 21160 21174 21212
rect 21012 21158 21036 21160
rect 21092 21158 21116 21160
rect 21172 21158 21196 21160
rect 20956 21138 21252 21158
rect 19432 20770 19484 20776
rect 19432 20712 19484 20718
rect 19616 20770 19668 20776
rect 19616 20712 19668 20718
rect 16762 18970 16818 18979
rect 16762 18905 16764 18914
rect 16816 18905 16818 18914
rect 18694 18970 18750 18979
rect 18694 18905 18750 18914
rect 16764 18876 16816 18882
rect 8852 18866 8904 18872
rect 8852 18808 8904 18814
rect 8576 18798 8628 18804
rect 8576 18740 8628 18746
rect 8588 18328 8616 18740
rect 8864 18396 8892 18808
rect 15660 18798 15712 18804
rect 15660 18740 15712 18746
rect 15384 18730 15436 18736
rect 15384 18672 15436 18678
rect 9956 18594 10008 18600
rect 9956 18536 10008 18542
rect 8852 18390 8904 18396
rect 8852 18332 8904 18338
rect 8576 18322 8628 18328
rect 8576 18264 8628 18270
rect 8588 18163 8616 18264
rect 8574 18154 8630 18163
rect 8574 18089 8630 18098
rect 7012 16214 7064 16220
rect 7012 16156 7064 16162
rect 9968 15987 9996 18536
rect 15396 18192 15424 18672
rect 15384 18186 15436 18192
rect 13082 18154 13138 18163
rect 15382 18154 15384 18163
rect 15436 18154 15438 18163
rect 13082 18089 13138 18098
rect 15200 18118 15252 18124
rect 10956 17950 11252 17970
rect 11012 17948 11036 17950
rect 11092 17948 11116 17950
rect 11172 17948 11196 17950
rect 11034 17896 11036 17948
rect 11098 17896 11110 17948
rect 11172 17896 11174 17948
rect 11012 17894 11036 17896
rect 11092 17894 11116 17896
rect 11172 17894 11196 17896
rect 10956 17874 11252 17894
rect 10956 16862 11252 16882
rect 11012 16860 11036 16862
rect 11092 16860 11116 16862
rect 11172 16860 11196 16862
rect 11034 16808 11036 16860
rect 11098 16808 11110 16860
rect 11172 16808 11174 16860
rect 11012 16806 11036 16808
rect 11092 16806 11116 16808
rect 11172 16806 11196 16808
rect 10956 16786 11252 16806
rect 13096 16628 13124 18089
rect 15672 18124 15700 18740
rect 15956 18494 16252 18514
rect 16012 18492 16036 18494
rect 16092 18492 16116 18494
rect 16172 18492 16196 18494
rect 16034 18440 16036 18492
rect 16098 18440 16110 18492
rect 16172 18440 16174 18492
rect 16012 18438 16036 18440
rect 16092 18438 16116 18440
rect 16172 18438 16196 18440
rect 15956 18418 16252 18438
rect 15382 18089 15438 18098
rect 15660 18118 15712 18124
rect 15200 18060 15252 18066
rect 15396 18063 15424 18089
rect 15660 18060 15712 18066
rect 13542 16930 13598 16939
rect 13542 16865 13598 16874
rect 13084 16622 13136 16628
rect 13084 16564 13136 16570
rect 13096 16220 13124 16564
rect 13084 16214 13136 16220
rect 13084 16156 13136 16162
rect 7194 15978 7250 15987
rect 7194 15913 7196 15922
rect 7248 15913 7250 15922
rect 9954 15978 10010 15987
rect 9954 15913 10010 15922
rect 7196 15884 7248 15890
rect 7208 15676 7236 15884
rect 8484 15874 8536 15880
rect 8484 15816 8536 15822
rect 13452 15874 13504 15880
rect 13452 15816 13504 15822
rect 7196 15670 7248 15676
rect 7196 15612 7248 15618
rect 5956 15230 6252 15250
rect 6012 15228 6036 15230
rect 6092 15228 6116 15230
rect 6172 15228 6196 15230
rect 6034 15176 6036 15228
rect 6098 15176 6110 15228
rect 6172 15176 6174 15228
rect 6012 15174 6036 15176
rect 6092 15174 6116 15176
rect 6172 15174 6196 15176
rect 5956 15154 6252 15174
rect 5956 14142 6252 14162
rect 6012 14140 6036 14142
rect 6092 14140 6116 14142
rect 6172 14140 6196 14142
rect 6034 14088 6036 14140
rect 6098 14088 6110 14140
rect 6172 14088 6174 14140
rect 6012 14086 6036 14088
rect 6092 14086 6116 14088
rect 6172 14086 6196 14088
rect 5956 14066 6252 14086
rect 5956 13054 6252 13074
rect 6012 13052 6036 13054
rect 6092 13052 6116 13054
rect 6172 13052 6196 13054
rect 6034 13000 6036 13052
rect 6098 13000 6110 13052
rect 6172 13000 6174 13052
rect 6012 12998 6036 13000
rect 6092 12998 6116 13000
rect 6172 12998 6196 13000
rect 5956 12978 6252 12998
rect 5956 11966 6252 11986
rect 6012 11964 6036 11966
rect 6092 11964 6116 11966
rect 6172 11964 6196 11966
rect 6034 11912 6036 11964
rect 6098 11912 6110 11964
rect 6172 11912 6174 11964
rect 6012 11910 6036 11912
rect 6092 11910 6116 11912
rect 6172 11910 6196 11912
rect 5956 11890 6252 11910
rect 7102 11354 7158 11363
rect 7102 11289 7158 11298
rect 5956 10878 6252 10898
rect 6012 10876 6036 10878
rect 6092 10876 6116 10878
rect 6172 10876 6196 10878
rect 6034 10824 6036 10876
rect 6098 10824 6110 10876
rect 6172 10824 6174 10876
rect 6012 10822 6036 10824
rect 6092 10822 6116 10824
rect 6172 10822 6196 10824
rect 5956 10802 6252 10822
rect 7116 10780 7144 11289
rect 7208 11188 7236 15612
rect 8496 15171 8524 15816
rect 10956 15774 11252 15794
rect 11012 15772 11036 15774
rect 11092 15772 11116 15774
rect 11172 15772 11196 15774
rect 11034 15720 11036 15772
rect 11098 15720 11110 15772
rect 11172 15720 11174 15772
rect 11012 15718 11036 15720
rect 11092 15718 11116 15720
rect 11172 15718 11196 15720
rect 10956 15698 11252 15718
rect 13464 15171 13492 15816
rect 8482 15162 8538 15171
rect 8482 15097 8538 15106
rect 13450 15162 13506 15171
rect 13450 15097 13506 15106
rect 8300 12406 8352 12412
rect 8300 12348 8352 12354
rect 7378 12170 7434 12179
rect 7378 12105 7434 12114
rect 7930 12170 7986 12179
rect 7930 12105 7932 12114
rect 7196 11182 7248 11188
rect 7196 11124 7248 11130
rect 7392 11120 7420 12105
rect 7984 12105 7986 12114
rect 7932 12076 7984 12082
rect 8114 11762 8170 11771
rect 8114 11697 8170 11706
rect 8128 11363 8156 11697
rect 8312 11528 8340 12348
rect 8496 12208 8524 15097
rect 10956 14686 11252 14706
rect 11012 14684 11036 14686
rect 11092 14684 11116 14686
rect 11172 14684 11196 14686
rect 11034 14632 11036 14684
rect 11098 14632 11110 14684
rect 11172 14632 11174 14684
rect 11012 14630 11036 14632
rect 11092 14630 11116 14632
rect 11172 14630 11196 14632
rect 10956 14610 11252 14630
rect 13464 14491 13492 15097
rect 13450 14482 13506 14491
rect 13450 14417 13506 14426
rect 10956 13598 11252 13618
rect 11012 13596 11036 13598
rect 11092 13596 11116 13598
rect 11172 13596 11196 13598
rect 11034 13544 11036 13596
rect 11098 13544 11110 13596
rect 11172 13544 11174 13596
rect 11012 13542 11036 13544
rect 11092 13542 11116 13544
rect 11172 13542 11196 13544
rect 10956 13522 11252 13542
rect 11978 13258 12034 13267
rect 11978 13193 12034 13202
rect 10956 12510 11252 12530
rect 11012 12508 11036 12510
rect 11092 12508 11116 12510
rect 11172 12508 11196 12510
rect 11034 12456 11036 12508
rect 11098 12456 11110 12508
rect 11172 12456 11174 12508
rect 11012 12454 11036 12456
rect 11092 12454 11116 12456
rect 11172 12454 11196 12456
rect 10956 12434 11252 12454
rect 8668 12270 8720 12276
rect 8668 12212 8720 12218
rect 8484 12202 8536 12208
rect 8484 12144 8536 12150
rect 8496 11868 8524 12144
rect 8484 11862 8536 11868
rect 8484 11804 8536 11810
rect 8680 11528 8708 12212
rect 11992 11868 12020 13193
rect 13084 12270 13136 12276
rect 13084 12212 13136 12218
rect 12072 12066 12124 12072
rect 12072 12008 12124 12014
rect 11980 11862 12032 11868
rect 11980 11804 12032 11810
rect 11992 11664 12020 11804
rect 12084 11732 12112 12008
rect 13096 11907 13124 12212
rect 13464 12140 13492 14417
rect 13556 13500 13584 16865
rect 15212 16764 15240 18060
rect 15956 17406 16252 17426
rect 16012 17404 16036 17406
rect 16092 17404 16116 17406
rect 16172 17404 16196 17406
rect 16034 17352 16036 17404
rect 16098 17352 16110 17404
rect 16172 17352 16174 17404
rect 16012 17350 16036 17352
rect 16092 17350 16116 17352
rect 16172 17350 16196 17352
rect 15956 17330 16252 17350
rect 18708 17172 18736 18905
rect 19340 18050 19392 18056
rect 19260 17998 19340 18004
rect 19260 17992 19392 17998
rect 19260 17976 19380 17992
rect 19260 17308 19288 17976
rect 19248 17302 19300 17308
rect 19248 17244 19300 17250
rect 18696 17166 18748 17172
rect 18696 17108 18748 17114
rect 17500 16962 17552 16968
rect 17498 16930 17500 16939
rect 18328 16962 18380 16968
rect 17552 16930 17554 16939
rect 18328 16904 18380 16910
rect 17498 16865 17554 16874
rect 18340 16764 18368 16904
rect 14096 16758 14148 16764
rect 14096 16700 14148 16706
rect 15200 16758 15252 16764
rect 15200 16700 15252 16706
rect 18328 16758 18380 16764
rect 18328 16700 18380 16706
rect 13636 16622 13688 16628
rect 13636 16564 13688 16570
rect 13648 15880 13676 16564
rect 13636 15874 13688 15880
rect 13636 15816 13688 15822
rect 14108 15035 14136 16700
rect 15956 16318 16252 16338
rect 16012 16316 16036 16318
rect 16092 16316 16116 16318
rect 16172 16316 16196 16318
rect 16034 16264 16036 16316
rect 16098 16264 16110 16316
rect 16172 16264 16174 16316
rect 16012 16262 16036 16264
rect 16092 16262 16116 16264
rect 16172 16262 16196 16264
rect 15956 16242 16252 16262
rect 15956 15230 16252 15250
rect 16012 15228 16036 15230
rect 16092 15228 16116 15230
rect 16172 15228 16196 15230
rect 16034 15176 16036 15228
rect 16098 15176 16110 15228
rect 16172 15176 16174 15228
rect 16012 15174 16036 15176
rect 16092 15174 16116 15176
rect 16172 15174 16196 15176
rect 15956 15154 16252 15174
rect 18340 15132 18368 16700
rect 19248 15330 19300 15336
rect 19248 15272 19300 15278
rect 18328 15126 18380 15132
rect 18328 15068 18380 15074
rect 14094 15026 14150 15035
rect 14094 14961 14150 14970
rect 18786 15026 18842 15035
rect 18786 14961 18788 14970
rect 13544 13494 13596 13500
rect 13544 13436 13596 13442
rect 13820 13358 13872 13364
rect 13820 13300 13872 13306
rect 13832 12684 13860 13300
rect 14108 13296 14136 14961
rect 18840 14961 18842 14970
rect 19260 15012 19288 15272
rect 19260 14984 19380 15012
rect 18788 14932 18840 14938
rect 15956 14142 16252 14162
rect 16012 14140 16036 14142
rect 16092 14140 16116 14142
rect 16172 14140 16196 14142
rect 16034 14088 16036 14140
rect 16098 14088 16110 14140
rect 16172 14088 16174 14140
rect 16012 14086 16036 14088
rect 16092 14086 16116 14088
rect 16172 14086 16196 14088
rect 15956 14066 16252 14086
rect 19260 13500 19288 14984
rect 19352 14928 19380 14984
rect 19340 14922 19392 14928
rect 19340 14864 19392 14870
rect 19444 14876 19472 20712
rect 19444 14848 19564 14876
rect 19432 14786 19484 14792
rect 19432 14728 19484 14734
rect 19444 14588 19472 14728
rect 19536 14588 19564 14848
rect 19432 14582 19484 14588
rect 19432 14524 19484 14530
rect 19524 14582 19576 14588
rect 19524 14524 19576 14530
rect 19536 14044 19564 14524
rect 19524 14038 19576 14044
rect 19524 13980 19576 13986
rect 19536 13539 19564 13980
rect 19522 13530 19578 13539
rect 19248 13494 19300 13500
rect 19522 13465 19578 13474
rect 19248 13436 19300 13442
rect 19524 13358 19576 13364
rect 19524 13300 19576 13306
rect 14096 13290 14148 13296
rect 14096 13232 14148 13238
rect 19156 13290 19208 13296
rect 19156 13232 19208 13238
rect 13912 13222 13964 13228
rect 13912 13164 13964 13170
rect 13820 12678 13872 12684
rect 13820 12620 13872 12626
rect 13832 12564 13860 12620
rect 13924 12616 13952 13164
rect 14108 12956 14136 13232
rect 15956 13054 16252 13074
rect 16012 13052 16036 13054
rect 16092 13052 16116 13054
rect 16172 13052 16196 13054
rect 16034 13000 16036 13052
rect 16098 13000 16110 13052
rect 16172 13000 16174 13052
rect 16012 12998 16036 13000
rect 16092 12998 16116 13000
rect 16172 12998 16196 13000
rect 15956 12978 16252 12998
rect 14096 12950 14148 12956
rect 14096 12892 14148 12898
rect 19168 12752 19196 13232
rect 19536 12820 19564 13300
rect 19628 13296 19656 20712
rect 24030 20466 24086 20475
rect 24030 20401 24086 20410
rect 20956 20126 21252 20146
rect 21012 20124 21036 20126
rect 21092 20124 21116 20126
rect 21172 20124 21196 20126
rect 21034 20072 21036 20124
rect 21098 20072 21110 20124
rect 21172 20072 21174 20124
rect 21012 20070 21036 20072
rect 21092 20070 21116 20072
rect 21172 20070 21196 20072
rect 20956 20050 21252 20070
rect 20810 19242 20866 19251
rect 20810 19177 20866 19186
rect 20824 18940 20852 19177
rect 23480 19138 23532 19144
rect 23480 19080 23532 19086
rect 20956 19038 21252 19058
rect 21012 19036 21036 19038
rect 21092 19036 21116 19038
rect 21172 19036 21196 19038
rect 21034 18984 21036 19036
rect 21098 18984 21110 19036
rect 21172 18984 21174 19036
rect 21012 18982 21036 18984
rect 21092 18982 21116 18984
rect 21172 18982 21196 18984
rect 20956 18962 21252 18982
rect 20812 18934 20864 18940
rect 20812 18876 20864 18882
rect 20628 18798 20680 18804
rect 20628 18740 20680 18746
rect 19890 18426 19946 18435
rect 19890 18361 19946 18370
rect 19904 14384 19932 18361
rect 20640 18056 20668 18740
rect 20628 18050 20680 18056
rect 20628 17992 20680 17998
rect 20956 17950 21252 17970
rect 21012 17948 21036 17950
rect 21092 17948 21116 17950
rect 21172 17948 21196 17950
rect 21034 17896 21036 17948
rect 21098 17896 21110 17948
rect 21172 17896 21174 17948
rect 21012 17894 21036 17896
rect 21092 17894 21116 17896
rect 21172 17894 21196 17896
rect 20956 17874 21252 17894
rect 20956 16862 21252 16882
rect 21012 16860 21036 16862
rect 21092 16860 21116 16862
rect 21172 16860 21196 16862
rect 21034 16808 21036 16860
rect 21098 16808 21110 16860
rect 21172 16808 21174 16860
rect 21012 16806 21036 16808
rect 21092 16806 21116 16808
rect 21172 16806 21196 16808
rect 20956 16786 21252 16806
rect 21454 15842 21510 15851
rect 20956 15774 21252 15794
rect 21454 15777 21510 15786
rect 21012 15772 21036 15774
rect 21092 15772 21116 15774
rect 21172 15772 21196 15774
rect 21034 15720 21036 15772
rect 21098 15720 21110 15772
rect 21172 15720 21174 15772
rect 21012 15718 21036 15720
rect 21092 15718 21116 15720
rect 21172 15718 21196 15720
rect 20956 15698 21252 15718
rect 20956 14686 21252 14706
rect 21012 14684 21036 14686
rect 21092 14684 21116 14686
rect 21172 14684 21196 14686
rect 21034 14632 21036 14684
rect 21098 14632 21110 14684
rect 21172 14632 21174 14684
rect 21012 14630 21036 14632
rect 21092 14630 21116 14632
rect 21172 14630 21196 14632
rect 20956 14610 21252 14630
rect 19982 14482 20038 14491
rect 19982 14417 20038 14426
rect 19996 14384 20024 14417
rect 19708 14378 19760 14384
rect 19708 14320 19760 14326
rect 19892 14378 19944 14384
rect 19892 14320 19944 14326
rect 19984 14378 20036 14384
rect 19984 14320 20036 14326
rect 19720 13840 19748 14320
rect 19996 14044 20024 14320
rect 19984 14038 20036 14044
rect 19984 13980 20036 13986
rect 19708 13834 19760 13840
rect 19708 13776 19760 13782
rect 19720 13403 19748 13776
rect 19706 13394 19762 13403
rect 19706 13329 19762 13338
rect 19996 13296 20024 13980
rect 20956 13598 21252 13618
rect 21012 13596 21036 13598
rect 21092 13596 21116 13598
rect 21172 13596 21196 13598
rect 21034 13544 21036 13596
rect 21098 13544 21110 13596
rect 21172 13544 21174 13596
rect 21012 13542 21036 13544
rect 21092 13542 21116 13544
rect 21172 13542 21196 13544
rect 20956 13522 21252 13542
rect 19616 13290 19668 13296
rect 19616 13232 19668 13238
rect 19984 13290 20036 13296
rect 19984 13232 20036 13238
rect 19996 12956 20024 13232
rect 19984 12950 20036 12956
rect 19984 12892 20036 12898
rect 19524 12814 19576 12820
rect 19524 12756 19576 12762
rect 19156 12746 19208 12752
rect 19154 12714 19156 12723
rect 19208 12714 19210 12723
rect 19154 12649 19210 12658
rect 13740 12536 13860 12564
rect 13912 12610 13964 12616
rect 13912 12552 13964 12558
rect 13740 12412 13768 12536
rect 13728 12406 13780 12412
rect 13728 12348 13780 12354
rect 13544 12202 13596 12208
rect 13924 12179 13952 12552
rect 20956 12510 21252 12530
rect 21012 12508 21036 12510
rect 21092 12508 21116 12510
rect 21172 12508 21196 12510
rect 21034 12456 21036 12508
rect 21098 12456 21110 12508
rect 21172 12456 21174 12508
rect 21012 12454 21036 12456
rect 21092 12454 21116 12456
rect 21172 12454 21196 12456
rect 20956 12434 21252 12454
rect 13544 12144 13596 12150
rect 13910 12170 13966 12179
rect 13452 12134 13504 12140
rect 13452 12076 13504 12082
rect 13082 11898 13138 11907
rect 13082 11833 13138 11842
rect 13096 11800 13124 11833
rect 13084 11794 13136 11800
rect 13084 11736 13136 11742
rect 13464 11732 13492 12076
rect 13556 11868 13584 12144
rect 13910 12105 13966 12114
rect 15956 11966 16252 11986
rect 16012 11964 16036 11966
rect 16092 11964 16116 11966
rect 16172 11964 16196 11966
rect 16034 11912 16036 11964
rect 16098 11912 16110 11964
rect 16172 11912 16174 11964
rect 16012 11910 16036 11912
rect 16092 11910 16116 11912
rect 16172 11910 16196 11912
rect 14738 11898 14794 11907
rect 13544 11862 13596 11868
rect 15956 11890 16252 11910
rect 14738 11833 14794 11842
rect 13544 11804 13596 11810
rect 12072 11726 12124 11732
rect 12072 11668 12124 11674
rect 13452 11726 13504 11732
rect 13452 11668 13504 11674
rect 11980 11658 12032 11664
rect 11980 11600 12032 11606
rect 8300 11522 8352 11528
rect 8300 11464 8352 11470
rect 8668 11522 8720 11528
rect 8668 11464 8720 11470
rect 8114 11354 8170 11363
rect 8312 11340 8340 11464
rect 8114 11289 8170 11298
rect 8220 11312 8340 11340
rect 8680 11324 8708 11464
rect 10956 11422 11252 11442
rect 11012 11420 11036 11422
rect 11092 11420 11116 11422
rect 11172 11420 11196 11422
rect 11034 11368 11036 11420
rect 11098 11368 11110 11420
rect 11172 11368 11174 11420
rect 11012 11366 11036 11368
rect 11092 11366 11116 11368
rect 11172 11366 11196 11368
rect 10956 11346 11252 11366
rect 8668 11318 8720 11324
rect 8128 11256 8156 11289
rect 8116 11250 8168 11256
rect 8116 11192 8168 11198
rect 7380 11114 7432 11120
rect 7380 11056 7432 11062
rect 7104 10774 7156 10780
rect 7104 10716 7156 10722
rect 7392 10440 7420 11056
rect 8220 10780 8248 11312
rect 8668 11260 8720 11266
rect 8300 11114 8352 11120
rect 8298 11082 8300 11091
rect 12084 11091 12112 11668
rect 12624 11658 12676 11664
rect 12162 11626 12218 11635
rect 12624 11600 12676 11606
rect 12162 11561 12218 11570
rect 12176 11528 12204 11561
rect 12164 11522 12216 11528
rect 12164 11464 12216 11470
rect 12176 11324 12204 11464
rect 12164 11318 12216 11324
rect 12164 11260 12216 11266
rect 8352 11082 8354 11091
rect 8298 11017 8354 11026
rect 12070 11082 12126 11091
rect 12070 11017 12126 11026
rect 8312 10780 8340 11017
rect 8208 10774 8260 10780
rect 8208 10716 8260 10722
rect 8300 10774 8352 10780
rect 8300 10716 8352 10722
rect 8576 10638 8628 10644
rect 8576 10580 8628 10586
rect 8298 10538 8354 10547
rect 8298 10473 8300 10482
rect 8352 10473 8354 10482
rect 8300 10444 8352 10450
rect 7380 10434 7432 10440
rect 7380 10376 7432 10382
rect 7840 10434 7892 10440
rect 7840 10376 7892 10382
rect 5956 9790 6252 9810
rect 6012 9788 6036 9790
rect 6092 9788 6116 9790
rect 6172 9788 6196 9790
rect 6034 9736 6036 9788
rect 6098 9736 6110 9788
rect 6172 9736 6174 9788
rect 6012 9734 6036 9736
rect 6092 9734 6116 9736
rect 6172 9734 6196 9736
rect 5956 9714 6252 9734
rect 4158 9586 4214 9595
rect 4158 9521 4214 9530
rect 3896 7640 4108 7668
rect 3790 7410 3846 7419
rect 3790 7345 3846 7354
rect 3606 7274 3662 7283
rect 3606 7209 3662 7218
rect 3514 5234 3570 5243
rect 3514 5169 3570 5178
rect 3896 4699 3924 7640
rect 4172 5748 4200 9521
rect 5956 8702 6252 8722
rect 6012 8700 6036 8702
rect 6092 8700 6116 8702
rect 6172 8700 6196 8702
rect 6034 8648 6036 8700
rect 6098 8648 6110 8700
rect 6172 8648 6174 8700
rect 6012 8646 6036 8648
rect 6092 8646 6116 8648
rect 6172 8646 6196 8648
rect 5956 8626 6252 8646
rect 5956 7614 6252 7634
rect 6012 7612 6036 7614
rect 6092 7612 6116 7614
rect 6172 7612 6196 7614
rect 6034 7560 6036 7612
rect 6098 7560 6110 7612
rect 6172 7560 6174 7612
rect 6012 7558 6036 7560
rect 6092 7558 6116 7560
rect 6172 7558 6196 7560
rect 5956 7538 6252 7558
rect 5956 6526 6252 6546
rect 6012 6524 6036 6526
rect 6092 6524 6116 6526
rect 6172 6524 6196 6526
rect 6034 6472 6036 6524
rect 6098 6472 6110 6524
rect 6172 6472 6174 6524
rect 6012 6470 6036 6472
rect 6092 6470 6116 6472
rect 6172 6470 6196 6472
rect 5956 6450 6252 6470
rect 4160 5742 4212 5748
rect 4160 5684 4212 5690
rect 4172 5340 4200 5684
rect 4342 5642 4398 5651
rect 4342 5577 4344 5586
rect 4396 5577 4398 5586
rect 4344 5548 4396 5554
rect 5956 5438 6252 5458
rect 6012 5436 6036 5438
rect 6092 5436 6116 5438
rect 6172 5436 6196 5438
rect 6034 5384 6036 5436
rect 6098 5384 6110 5436
rect 6172 5384 6174 5436
rect 6012 5382 6036 5384
rect 6092 5382 6116 5384
rect 6172 5382 6196 5384
rect 5956 5362 6252 5382
rect 4160 5334 4212 5340
rect 4160 5276 4212 5282
rect 3882 4690 3938 4699
rect 3882 4625 3938 4634
rect 5956 4350 6252 4370
rect 6012 4348 6036 4350
rect 6092 4348 6116 4350
rect 6172 4348 6196 4350
rect 6034 4296 6036 4348
rect 6098 4296 6110 4348
rect 6172 4296 6174 4348
rect 6012 4294 6036 4296
rect 6092 4294 6116 4296
rect 6172 4294 6196 4296
rect 5956 4274 6252 4294
rect 3422 4010 3478 4019
rect 3422 3945 3478 3954
rect 5956 3262 6252 3282
rect 6012 3260 6036 3262
rect 6092 3260 6116 3262
rect 6172 3260 6196 3262
rect 6034 3208 6036 3260
rect 6098 3208 6110 3260
rect 6172 3208 6174 3260
rect 6012 3206 6036 3208
rect 6092 3206 6116 3208
rect 6172 3206 6196 3208
rect 5956 3186 6252 3206
rect 7392 3067 7420 10376
rect 7852 10275 7880 10376
rect 7838 10266 7894 10275
rect 8312 10236 8340 10444
rect 8392 10434 8444 10440
rect 8392 10376 8444 10382
rect 7838 10201 7894 10210
rect 8300 10230 8352 10236
rect 8300 10172 8352 10178
rect 8312 10003 8340 10172
rect 8298 9994 8354 10003
rect 8298 9929 8354 9938
rect 7378 3058 7434 3067
rect 7378 2993 7434 3002
rect 8404 2523 8432 10376
rect 8588 10236 8616 10580
rect 10956 10334 11252 10354
rect 11012 10332 11036 10334
rect 11092 10332 11116 10334
rect 11172 10332 11196 10334
rect 11034 10280 11036 10332
rect 11098 10280 11110 10332
rect 11172 10280 11174 10332
rect 11012 10278 11036 10280
rect 11092 10278 11116 10280
rect 11172 10278 11196 10280
rect 10956 10258 11252 10278
rect 8576 10230 8628 10236
rect 8576 10172 8628 10178
rect 10956 9246 11252 9266
rect 11012 9244 11036 9246
rect 11092 9244 11116 9246
rect 11172 9244 11196 9246
rect 11034 9192 11036 9244
rect 11098 9192 11110 9244
rect 11172 9192 11174 9244
rect 11012 9190 11036 9192
rect 11092 9190 11116 9192
rect 11172 9190 11196 9192
rect 10956 9170 11252 9190
rect 10956 8158 11252 8178
rect 11012 8156 11036 8158
rect 11092 8156 11116 8158
rect 11172 8156 11196 8158
rect 11034 8104 11036 8156
rect 11098 8104 11110 8156
rect 11172 8104 11174 8156
rect 11012 8102 11036 8104
rect 11092 8102 11116 8104
rect 11172 8102 11196 8104
rect 10956 8082 11252 8102
rect 10956 7070 11252 7090
rect 11012 7068 11036 7070
rect 11092 7068 11116 7070
rect 11172 7068 11196 7070
rect 11034 7016 11036 7068
rect 11098 7016 11110 7068
rect 11172 7016 11174 7068
rect 11012 7014 11036 7016
rect 11092 7014 11116 7016
rect 11172 7014 11196 7016
rect 10956 6994 11252 7014
rect 12636 6852 12664 11600
rect 13082 7818 13138 7827
rect 13082 7753 13138 7762
rect 13096 7312 13124 7753
rect 13084 7306 13136 7312
rect 13084 7248 13136 7254
rect 13268 7170 13320 7176
rect 13266 7138 13268 7147
rect 13320 7138 13322 7147
rect 13266 7073 13322 7082
rect 12636 6824 12756 6852
rect 14752 6836 14780 11833
rect 20956 11422 21252 11442
rect 21012 11420 21036 11422
rect 21092 11420 21116 11422
rect 21172 11420 21196 11422
rect 21034 11368 21036 11420
rect 21098 11368 21110 11420
rect 21172 11368 21174 11420
rect 21012 11366 21036 11368
rect 21092 11366 21116 11368
rect 21172 11366 21196 11368
rect 20956 11346 21252 11366
rect 15956 10878 16252 10898
rect 16012 10876 16036 10878
rect 16092 10876 16116 10878
rect 16172 10876 16196 10878
rect 16034 10824 16036 10876
rect 16098 10824 16110 10876
rect 16172 10824 16174 10876
rect 16012 10822 16036 10824
rect 16092 10822 16116 10824
rect 16172 10822 16196 10824
rect 15956 10802 16252 10822
rect 20956 10334 21252 10354
rect 21012 10332 21036 10334
rect 21092 10332 21116 10334
rect 21172 10332 21196 10334
rect 21034 10280 21036 10332
rect 21098 10280 21110 10332
rect 21172 10280 21174 10332
rect 21012 10278 21036 10280
rect 21092 10278 21116 10280
rect 21172 10278 21196 10280
rect 20956 10258 21252 10278
rect 15956 9790 16252 9810
rect 16012 9788 16036 9790
rect 16092 9788 16116 9790
rect 16172 9788 16196 9790
rect 16034 9736 16036 9788
rect 16098 9736 16110 9788
rect 16172 9736 16174 9788
rect 16012 9734 16036 9736
rect 16092 9734 16116 9736
rect 16172 9734 16196 9736
rect 15956 9714 16252 9734
rect 20956 9246 21252 9266
rect 21012 9244 21036 9246
rect 21092 9244 21116 9246
rect 21172 9244 21196 9246
rect 21034 9192 21036 9244
rect 21098 9192 21110 9244
rect 21172 9192 21174 9244
rect 21012 9190 21036 9192
rect 21092 9190 21116 9192
rect 21172 9190 21196 9192
rect 20956 9170 21252 9190
rect 15956 8702 16252 8722
rect 16012 8700 16036 8702
rect 16092 8700 16116 8702
rect 16172 8700 16196 8702
rect 16034 8648 16036 8700
rect 16098 8648 16110 8700
rect 16172 8648 16174 8700
rect 16012 8646 16036 8648
rect 16092 8646 16116 8648
rect 16172 8646 16196 8648
rect 15956 8626 16252 8646
rect 20956 8158 21252 8178
rect 21012 8156 21036 8158
rect 21092 8156 21116 8158
rect 21172 8156 21196 8158
rect 21034 8104 21036 8156
rect 21098 8104 21110 8156
rect 21172 8104 21174 8156
rect 21012 8102 21036 8104
rect 21092 8102 21116 8104
rect 21172 8102 21196 8104
rect 20956 8082 21252 8102
rect 15956 7614 16252 7634
rect 16012 7612 16036 7614
rect 16092 7612 16116 7614
rect 16172 7612 16196 7614
rect 16034 7560 16036 7612
rect 16098 7560 16110 7612
rect 16172 7560 16174 7612
rect 16012 7558 16036 7560
rect 16092 7558 16116 7560
rect 16172 7558 16196 7560
rect 15956 7538 16252 7558
rect 20534 7546 20590 7555
rect 20534 7481 20590 7490
rect 18604 7442 18656 7448
rect 18418 7410 18474 7419
rect 18418 7345 18474 7354
rect 18602 7410 18604 7419
rect 18656 7410 18658 7419
rect 18602 7345 18658 7354
rect 18432 7312 18460 7345
rect 18420 7306 18472 7312
rect 20548 7283 20576 7481
rect 18420 7248 18472 7254
rect 20534 7274 20590 7283
rect 20534 7209 20590 7218
rect 20956 7070 21252 7090
rect 21012 7068 21036 7070
rect 21092 7068 21116 7070
rect 21172 7068 21196 7070
rect 21034 7016 21036 7068
rect 21098 7016 21110 7068
rect 21172 7016 21174 7068
rect 21012 7014 21036 7016
rect 21092 7014 21116 7016
rect 21172 7014 21196 7016
rect 20956 6994 21252 7014
rect 14922 6866 14978 6875
rect 10956 5982 11252 6002
rect 11012 5980 11036 5982
rect 11092 5980 11116 5982
rect 11172 5980 11196 5982
rect 11034 5928 11036 5980
rect 11098 5928 11110 5980
rect 11172 5928 11174 5980
rect 11012 5926 11036 5928
rect 11092 5926 11116 5928
rect 11172 5926 11196 5928
rect 10956 5906 11252 5926
rect 12622 5234 12678 5243
rect 12622 5169 12678 5178
rect 12636 5136 12664 5169
rect 12624 5130 12676 5136
rect 12624 5072 12676 5078
rect 10956 4894 11252 4914
rect 11012 4892 11036 4894
rect 11092 4892 11116 4894
rect 11172 4892 11196 4894
rect 11034 4840 11036 4892
rect 11098 4840 11110 4892
rect 11172 4840 11174 4892
rect 11012 4838 11036 4840
rect 11092 4838 11116 4840
rect 11172 4838 11196 4840
rect 10956 4818 11252 4838
rect 10956 3806 11252 3826
rect 11012 3804 11036 3806
rect 11092 3804 11116 3806
rect 11172 3804 11196 3806
rect 11034 3752 11036 3804
rect 11098 3752 11110 3804
rect 11172 3752 11174 3804
rect 11012 3750 11036 3752
rect 11092 3750 11116 3752
rect 11172 3750 11196 3752
rect 10956 3730 11252 3750
rect 9496 2818 9548 2824
rect 9496 2760 9548 2766
rect 8390 2514 8446 2523
rect 8390 2449 8446 2458
rect 5956 2174 6252 2194
rect 6012 2172 6036 2174
rect 6092 2172 6116 2174
rect 6172 2172 6196 2174
rect 6034 2120 6036 2172
rect 6098 2120 6110 2172
rect 6172 2120 6174 2172
rect 6012 2118 6036 2120
rect 6092 2118 6116 2120
rect 6172 2118 6196 2120
rect 5956 2098 6252 2118
rect 2134 1426 2190 1435
rect 2134 1361 2190 1370
rect 1582 882 1638 891
rect 1582 817 1638 826
rect 1398 338 1454 347
rect 1398 273 1454 282
rect 9508 75 9536 2760
rect 10956 2718 11252 2738
rect 11012 2716 11036 2718
rect 11092 2716 11116 2718
rect 11172 2716 11196 2718
rect 11034 2664 11036 2716
rect 11098 2664 11110 2716
rect 11172 2664 11174 2716
rect 11012 2662 11036 2664
rect 11092 2662 11116 2664
rect 11172 2662 11196 2664
rect 10956 2642 11252 2662
rect 12728 1979 12756 6824
rect 14740 6830 14792 6836
rect 14922 6801 14978 6810
rect 14740 6772 14792 6778
rect 14752 6428 14780 6772
rect 14936 6700 14964 6801
rect 14924 6694 14976 6700
rect 14924 6636 14976 6642
rect 15956 6526 16252 6546
rect 16012 6524 16036 6526
rect 16092 6524 16116 6526
rect 16172 6524 16196 6526
rect 16034 6472 16036 6524
rect 16098 6472 16110 6524
rect 16172 6472 16174 6524
rect 16012 6470 16036 6472
rect 16092 6470 16116 6472
rect 16172 6470 16196 6472
rect 15956 6450 16252 6470
rect 14740 6422 14792 6428
rect 14740 6364 14792 6370
rect 20956 5982 21252 6002
rect 21012 5980 21036 5982
rect 21092 5980 21116 5982
rect 21172 5980 21196 5982
rect 21034 5928 21036 5980
rect 21098 5928 21110 5980
rect 21172 5928 21174 5980
rect 21012 5926 21036 5928
rect 21092 5926 21116 5928
rect 21172 5926 21196 5928
rect 20956 5906 21252 5926
rect 13084 5878 13136 5884
rect 13084 5820 13136 5826
rect 13096 5787 13124 5820
rect 13082 5778 13138 5787
rect 13082 5713 13138 5722
rect 13634 5778 13690 5787
rect 13634 5713 13636 5722
rect 13688 5713 13690 5722
rect 13636 5684 13688 5690
rect 13648 5340 13676 5684
rect 15956 5438 16252 5458
rect 16012 5436 16036 5438
rect 16092 5436 16116 5438
rect 16172 5436 16196 5438
rect 16034 5384 16036 5436
rect 16098 5384 16110 5436
rect 16172 5384 16174 5436
rect 16012 5382 16036 5384
rect 16092 5382 16116 5384
rect 16172 5382 16196 5384
rect 15956 5362 16252 5382
rect 13636 5334 13688 5340
rect 13636 5276 13688 5282
rect 15566 5234 15622 5243
rect 15566 5169 15622 5178
rect 12808 4994 12860 5000
rect 12808 4936 12860 4942
rect 12820 4155 12848 4936
rect 15580 4660 15608 5169
rect 20956 4894 21252 4914
rect 21012 4892 21036 4894
rect 21092 4892 21116 4894
rect 21172 4892 21196 4894
rect 21034 4840 21036 4892
rect 21098 4840 21110 4892
rect 21172 4840 21174 4892
rect 21012 4838 21036 4840
rect 21092 4838 21116 4840
rect 21172 4838 21196 4840
rect 20956 4818 21252 4838
rect 20442 4690 20498 4699
rect 15568 4654 15620 4660
rect 20442 4625 20444 4634
rect 15568 4596 15620 4602
rect 20496 4625 20498 4634
rect 20444 4596 20496 4602
rect 15580 4252 15608 4596
rect 15750 4554 15806 4563
rect 15750 4489 15752 4498
rect 15804 4489 15806 4498
rect 15752 4460 15804 4466
rect 15956 4350 16252 4370
rect 16012 4348 16036 4350
rect 16092 4348 16116 4350
rect 16172 4348 16196 4350
rect 16034 4296 16036 4348
rect 16098 4296 16110 4348
rect 16172 4296 16174 4348
rect 16012 4294 16036 4296
rect 16092 4294 16116 4296
rect 16172 4294 16196 4296
rect 15956 4274 16252 4294
rect 20456 4252 20484 4596
rect 20626 4554 20682 4563
rect 20626 4489 20628 4498
rect 20680 4489 20682 4498
rect 20628 4460 20680 4466
rect 15568 4246 15620 4252
rect 15568 4188 15620 4194
rect 20444 4246 20496 4252
rect 20444 4188 20496 4194
rect 12806 4146 12862 4155
rect 21468 4116 21496 15777
rect 22926 13802 22982 13811
rect 22926 13737 22982 13746
rect 22466 7682 22522 7691
rect 22466 7617 22522 7626
rect 22480 7516 22508 7617
rect 22940 7516 22968 13737
rect 23492 12315 23520 19080
rect 23938 18834 23994 18843
rect 23938 18769 23940 18778
rect 23992 18769 23994 18778
rect 23940 18740 23992 18746
rect 23952 18396 23980 18740
rect 23940 18390 23992 18396
rect 23940 18332 23992 18338
rect 23938 18290 23994 18299
rect 23938 18225 23994 18234
rect 23952 18192 23980 18225
rect 23940 18186 23992 18192
rect 23940 18128 23992 18134
rect 23754 17882 23810 17891
rect 23754 17817 23810 17826
rect 23664 15874 23716 15880
rect 23664 15816 23716 15822
rect 23572 14242 23624 14248
rect 23572 14184 23624 14190
rect 23478 12306 23534 12315
rect 23478 12241 23534 12250
rect 23480 8530 23532 8536
rect 23480 8472 23532 8478
rect 23492 7963 23520 8472
rect 23584 8371 23612 14184
rect 23676 9459 23704 15816
rect 23662 9450 23718 9459
rect 23662 9385 23718 9394
rect 23768 8604 23796 17817
rect 23938 17746 23994 17755
rect 23938 17681 23940 17690
rect 23992 17681 23994 17690
rect 23940 17652 23992 17658
rect 23952 17308 23980 17652
rect 23940 17302 23992 17308
rect 23940 17244 23992 17250
rect 24044 14452 24072 20401
rect 24124 18594 24176 18600
rect 24124 18536 24176 18542
rect 24032 14446 24084 14452
rect 24032 14388 24084 14394
rect 24044 14044 24072 14388
rect 24032 14038 24084 14044
rect 24032 13980 24084 13986
rect 23938 13394 23994 13403
rect 23938 13329 23994 13338
rect 23952 11188 23980 13329
rect 24030 12442 24086 12451
rect 24030 12377 24086 12386
rect 23940 11182 23992 11188
rect 23940 11124 23992 11130
rect 23952 10780 23980 11124
rect 23940 10774 23992 10780
rect 23940 10716 23992 10722
rect 23938 9586 23994 9595
rect 23938 9521 23994 9530
rect 23952 9488 23980 9521
rect 23940 9482 23992 9488
rect 23940 9424 23992 9430
rect 23938 9042 23994 9051
rect 23938 8977 23940 8986
rect 23992 8977 23994 8986
rect 23940 8948 23992 8954
rect 23952 8604 23980 8948
rect 23756 8598 23808 8604
rect 23756 8540 23808 8546
rect 23940 8598 23992 8604
rect 23940 8540 23992 8546
rect 23768 8400 23796 8540
rect 23756 8394 23808 8400
rect 23570 8362 23626 8371
rect 23756 8336 23808 8342
rect 23570 8297 23626 8306
rect 23478 7954 23534 7963
rect 23478 7889 23534 7898
rect 23940 7918 23992 7924
rect 23940 7860 23992 7866
rect 23952 7555 23980 7860
rect 23938 7546 23994 7555
rect 22468 7510 22520 7516
rect 22468 7452 22520 7458
rect 22928 7510 22980 7516
rect 23938 7481 23940 7490
rect 22928 7452 22980 7458
rect 23992 7481 23994 7490
rect 23940 7452 23992 7458
rect 22940 7312 22968 7452
rect 22928 7306 22980 7312
rect 22928 7248 22980 7254
rect 24044 6836 24072 12377
rect 24136 11635 24164 18536
rect 24308 18050 24360 18056
rect 24308 17992 24360 17998
rect 24216 17506 24268 17512
rect 24216 17448 24268 17454
rect 24122 11626 24178 11635
rect 24122 11561 24178 11570
rect 24124 11522 24176 11528
rect 24124 11464 24176 11470
rect 24136 10683 24164 11464
rect 24122 10674 24178 10683
rect 24122 10609 24178 10618
rect 24228 10411 24256 17448
rect 24320 11091 24348 17992
rect 24412 11868 24440 22305
rect 24490 21282 24546 21291
rect 24490 21217 24546 21226
rect 24504 16220 24532 21217
rect 24780 19280 24808 23529
rect 26146 23490 26202 23970
rect 25042 23050 25098 23059
rect 25042 22985 25098 22994
rect 24858 21554 24914 21563
rect 24858 21489 24914 21498
rect 24872 20776 24900 21489
rect 24860 20770 24912 20776
rect 24860 20712 24912 20718
rect 24858 20058 24914 20067
rect 24858 19993 24914 20002
rect 24768 19274 24820 19280
rect 24768 19216 24820 19222
rect 24872 17891 24900 19993
rect 24950 18834 25006 18843
rect 25056 18804 25084 22985
rect 26160 21948 26188 23490
rect 25884 21920 26188 21948
rect 25502 19378 25558 19387
rect 25502 19313 25558 19322
rect 24950 18769 25006 18778
rect 25044 18798 25096 18804
rect 24858 17882 24914 17891
rect 24858 17817 24914 17826
rect 24766 17066 24822 17075
rect 24766 17001 24822 17010
rect 24492 16214 24544 16220
rect 24492 16156 24544 16162
rect 24504 16016 24532 16156
rect 24492 16010 24544 16016
rect 24492 15952 24544 15958
rect 24674 15434 24730 15443
rect 24674 15369 24730 15378
rect 24400 11862 24452 11868
rect 24400 11804 24452 11810
rect 24412 11664 24440 11804
rect 24400 11658 24452 11664
rect 24400 11600 24452 11606
rect 24306 11082 24362 11091
rect 24306 11017 24362 11026
rect 24214 10402 24270 10411
rect 24214 10337 24270 10346
rect 24124 9346 24176 9352
rect 24122 9314 24124 9323
rect 24176 9314 24178 9323
rect 24122 9249 24178 9258
rect 24124 8802 24176 8808
rect 24124 8744 24176 8750
rect 24136 8507 24164 8744
rect 24122 8498 24178 8507
rect 24122 8433 24178 8442
rect 24122 8090 24178 8099
rect 24122 8025 24124 8034
rect 24176 8025 24178 8034
rect 24124 7996 24176 8002
rect 24032 6830 24084 6836
rect 24032 6772 24084 6778
rect 24044 6428 24072 6772
rect 24122 6730 24178 6739
rect 24122 6665 24124 6674
rect 24176 6665 24178 6674
rect 24124 6636 24176 6642
rect 24032 6422 24084 6428
rect 24032 6364 24084 6370
rect 24122 5098 24178 5107
rect 24122 5033 24178 5042
rect 24306 5098 24362 5107
rect 24306 5033 24362 5042
rect 24136 5000 24164 5033
rect 24124 4994 24176 5000
rect 24124 4936 24176 4942
rect 24320 4155 24348 5033
rect 24306 4146 24362 4155
rect 12806 4081 12862 4090
rect 21456 4110 21508 4116
rect 24306 4081 24362 4090
rect 21456 4052 21508 4058
rect 23940 4042 23992 4048
rect 23938 4010 23940 4019
rect 23992 4010 23994 4019
rect 23938 3945 23994 3954
rect 20720 3906 20772 3912
rect 24124 3906 24176 3912
rect 20720 3848 20772 3854
rect 24122 3874 24124 3883
rect 24176 3874 24178 3883
rect 20732 3611 20760 3848
rect 20956 3806 21252 3826
rect 24122 3809 24178 3818
rect 21012 3804 21036 3806
rect 21092 3804 21116 3806
rect 21172 3804 21196 3806
rect 21034 3752 21036 3804
rect 21098 3752 21110 3804
rect 21172 3752 21174 3804
rect 21012 3750 21036 3752
rect 21092 3750 21116 3752
rect 21172 3750 21196 3752
rect 20956 3730 21252 3750
rect 20718 3602 20774 3611
rect 24688 3572 24716 15369
rect 24780 5340 24808 17001
rect 24858 13394 24914 13403
rect 24858 13329 24914 13338
rect 24872 11907 24900 13329
rect 24964 12451 24992 18769
rect 25044 18740 25096 18746
rect 25056 18396 25084 18740
rect 25228 18594 25280 18600
rect 25228 18536 25280 18542
rect 25044 18390 25096 18396
rect 25044 18332 25096 18338
rect 25240 18027 25268 18536
rect 25226 18018 25282 18027
rect 25226 17953 25282 17962
rect 25134 14618 25190 14627
rect 25134 14553 25190 14562
rect 25042 13938 25098 13947
rect 25042 13873 25098 13882
rect 24950 12442 25006 12451
rect 24950 12377 25006 12386
rect 24950 12306 25006 12315
rect 24950 12241 25006 12250
rect 24858 11898 24914 11907
rect 24858 11833 24914 11842
rect 24860 11046 24912 11052
rect 24860 10988 24912 10994
rect 24872 10003 24900 10988
rect 24964 10547 24992 12241
rect 25056 11227 25084 13873
rect 25148 11771 25176 14553
rect 25516 13811 25544 19313
rect 25884 19251 25912 21920
rect 25956 21758 26252 21778
rect 26012 21756 26036 21758
rect 26092 21756 26116 21758
rect 26172 21756 26196 21758
rect 26034 21704 26036 21756
rect 26098 21704 26110 21756
rect 26172 21704 26174 21756
rect 26012 21702 26036 21704
rect 26092 21702 26116 21704
rect 26172 21702 26196 21704
rect 25956 21682 26252 21702
rect 25956 20670 26252 20690
rect 26012 20668 26036 20670
rect 26092 20668 26116 20670
rect 26172 20668 26196 20670
rect 26034 20616 26036 20668
rect 26098 20616 26110 20668
rect 26172 20616 26174 20668
rect 26012 20614 26036 20616
rect 26092 20614 26116 20616
rect 26172 20614 26196 20616
rect 25956 20594 26252 20614
rect 25956 19582 26252 19602
rect 26012 19580 26036 19582
rect 26092 19580 26116 19582
rect 26172 19580 26196 19582
rect 26034 19528 26036 19580
rect 26098 19528 26110 19580
rect 26172 19528 26174 19580
rect 26012 19526 26036 19528
rect 26092 19526 26116 19528
rect 26172 19526 26196 19528
rect 25956 19506 26252 19526
rect 25870 19242 25926 19251
rect 25870 19177 25926 19186
rect 25956 18494 26252 18514
rect 26012 18492 26036 18494
rect 26092 18492 26116 18494
rect 26172 18492 26196 18494
rect 26034 18440 26036 18492
rect 26098 18440 26110 18492
rect 26172 18440 26174 18492
rect 26012 18438 26036 18440
rect 26092 18438 26116 18440
rect 26172 18438 26196 18440
rect 25956 18418 26252 18438
rect 25594 17610 25650 17619
rect 25594 17545 25650 17554
rect 25502 13802 25558 13811
rect 25502 13737 25558 13746
rect 25502 12850 25558 12859
rect 25502 12785 25558 12794
rect 25134 11762 25190 11771
rect 25134 11697 25190 11706
rect 25042 11218 25098 11227
rect 25042 11153 25098 11162
rect 24950 10538 25006 10547
rect 24950 10473 25006 10482
rect 24858 9994 24914 10003
rect 24858 9929 24914 9938
rect 24768 5334 24820 5340
rect 24768 5276 24820 5282
rect 20718 3537 20774 3546
rect 23848 3566 23900 3572
rect 23848 3508 23900 3514
rect 24676 3566 24728 3572
rect 24676 3508 24728 3514
rect 15956 3262 16252 3282
rect 16012 3260 16036 3262
rect 16092 3260 16116 3262
rect 16172 3260 16196 3262
rect 16034 3208 16036 3260
rect 16098 3208 16110 3260
rect 16172 3208 16174 3260
rect 16012 3206 16036 3208
rect 16092 3206 16116 3208
rect 16172 3206 16196 3208
rect 15956 3186 16252 3206
rect 23860 3164 23888 3508
rect 24122 3466 24178 3475
rect 24122 3401 24124 3410
rect 24176 3401 24178 3410
rect 24124 3372 24176 3378
rect 23848 3158 23900 3164
rect 23848 3100 23900 3106
rect 23938 3058 23994 3067
rect 23938 2993 23994 3002
rect 23952 2960 23980 2993
rect 23940 2954 23992 2960
rect 23940 2896 23992 2902
rect 24860 2818 24912 2824
rect 24860 2760 24912 2766
rect 20956 2718 21252 2738
rect 21012 2716 21036 2718
rect 21092 2716 21116 2718
rect 21172 2716 21196 2718
rect 21034 2664 21036 2716
rect 21098 2664 21110 2716
rect 21172 2664 21174 2716
rect 21012 2662 21036 2664
rect 21092 2662 21116 2664
rect 21172 2662 21196 2664
rect 20956 2642 21252 2662
rect 24214 2650 24270 2659
rect 24214 2585 24216 2594
rect 24268 2585 24270 2594
rect 24216 2556 24268 2562
rect 24032 2478 24084 2484
rect 24032 2420 24084 2426
rect 15956 2174 16252 2194
rect 16012 2172 16036 2174
rect 16092 2172 16116 2174
rect 16172 2172 16196 2174
rect 16034 2120 16036 2172
rect 16098 2120 16110 2172
rect 16172 2120 16174 2172
rect 16012 2118 16036 2120
rect 16092 2118 16116 2120
rect 16172 2118 16196 2120
rect 15956 2098 16252 2118
rect 24044 1979 24072 2420
rect 12714 1970 12770 1979
rect 12714 1905 12770 1914
rect 24030 1970 24086 1979
rect 24030 1905 24086 1914
rect 12346 1698 12402 1707
rect 12530 1698 12586 1707
rect 12402 1656 12530 1684
rect 12346 1633 12402 1642
rect 12530 1633 12586 1642
rect 24872 1571 24900 2760
rect 25134 2514 25190 2523
rect 25134 2449 25136 2458
rect 25188 2449 25190 2458
rect 25136 2420 25188 2426
rect 25516 2387 25544 12785
rect 25608 5787 25636 17545
rect 25956 17406 26252 17426
rect 26012 17404 26036 17406
rect 26092 17404 26116 17406
rect 26172 17404 26196 17406
rect 26034 17352 26036 17404
rect 26098 17352 26110 17404
rect 26172 17352 26174 17404
rect 26012 17350 26036 17352
rect 26092 17350 26116 17352
rect 26172 17350 26196 17352
rect 25956 17330 26252 17350
rect 25956 16318 26252 16338
rect 26012 16316 26036 16318
rect 26092 16316 26116 16318
rect 26172 16316 26196 16318
rect 26034 16264 26036 16316
rect 26098 16264 26110 16316
rect 26172 16264 26174 16316
rect 26012 16262 26036 16264
rect 26092 16262 26116 16264
rect 26172 16262 26196 16264
rect 25956 16242 26252 16262
rect 25686 16114 25742 16123
rect 25686 16049 25742 16058
rect 25594 5778 25650 5787
rect 25594 5713 25650 5722
rect 25700 5243 25728 16049
rect 25956 15230 26252 15250
rect 26012 15228 26036 15230
rect 26092 15228 26116 15230
rect 26172 15228 26196 15230
rect 26034 15176 26036 15228
rect 26098 15176 26110 15228
rect 26172 15176 26174 15228
rect 26012 15174 26036 15176
rect 26092 15174 26116 15176
rect 26172 15174 26196 15176
rect 25956 15154 26252 15174
rect 25956 14142 26252 14162
rect 26012 14140 26036 14142
rect 26092 14140 26116 14142
rect 26172 14140 26196 14142
rect 26034 14088 26036 14140
rect 26098 14088 26110 14140
rect 26172 14088 26174 14140
rect 26012 14086 26036 14088
rect 26092 14086 26116 14088
rect 26172 14086 26196 14088
rect 25956 14066 26252 14086
rect 25956 13054 26252 13074
rect 26012 13052 26036 13054
rect 26092 13052 26116 13054
rect 26172 13052 26196 13054
rect 26034 13000 26036 13052
rect 26098 13000 26110 13052
rect 26172 13000 26174 13052
rect 26012 12998 26036 13000
rect 26092 12998 26116 13000
rect 26172 12998 26196 13000
rect 25956 12978 26252 12998
rect 25956 11966 26252 11986
rect 26012 11964 26036 11966
rect 26092 11964 26116 11966
rect 26172 11964 26196 11966
rect 26034 11912 26036 11964
rect 26098 11912 26110 11964
rect 26172 11912 26174 11964
rect 26012 11910 26036 11912
rect 26092 11910 26116 11912
rect 26172 11910 26196 11912
rect 25956 11890 26252 11910
rect 25956 10878 26252 10898
rect 26012 10876 26036 10878
rect 26092 10876 26116 10878
rect 26172 10876 26196 10878
rect 26034 10824 26036 10876
rect 26098 10824 26110 10876
rect 26172 10824 26174 10876
rect 26012 10822 26036 10824
rect 26092 10822 26116 10824
rect 26172 10822 26196 10824
rect 25956 10802 26252 10822
rect 25956 9790 26252 9810
rect 26012 9788 26036 9790
rect 26092 9788 26116 9790
rect 26172 9788 26196 9790
rect 26034 9736 26036 9788
rect 26098 9736 26110 9788
rect 26172 9736 26174 9788
rect 26012 9734 26036 9736
rect 26092 9734 26116 9736
rect 26172 9734 26196 9736
rect 25956 9714 26252 9734
rect 25956 8702 26252 8722
rect 26012 8700 26036 8702
rect 26092 8700 26116 8702
rect 26172 8700 26196 8702
rect 26034 8648 26036 8700
rect 26098 8648 26110 8700
rect 26172 8648 26174 8700
rect 26012 8646 26036 8648
rect 26092 8646 26116 8648
rect 26172 8646 26196 8648
rect 25956 8626 26252 8646
rect 25956 7614 26252 7634
rect 26012 7612 26036 7614
rect 26092 7612 26116 7614
rect 26172 7612 26196 7614
rect 26034 7560 26036 7612
rect 26098 7560 26110 7612
rect 26172 7560 26174 7612
rect 26012 7558 26036 7560
rect 26092 7558 26116 7560
rect 26172 7558 26196 7560
rect 25956 7538 26252 7558
rect 25956 6526 26252 6546
rect 26012 6524 26036 6526
rect 26092 6524 26116 6526
rect 26172 6524 26196 6526
rect 26034 6472 26036 6524
rect 26098 6472 26110 6524
rect 26172 6472 26174 6524
rect 26012 6470 26036 6472
rect 26092 6470 26116 6472
rect 26172 6470 26196 6472
rect 25956 6450 26252 6470
rect 25956 5438 26252 5458
rect 26012 5436 26036 5438
rect 26092 5436 26116 5438
rect 26172 5436 26196 5438
rect 26034 5384 26036 5436
rect 26098 5384 26110 5436
rect 26172 5384 26174 5436
rect 26012 5382 26036 5384
rect 26092 5382 26116 5384
rect 26172 5382 26196 5384
rect 25956 5362 26252 5382
rect 25686 5234 25742 5243
rect 25686 5169 25742 5178
rect 25956 4350 26252 4370
rect 26012 4348 26036 4350
rect 26092 4348 26116 4350
rect 26172 4348 26196 4350
rect 26034 4296 26036 4348
rect 26098 4296 26110 4348
rect 26172 4296 26174 4348
rect 26012 4294 26036 4296
rect 26092 4294 26116 4296
rect 26172 4294 26196 4296
rect 25956 4274 26252 4294
rect 25956 3262 26252 3282
rect 26012 3260 26036 3262
rect 26092 3260 26116 3262
rect 26172 3260 26196 3262
rect 26034 3208 26036 3260
rect 26098 3208 26110 3260
rect 26172 3208 26174 3260
rect 26012 3206 26036 3208
rect 26092 3206 26116 3208
rect 26172 3206 26196 3208
rect 25956 3186 26252 3206
rect 25502 2378 25558 2387
rect 25502 2313 25558 2322
rect 25320 2274 25372 2280
rect 25320 2216 25372 2222
rect 24858 1562 24914 1571
rect 24858 1497 24914 1506
rect 25332 347 25360 2216
rect 25956 2174 26252 2194
rect 26012 2172 26036 2174
rect 26092 2172 26116 2174
rect 26172 2172 26196 2174
rect 26034 2120 26036 2172
rect 26098 2120 26110 2172
rect 26172 2120 26174 2172
rect 26012 2118 26036 2120
rect 26092 2118 26116 2120
rect 26172 2118 26196 2120
rect 25956 2098 26252 2118
rect 12346 338 12402 347
rect 12530 338 12586 347
rect 12402 296 12530 324
rect 12346 273 12402 282
rect 12530 273 12586 282
rect 25318 338 25374 347
rect 25318 273 25374 282
rect 9494 66 9550 75
rect 9494 1 9550 10
<< via2 >>
rect 3882 23538 3938 23594
rect 3330 22994 3386 23050
rect 3146 21226 3202 21282
rect 3238 18778 3294 18834
rect 2870 18234 2926 18290
rect 1398 15242 1454 15298
rect 1582 14018 1638 14074
rect 1490 13358 1546 13394
rect 1490 13338 1492 13358
rect 1492 13338 1544 13358
rect 1544 13338 1546 13358
rect 1398 9938 1454 9994
rect 1582 9838 1584 9858
rect 1584 9838 1636 9858
rect 1636 9838 1638 9858
rect 1582 9802 1638 9838
rect 1306 6266 1362 6322
rect 1674 2866 1730 2922
rect 2778 12794 2834 12850
rect 2226 12658 2282 12714
rect 2042 11182 2098 11218
rect 2042 11162 2044 11182
rect 2044 11162 2096 11182
rect 2096 11162 2098 11182
rect 1766 2594 1822 2650
rect 2042 2458 2098 2514
rect 2042 2358 2044 2378
rect 2044 2358 2096 2378
rect 2096 2358 2098 2378
rect 2042 2322 2098 2358
rect 1490 1370 1546 1426
rect 2410 11434 2466 11490
rect 2502 11298 2558 11354
rect 3054 15786 3110 15842
rect 2870 11706 2926 11762
rect 3514 22314 3570 22370
rect 3422 21770 3478 21826
rect 3330 18234 3386 18290
rect 3606 20002 3662 20058
rect 3514 17690 3570 17746
rect 3330 17554 3386 17610
rect 3238 13202 3294 13258
rect 3146 12250 3202 12306
rect 3514 17010 3570 17066
rect 3422 14562 3478 14618
rect 3422 13202 3478 13258
rect 3330 12250 3386 12306
rect 3238 12114 3294 12170
rect 3330 11570 3386 11626
rect 3146 10210 3202 10266
rect 3422 9530 3478 9586
rect 3790 19322 3846 19378
rect 3698 18914 3754 18970
rect 3698 9394 3754 9450
rect 24766 23538 24822 23594
rect 5956 21756 6012 21758
rect 6036 21756 6092 21758
rect 6116 21756 6172 21758
rect 6196 21756 6252 21758
rect 5956 21704 5982 21756
rect 5982 21704 6012 21756
rect 6036 21704 6046 21756
rect 6046 21704 6092 21756
rect 6116 21704 6162 21756
rect 6162 21704 6172 21756
rect 6196 21704 6226 21756
rect 6226 21704 6252 21756
rect 5956 21702 6012 21704
rect 6036 21702 6092 21704
rect 6116 21702 6172 21704
rect 6196 21702 6252 21704
rect 15956 21756 16012 21758
rect 16036 21756 16092 21758
rect 16116 21756 16172 21758
rect 16196 21756 16252 21758
rect 15956 21704 15982 21756
rect 15982 21704 16012 21756
rect 16036 21704 16046 21756
rect 16046 21704 16092 21756
rect 16116 21704 16162 21756
rect 16162 21704 16172 21756
rect 16196 21704 16226 21756
rect 16226 21704 16252 21756
rect 15956 21702 16012 21704
rect 16036 21702 16092 21704
rect 16116 21702 16172 21704
rect 16196 21702 16252 21704
rect 10956 21212 11012 21214
rect 11036 21212 11092 21214
rect 11116 21212 11172 21214
rect 11196 21212 11252 21214
rect 10956 21160 10982 21212
rect 10982 21160 11012 21212
rect 11036 21160 11046 21212
rect 11046 21160 11092 21212
rect 11116 21160 11162 21212
rect 11162 21160 11172 21212
rect 11196 21160 11226 21212
rect 11226 21160 11252 21212
rect 10956 21158 11012 21160
rect 11036 21158 11092 21160
rect 11116 21158 11172 21160
rect 11196 21158 11252 21160
rect 5956 20668 6012 20670
rect 6036 20668 6092 20670
rect 6116 20668 6172 20670
rect 6196 20668 6252 20670
rect 5956 20616 5982 20668
rect 5982 20616 6012 20668
rect 6036 20616 6046 20668
rect 6046 20616 6092 20668
rect 6116 20616 6162 20668
rect 6162 20616 6172 20668
rect 6196 20616 6226 20668
rect 6226 20616 6252 20668
rect 5956 20614 6012 20616
rect 6036 20614 6092 20616
rect 6116 20614 6172 20616
rect 6196 20614 6252 20616
rect 3974 20546 4030 20602
rect 3882 18778 3938 18834
rect 10956 20124 11012 20126
rect 11036 20124 11092 20126
rect 11116 20124 11172 20126
rect 11196 20124 11252 20126
rect 10956 20072 10982 20124
rect 10982 20072 11012 20124
rect 11036 20072 11046 20124
rect 11046 20072 11092 20124
rect 11116 20072 11162 20124
rect 11162 20072 11172 20124
rect 11196 20072 11226 20124
rect 11226 20072 11252 20124
rect 10956 20070 11012 20072
rect 11036 20070 11092 20072
rect 11116 20070 11172 20072
rect 11196 20070 11252 20072
rect 5956 19580 6012 19582
rect 6036 19580 6092 19582
rect 6116 19580 6172 19582
rect 6196 19580 6252 19582
rect 5956 19528 5982 19580
rect 5982 19528 6012 19580
rect 6036 19528 6046 19580
rect 6046 19528 6092 19580
rect 6116 19528 6162 19580
rect 6162 19528 6172 19580
rect 6196 19528 6226 19580
rect 6226 19528 6252 19580
rect 5956 19526 6012 19528
rect 6036 19526 6092 19528
rect 6116 19526 6172 19528
rect 6196 19526 6252 19528
rect 15956 20668 16012 20670
rect 16036 20668 16092 20670
rect 16116 20668 16172 20670
rect 16196 20668 16252 20670
rect 15956 20616 15982 20668
rect 15982 20616 16012 20668
rect 16036 20616 16046 20668
rect 16046 20616 16092 20668
rect 16116 20616 16162 20668
rect 16162 20616 16172 20668
rect 16196 20616 16226 20668
rect 16226 20616 16252 20668
rect 15956 20614 16012 20616
rect 16036 20614 16092 20616
rect 16116 20614 16172 20616
rect 16196 20614 16252 20616
rect 15956 19580 16012 19582
rect 16036 19580 16092 19582
rect 16116 19580 16172 19582
rect 16196 19580 16252 19582
rect 15956 19528 15982 19580
rect 15982 19528 16012 19580
rect 16036 19528 16046 19580
rect 16046 19528 16092 19580
rect 16116 19528 16162 19580
rect 16162 19528 16172 19580
rect 16196 19528 16226 19580
rect 16226 19528 16252 19580
rect 15956 19526 16012 19528
rect 16036 19526 16092 19528
rect 16116 19526 16172 19528
rect 16196 19526 16252 19528
rect 8850 19322 8906 19378
rect 11334 19322 11390 19378
rect 7010 18914 7066 18970
rect 8574 18914 8630 18970
rect 5956 18492 6012 18494
rect 6036 18492 6092 18494
rect 6116 18492 6172 18494
rect 6196 18492 6252 18494
rect 5956 18440 5982 18492
rect 5982 18440 6012 18492
rect 6036 18440 6046 18492
rect 6046 18440 6092 18492
rect 6116 18440 6162 18492
rect 6162 18440 6172 18492
rect 6196 18440 6226 18492
rect 6226 18440 6252 18492
rect 5956 18438 6012 18440
rect 6036 18438 6092 18440
rect 6116 18438 6172 18440
rect 6196 18438 6252 18440
rect 5956 17404 6012 17406
rect 6036 17404 6092 17406
rect 6116 17404 6172 17406
rect 6196 17404 6252 17406
rect 5956 17352 5982 17404
rect 5982 17352 6012 17404
rect 6036 17352 6046 17404
rect 6046 17352 6092 17404
rect 6116 17352 6162 17404
rect 6162 17352 6172 17404
rect 6196 17352 6226 17404
rect 6226 17352 6252 17404
rect 5956 17350 6012 17352
rect 6036 17350 6092 17352
rect 6116 17350 6172 17352
rect 6196 17350 6252 17352
rect 4066 16330 4122 16386
rect 3974 8986 4030 9042
rect 3882 7762 3938 7818
rect 5956 16316 6012 16318
rect 6036 16316 6092 16318
rect 6116 16316 6172 16318
rect 6196 16316 6252 16318
rect 5956 16264 5982 16316
rect 5982 16264 6012 16316
rect 6036 16264 6046 16316
rect 6046 16264 6092 16316
rect 6116 16264 6162 16316
rect 6162 16264 6172 16316
rect 6196 16264 6226 16316
rect 6226 16264 6252 16316
rect 5956 16262 6012 16264
rect 6036 16262 6092 16264
rect 6116 16262 6172 16264
rect 6196 16262 6252 16264
rect 10956 19036 11012 19038
rect 11036 19036 11092 19038
rect 11116 19036 11172 19038
rect 11196 19036 11252 19038
rect 10956 18984 10982 19036
rect 10982 18984 11012 19036
rect 11036 18984 11046 19036
rect 11046 18984 11092 19036
rect 11116 18984 11162 19036
rect 11162 18984 11172 19036
rect 11196 18984 11226 19036
rect 11226 18984 11252 19036
rect 10956 18982 11012 18984
rect 11036 18982 11092 18984
rect 11116 18982 11172 18984
rect 11196 18982 11252 18984
rect 24398 22314 24454 22370
rect 20956 21212 21012 21214
rect 21036 21212 21092 21214
rect 21116 21212 21172 21214
rect 21196 21212 21252 21214
rect 20956 21160 20982 21212
rect 20982 21160 21012 21212
rect 21036 21160 21046 21212
rect 21046 21160 21092 21212
rect 21116 21160 21162 21212
rect 21162 21160 21172 21212
rect 21196 21160 21226 21212
rect 21226 21160 21252 21212
rect 20956 21158 21012 21160
rect 21036 21158 21092 21160
rect 21116 21158 21172 21160
rect 21196 21158 21252 21160
rect 16762 18934 16818 18970
rect 16762 18914 16764 18934
rect 16764 18914 16816 18934
rect 16816 18914 16818 18934
rect 18694 18914 18750 18970
rect 8574 18098 8630 18154
rect 13082 18098 13138 18154
rect 15382 18134 15384 18154
rect 15384 18134 15436 18154
rect 15436 18134 15438 18154
rect 10956 17948 11012 17950
rect 11036 17948 11092 17950
rect 11116 17948 11172 17950
rect 11196 17948 11252 17950
rect 10956 17896 10982 17948
rect 10982 17896 11012 17948
rect 11036 17896 11046 17948
rect 11046 17896 11092 17948
rect 11116 17896 11162 17948
rect 11162 17896 11172 17948
rect 11196 17896 11226 17948
rect 11226 17896 11252 17948
rect 10956 17894 11012 17896
rect 11036 17894 11092 17896
rect 11116 17894 11172 17896
rect 11196 17894 11252 17896
rect 10956 16860 11012 16862
rect 11036 16860 11092 16862
rect 11116 16860 11172 16862
rect 11196 16860 11252 16862
rect 10956 16808 10982 16860
rect 10982 16808 11012 16860
rect 11036 16808 11046 16860
rect 11046 16808 11092 16860
rect 11116 16808 11162 16860
rect 11162 16808 11172 16860
rect 11196 16808 11226 16860
rect 11226 16808 11252 16860
rect 10956 16806 11012 16808
rect 11036 16806 11092 16808
rect 11116 16806 11172 16808
rect 11196 16806 11252 16808
rect 15382 18098 15438 18134
rect 15956 18492 16012 18494
rect 16036 18492 16092 18494
rect 16116 18492 16172 18494
rect 16196 18492 16252 18494
rect 15956 18440 15982 18492
rect 15982 18440 16012 18492
rect 16036 18440 16046 18492
rect 16046 18440 16092 18492
rect 16116 18440 16162 18492
rect 16162 18440 16172 18492
rect 16196 18440 16226 18492
rect 16226 18440 16252 18492
rect 15956 18438 16012 18440
rect 16036 18438 16092 18440
rect 16116 18438 16172 18440
rect 16196 18438 16252 18440
rect 13542 16874 13598 16930
rect 7194 15942 7250 15978
rect 7194 15922 7196 15942
rect 7196 15922 7248 15942
rect 7248 15922 7250 15942
rect 9954 15922 10010 15978
rect 5956 15228 6012 15230
rect 6036 15228 6092 15230
rect 6116 15228 6172 15230
rect 6196 15228 6252 15230
rect 5956 15176 5982 15228
rect 5982 15176 6012 15228
rect 6036 15176 6046 15228
rect 6046 15176 6092 15228
rect 6116 15176 6162 15228
rect 6162 15176 6172 15228
rect 6196 15176 6226 15228
rect 6226 15176 6252 15228
rect 5956 15174 6012 15176
rect 6036 15174 6092 15176
rect 6116 15174 6172 15176
rect 6196 15174 6252 15176
rect 5956 14140 6012 14142
rect 6036 14140 6092 14142
rect 6116 14140 6172 14142
rect 6196 14140 6252 14142
rect 5956 14088 5982 14140
rect 5982 14088 6012 14140
rect 6036 14088 6046 14140
rect 6046 14088 6092 14140
rect 6116 14088 6162 14140
rect 6162 14088 6172 14140
rect 6196 14088 6226 14140
rect 6226 14088 6252 14140
rect 5956 14086 6012 14088
rect 6036 14086 6092 14088
rect 6116 14086 6172 14088
rect 6196 14086 6252 14088
rect 5956 13052 6012 13054
rect 6036 13052 6092 13054
rect 6116 13052 6172 13054
rect 6196 13052 6252 13054
rect 5956 13000 5982 13052
rect 5982 13000 6012 13052
rect 6036 13000 6046 13052
rect 6046 13000 6092 13052
rect 6116 13000 6162 13052
rect 6162 13000 6172 13052
rect 6196 13000 6226 13052
rect 6226 13000 6252 13052
rect 5956 12998 6012 13000
rect 6036 12998 6092 13000
rect 6116 12998 6172 13000
rect 6196 12998 6252 13000
rect 5956 11964 6012 11966
rect 6036 11964 6092 11966
rect 6116 11964 6172 11966
rect 6196 11964 6252 11966
rect 5956 11912 5982 11964
rect 5982 11912 6012 11964
rect 6036 11912 6046 11964
rect 6046 11912 6092 11964
rect 6116 11912 6162 11964
rect 6162 11912 6172 11964
rect 6196 11912 6226 11964
rect 6226 11912 6252 11964
rect 5956 11910 6012 11912
rect 6036 11910 6092 11912
rect 6116 11910 6172 11912
rect 6196 11910 6252 11912
rect 7102 11298 7158 11354
rect 5956 10876 6012 10878
rect 6036 10876 6092 10878
rect 6116 10876 6172 10878
rect 6196 10876 6252 10878
rect 5956 10824 5982 10876
rect 5982 10824 6012 10876
rect 6036 10824 6046 10876
rect 6046 10824 6092 10876
rect 6116 10824 6162 10876
rect 6162 10824 6172 10876
rect 6196 10824 6226 10876
rect 6226 10824 6252 10876
rect 5956 10822 6012 10824
rect 6036 10822 6092 10824
rect 6116 10822 6172 10824
rect 6196 10822 6252 10824
rect 10956 15772 11012 15774
rect 11036 15772 11092 15774
rect 11116 15772 11172 15774
rect 11196 15772 11252 15774
rect 10956 15720 10982 15772
rect 10982 15720 11012 15772
rect 11036 15720 11046 15772
rect 11046 15720 11092 15772
rect 11116 15720 11162 15772
rect 11162 15720 11172 15772
rect 11196 15720 11226 15772
rect 11226 15720 11252 15772
rect 10956 15718 11012 15720
rect 11036 15718 11092 15720
rect 11116 15718 11172 15720
rect 11196 15718 11252 15720
rect 8482 15106 8538 15162
rect 13450 15106 13506 15162
rect 7378 12114 7434 12170
rect 7930 12134 7986 12170
rect 7930 12114 7932 12134
rect 7932 12114 7984 12134
rect 7984 12114 7986 12134
rect 8114 11706 8170 11762
rect 10956 14684 11012 14686
rect 11036 14684 11092 14686
rect 11116 14684 11172 14686
rect 11196 14684 11252 14686
rect 10956 14632 10982 14684
rect 10982 14632 11012 14684
rect 11036 14632 11046 14684
rect 11046 14632 11092 14684
rect 11116 14632 11162 14684
rect 11162 14632 11172 14684
rect 11196 14632 11226 14684
rect 11226 14632 11252 14684
rect 10956 14630 11012 14632
rect 11036 14630 11092 14632
rect 11116 14630 11172 14632
rect 11196 14630 11252 14632
rect 13450 14426 13506 14482
rect 10956 13596 11012 13598
rect 11036 13596 11092 13598
rect 11116 13596 11172 13598
rect 11196 13596 11252 13598
rect 10956 13544 10982 13596
rect 10982 13544 11012 13596
rect 11036 13544 11046 13596
rect 11046 13544 11092 13596
rect 11116 13544 11162 13596
rect 11162 13544 11172 13596
rect 11196 13544 11226 13596
rect 11226 13544 11252 13596
rect 10956 13542 11012 13544
rect 11036 13542 11092 13544
rect 11116 13542 11172 13544
rect 11196 13542 11252 13544
rect 11978 13202 12034 13258
rect 10956 12508 11012 12510
rect 11036 12508 11092 12510
rect 11116 12508 11172 12510
rect 11196 12508 11252 12510
rect 10956 12456 10982 12508
rect 10982 12456 11012 12508
rect 11036 12456 11046 12508
rect 11046 12456 11092 12508
rect 11116 12456 11162 12508
rect 11162 12456 11172 12508
rect 11196 12456 11226 12508
rect 11226 12456 11252 12508
rect 10956 12454 11012 12456
rect 11036 12454 11092 12456
rect 11116 12454 11172 12456
rect 11196 12454 11252 12456
rect 15956 17404 16012 17406
rect 16036 17404 16092 17406
rect 16116 17404 16172 17406
rect 16196 17404 16252 17406
rect 15956 17352 15982 17404
rect 15982 17352 16012 17404
rect 16036 17352 16046 17404
rect 16046 17352 16092 17404
rect 16116 17352 16162 17404
rect 16162 17352 16172 17404
rect 16196 17352 16226 17404
rect 16226 17352 16252 17404
rect 15956 17350 16012 17352
rect 16036 17350 16092 17352
rect 16116 17350 16172 17352
rect 16196 17350 16252 17352
rect 17498 16910 17500 16930
rect 17500 16910 17552 16930
rect 17552 16910 17554 16930
rect 17498 16874 17554 16910
rect 15956 16316 16012 16318
rect 16036 16316 16092 16318
rect 16116 16316 16172 16318
rect 16196 16316 16252 16318
rect 15956 16264 15982 16316
rect 15982 16264 16012 16316
rect 16036 16264 16046 16316
rect 16046 16264 16092 16316
rect 16116 16264 16162 16316
rect 16162 16264 16172 16316
rect 16196 16264 16226 16316
rect 16226 16264 16252 16316
rect 15956 16262 16012 16264
rect 16036 16262 16092 16264
rect 16116 16262 16172 16264
rect 16196 16262 16252 16264
rect 15956 15228 16012 15230
rect 16036 15228 16092 15230
rect 16116 15228 16172 15230
rect 16196 15228 16252 15230
rect 15956 15176 15982 15228
rect 15982 15176 16012 15228
rect 16036 15176 16046 15228
rect 16046 15176 16092 15228
rect 16116 15176 16162 15228
rect 16162 15176 16172 15228
rect 16196 15176 16226 15228
rect 16226 15176 16252 15228
rect 15956 15174 16012 15176
rect 16036 15174 16092 15176
rect 16116 15174 16172 15176
rect 16196 15174 16252 15176
rect 14094 14970 14150 15026
rect 18786 14990 18842 15026
rect 18786 14970 18788 14990
rect 18788 14970 18840 14990
rect 18840 14970 18842 14990
rect 15956 14140 16012 14142
rect 16036 14140 16092 14142
rect 16116 14140 16172 14142
rect 16196 14140 16252 14142
rect 15956 14088 15982 14140
rect 15982 14088 16012 14140
rect 16036 14088 16046 14140
rect 16046 14088 16092 14140
rect 16116 14088 16162 14140
rect 16162 14088 16172 14140
rect 16196 14088 16226 14140
rect 16226 14088 16252 14140
rect 15956 14086 16012 14088
rect 16036 14086 16092 14088
rect 16116 14086 16172 14088
rect 16196 14086 16252 14088
rect 19522 13474 19578 13530
rect 15956 13052 16012 13054
rect 16036 13052 16092 13054
rect 16116 13052 16172 13054
rect 16196 13052 16252 13054
rect 15956 13000 15982 13052
rect 15982 13000 16012 13052
rect 16036 13000 16046 13052
rect 16046 13000 16092 13052
rect 16116 13000 16162 13052
rect 16162 13000 16172 13052
rect 16196 13000 16226 13052
rect 16226 13000 16252 13052
rect 15956 12998 16012 13000
rect 16036 12998 16092 13000
rect 16116 12998 16172 13000
rect 16196 12998 16252 13000
rect 24030 20410 24086 20466
rect 20956 20124 21012 20126
rect 21036 20124 21092 20126
rect 21116 20124 21172 20126
rect 21196 20124 21252 20126
rect 20956 20072 20982 20124
rect 20982 20072 21012 20124
rect 21036 20072 21046 20124
rect 21046 20072 21092 20124
rect 21116 20072 21162 20124
rect 21162 20072 21172 20124
rect 21196 20072 21226 20124
rect 21226 20072 21252 20124
rect 20956 20070 21012 20072
rect 21036 20070 21092 20072
rect 21116 20070 21172 20072
rect 21196 20070 21252 20072
rect 20810 19186 20866 19242
rect 20956 19036 21012 19038
rect 21036 19036 21092 19038
rect 21116 19036 21172 19038
rect 21196 19036 21252 19038
rect 20956 18984 20982 19036
rect 20982 18984 21012 19036
rect 21036 18984 21046 19036
rect 21046 18984 21092 19036
rect 21116 18984 21162 19036
rect 21162 18984 21172 19036
rect 21196 18984 21226 19036
rect 21226 18984 21252 19036
rect 20956 18982 21012 18984
rect 21036 18982 21092 18984
rect 21116 18982 21172 18984
rect 21196 18982 21252 18984
rect 19890 18370 19946 18426
rect 20956 17948 21012 17950
rect 21036 17948 21092 17950
rect 21116 17948 21172 17950
rect 21196 17948 21252 17950
rect 20956 17896 20982 17948
rect 20982 17896 21012 17948
rect 21036 17896 21046 17948
rect 21046 17896 21092 17948
rect 21116 17896 21162 17948
rect 21162 17896 21172 17948
rect 21196 17896 21226 17948
rect 21226 17896 21252 17948
rect 20956 17894 21012 17896
rect 21036 17894 21092 17896
rect 21116 17894 21172 17896
rect 21196 17894 21252 17896
rect 20956 16860 21012 16862
rect 21036 16860 21092 16862
rect 21116 16860 21172 16862
rect 21196 16860 21252 16862
rect 20956 16808 20982 16860
rect 20982 16808 21012 16860
rect 21036 16808 21046 16860
rect 21046 16808 21092 16860
rect 21116 16808 21162 16860
rect 21162 16808 21172 16860
rect 21196 16808 21226 16860
rect 21226 16808 21252 16860
rect 20956 16806 21012 16808
rect 21036 16806 21092 16808
rect 21116 16806 21172 16808
rect 21196 16806 21252 16808
rect 21454 15786 21510 15842
rect 20956 15772 21012 15774
rect 21036 15772 21092 15774
rect 21116 15772 21172 15774
rect 21196 15772 21252 15774
rect 20956 15720 20982 15772
rect 20982 15720 21012 15772
rect 21036 15720 21046 15772
rect 21046 15720 21092 15772
rect 21116 15720 21162 15772
rect 21162 15720 21172 15772
rect 21196 15720 21226 15772
rect 21226 15720 21252 15772
rect 20956 15718 21012 15720
rect 21036 15718 21092 15720
rect 21116 15718 21172 15720
rect 21196 15718 21252 15720
rect 20956 14684 21012 14686
rect 21036 14684 21092 14686
rect 21116 14684 21172 14686
rect 21196 14684 21252 14686
rect 20956 14632 20982 14684
rect 20982 14632 21012 14684
rect 21036 14632 21046 14684
rect 21046 14632 21092 14684
rect 21116 14632 21162 14684
rect 21162 14632 21172 14684
rect 21196 14632 21226 14684
rect 21226 14632 21252 14684
rect 20956 14630 21012 14632
rect 21036 14630 21092 14632
rect 21116 14630 21172 14632
rect 21196 14630 21252 14632
rect 19982 14426 20038 14482
rect 19706 13338 19762 13394
rect 20956 13596 21012 13598
rect 21036 13596 21092 13598
rect 21116 13596 21172 13598
rect 21196 13596 21252 13598
rect 20956 13544 20982 13596
rect 20982 13544 21012 13596
rect 21036 13544 21046 13596
rect 21046 13544 21092 13596
rect 21116 13544 21162 13596
rect 21162 13544 21172 13596
rect 21196 13544 21226 13596
rect 21226 13544 21252 13596
rect 20956 13542 21012 13544
rect 21036 13542 21092 13544
rect 21116 13542 21172 13544
rect 21196 13542 21252 13544
rect 19154 12694 19156 12714
rect 19156 12694 19208 12714
rect 19208 12694 19210 12714
rect 19154 12658 19210 12694
rect 20956 12508 21012 12510
rect 21036 12508 21092 12510
rect 21116 12508 21172 12510
rect 21196 12508 21252 12510
rect 20956 12456 20982 12508
rect 20982 12456 21012 12508
rect 21036 12456 21046 12508
rect 21046 12456 21092 12508
rect 21116 12456 21162 12508
rect 21162 12456 21172 12508
rect 21196 12456 21226 12508
rect 21226 12456 21252 12508
rect 20956 12454 21012 12456
rect 21036 12454 21092 12456
rect 21116 12454 21172 12456
rect 21196 12454 21252 12456
rect 13082 11842 13138 11898
rect 13910 12114 13966 12170
rect 15956 11964 16012 11966
rect 16036 11964 16092 11966
rect 16116 11964 16172 11966
rect 16196 11964 16252 11966
rect 15956 11912 15982 11964
rect 15982 11912 16012 11964
rect 16036 11912 16046 11964
rect 16046 11912 16092 11964
rect 16116 11912 16162 11964
rect 16162 11912 16172 11964
rect 16196 11912 16226 11964
rect 16226 11912 16252 11964
rect 15956 11910 16012 11912
rect 16036 11910 16092 11912
rect 16116 11910 16172 11912
rect 16196 11910 16252 11912
rect 14738 11842 14794 11898
rect 8114 11298 8170 11354
rect 10956 11420 11012 11422
rect 11036 11420 11092 11422
rect 11116 11420 11172 11422
rect 11196 11420 11252 11422
rect 10956 11368 10982 11420
rect 10982 11368 11012 11420
rect 11036 11368 11046 11420
rect 11046 11368 11092 11420
rect 11116 11368 11162 11420
rect 11162 11368 11172 11420
rect 11196 11368 11226 11420
rect 11226 11368 11252 11420
rect 10956 11366 11012 11368
rect 11036 11366 11092 11368
rect 11116 11366 11172 11368
rect 11196 11366 11252 11368
rect 12162 11570 12218 11626
rect 8298 11062 8300 11082
rect 8300 11062 8352 11082
rect 8352 11062 8354 11082
rect 8298 11026 8354 11062
rect 12070 11026 12126 11082
rect 8298 10502 8354 10538
rect 8298 10482 8300 10502
rect 8300 10482 8352 10502
rect 8352 10482 8354 10502
rect 5956 9788 6012 9790
rect 6036 9788 6092 9790
rect 6116 9788 6172 9790
rect 6196 9788 6252 9790
rect 5956 9736 5982 9788
rect 5982 9736 6012 9788
rect 6036 9736 6046 9788
rect 6046 9736 6092 9788
rect 6116 9736 6162 9788
rect 6162 9736 6172 9788
rect 6196 9736 6226 9788
rect 6226 9736 6252 9788
rect 5956 9734 6012 9736
rect 6036 9734 6092 9736
rect 6116 9734 6172 9736
rect 6196 9734 6252 9736
rect 4158 9530 4214 9586
rect 3790 7354 3846 7410
rect 3606 7218 3662 7274
rect 3514 5178 3570 5234
rect 5956 8700 6012 8702
rect 6036 8700 6092 8702
rect 6116 8700 6172 8702
rect 6196 8700 6252 8702
rect 5956 8648 5982 8700
rect 5982 8648 6012 8700
rect 6036 8648 6046 8700
rect 6046 8648 6092 8700
rect 6116 8648 6162 8700
rect 6162 8648 6172 8700
rect 6196 8648 6226 8700
rect 6226 8648 6252 8700
rect 5956 8646 6012 8648
rect 6036 8646 6092 8648
rect 6116 8646 6172 8648
rect 6196 8646 6252 8648
rect 5956 7612 6012 7614
rect 6036 7612 6092 7614
rect 6116 7612 6172 7614
rect 6196 7612 6252 7614
rect 5956 7560 5982 7612
rect 5982 7560 6012 7612
rect 6036 7560 6046 7612
rect 6046 7560 6092 7612
rect 6116 7560 6162 7612
rect 6162 7560 6172 7612
rect 6196 7560 6226 7612
rect 6226 7560 6252 7612
rect 5956 7558 6012 7560
rect 6036 7558 6092 7560
rect 6116 7558 6172 7560
rect 6196 7558 6252 7560
rect 5956 6524 6012 6526
rect 6036 6524 6092 6526
rect 6116 6524 6172 6526
rect 6196 6524 6252 6526
rect 5956 6472 5982 6524
rect 5982 6472 6012 6524
rect 6036 6472 6046 6524
rect 6046 6472 6092 6524
rect 6116 6472 6162 6524
rect 6162 6472 6172 6524
rect 6196 6472 6226 6524
rect 6226 6472 6252 6524
rect 5956 6470 6012 6472
rect 6036 6470 6092 6472
rect 6116 6470 6172 6472
rect 6196 6470 6252 6472
rect 4342 5606 4398 5642
rect 4342 5586 4344 5606
rect 4344 5586 4396 5606
rect 4396 5586 4398 5606
rect 5956 5436 6012 5438
rect 6036 5436 6092 5438
rect 6116 5436 6172 5438
rect 6196 5436 6252 5438
rect 5956 5384 5982 5436
rect 5982 5384 6012 5436
rect 6036 5384 6046 5436
rect 6046 5384 6092 5436
rect 6116 5384 6162 5436
rect 6162 5384 6172 5436
rect 6196 5384 6226 5436
rect 6226 5384 6252 5436
rect 5956 5382 6012 5384
rect 6036 5382 6092 5384
rect 6116 5382 6172 5384
rect 6196 5382 6252 5384
rect 3882 4634 3938 4690
rect 5956 4348 6012 4350
rect 6036 4348 6092 4350
rect 6116 4348 6172 4350
rect 6196 4348 6252 4350
rect 5956 4296 5982 4348
rect 5982 4296 6012 4348
rect 6036 4296 6046 4348
rect 6046 4296 6092 4348
rect 6116 4296 6162 4348
rect 6162 4296 6172 4348
rect 6196 4296 6226 4348
rect 6226 4296 6252 4348
rect 5956 4294 6012 4296
rect 6036 4294 6092 4296
rect 6116 4294 6172 4296
rect 6196 4294 6252 4296
rect 3422 3954 3478 4010
rect 5956 3260 6012 3262
rect 6036 3260 6092 3262
rect 6116 3260 6172 3262
rect 6196 3260 6252 3262
rect 5956 3208 5982 3260
rect 5982 3208 6012 3260
rect 6036 3208 6046 3260
rect 6046 3208 6092 3260
rect 6116 3208 6162 3260
rect 6162 3208 6172 3260
rect 6196 3208 6226 3260
rect 6226 3208 6252 3260
rect 5956 3206 6012 3208
rect 6036 3206 6092 3208
rect 6116 3206 6172 3208
rect 6196 3206 6252 3208
rect 7838 10210 7894 10266
rect 8298 9938 8354 9994
rect 7378 3002 7434 3058
rect 10956 10332 11012 10334
rect 11036 10332 11092 10334
rect 11116 10332 11172 10334
rect 11196 10332 11252 10334
rect 10956 10280 10982 10332
rect 10982 10280 11012 10332
rect 11036 10280 11046 10332
rect 11046 10280 11092 10332
rect 11116 10280 11162 10332
rect 11162 10280 11172 10332
rect 11196 10280 11226 10332
rect 11226 10280 11252 10332
rect 10956 10278 11012 10280
rect 11036 10278 11092 10280
rect 11116 10278 11172 10280
rect 11196 10278 11252 10280
rect 10956 9244 11012 9246
rect 11036 9244 11092 9246
rect 11116 9244 11172 9246
rect 11196 9244 11252 9246
rect 10956 9192 10982 9244
rect 10982 9192 11012 9244
rect 11036 9192 11046 9244
rect 11046 9192 11092 9244
rect 11116 9192 11162 9244
rect 11162 9192 11172 9244
rect 11196 9192 11226 9244
rect 11226 9192 11252 9244
rect 10956 9190 11012 9192
rect 11036 9190 11092 9192
rect 11116 9190 11172 9192
rect 11196 9190 11252 9192
rect 10956 8156 11012 8158
rect 11036 8156 11092 8158
rect 11116 8156 11172 8158
rect 11196 8156 11252 8158
rect 10956 8104 10982 8156
rect 10982 8104 11012 8156
rect 11036 8104 11046 8156
rect 11046 8104 11092 8156
rect 11116 8104 11162 8156
rect 11162 8104 11172 8156
rect 11196 8104 11226 8156
rect 11226 8104 11252 8156
rect 10956 8102 11012 8104
rect 11036 8102 11092 8104
rect 11116 8102 11172 8104
rect 11196 8102 11252 8104
rect 10956 7068 11012 7070
rect 11036 7068 11092 7070
rect 11116 7068 11172 7070
rect 11196 7068 11252 7070
rect 10956 7016 10982 7068
rect 10982 7016 11012 7068
rect 11036 7016 11046 7068
rect 11046 7016 11092 7068
rect 11116 7016 11162 7068
rect 11162 7016 11172 7068
rect 11196 7016 11226 7068
rect 11226 7016 11252 7068
rect 10956 7014 11012 7016
rect 11036 7014 11092 7016
rect 11116 7014 11172 7016
rect 11196 7014 11252 7016
rect 13082 7762 13138 7818
rect 13266 7118 13268 7138
rect 13268 7118 13320 7138
rect 13320 7118 13322 7138
rect 13266 7082 13322 7118
rect 20956 11420 21012 11422
rect 21036 11420 21092 11422
rect 21116 11420 21172 11422
rect 21196 11420 21252 11422
rect 20956 11368 20982 11420
rect 20982 11368 21012 11420
rect 21036 11368 21046 11420
rect 21046 11368 21092 11420
rect 21116 11368 21162 11420
rect 21162 11368 21172 11420
rect 21196 11368 21226 11420
rect 21226 11368 21252 11420
rect 20956 11366 21012 11368
rect 21036 11366 21092 11368
rect 21116 11366 21172 11368
rect 21196 11366 21252 11368
rect 15956 10876 16012 10878
rect 16036 10876 16092 10878
rect 16116 10876 16172 10878
rect 16196 10876 16252 10878
rect 15956 10824 15982 10876
rect 15982 10824 16012 10876
rect 16036 10824 16046 10876
rect 16046 10824 16092 10876
rect 16116 10824 16162 10876
rect 16162 10824 16172 10876
rect 16196 10824 16226 10876
rect 16226 10824 16252 10876
rect 15956 10822 16012 10824
rect 16036 10822 16092 10824
rect 16116 10822 16172 10824
rect 16196 10822 16252 10824
rect 20956 10332 21012 10334
rect 21036 10332 21092 10334
rect 21116 10332 21172 10334
rect 21196 10332 21252 10334
rect 20956 10280 20982 10332
rect 20982 10280 21012 10332
rect 21036 10280 21046 10332
rect 21046 10280 21092 10332
rect 21116 10280 21162 10332
rect 21162 10280 21172 10332
rect 21196 10280 21226 10332
rect 21226 10280 21252 10332
rect 20956 10278 21012 10280
rect 21036 10278 21092 10280
rect 21116 10278 21172 10280
rect 21196 10278 21252 10280
rect 15956 9788 16012 9790
rect 16036 9788 16092 9790
rect 16116 9788 16172 9790
rect 16196 9788 16252 9790
rect 15956 9736 15982 9788
rect 15982 9736 16012 9788
rect 16036 9736 16046 9788
rect 16046 9736 16092 9788
rect 16116 9736 16162 9788
rect 16162 9736 16172 9788
rect 16196 9736 16226 9788
rect 16226 9736 16252 9788
rect 15956 9734 16012 9736
rect 16036 9734 16092 9736
rect 16116 9734 16172 9736
rect 16196 9734 16252 9736
rect 20956 9244 21012 9246
rect 21036 9244 21092 9246
rect 21116 9244 21172 9246
rect 21196 9244 21252 9246
rect 20956 9192 20982 9244
rect 20982 9192 21012 9244
rect 21036 9192 21046 9244
rect 21046 9192 21092 9244
rect 21116 9192 21162 9244
rect 21162 9192 21172 9244
rect 21196 9192 21226 9244
rect 21226 9192 21252 9244
rect 20956 9190 21012 9192
rect 21036 9190 21092 9192
rect 21116 9190 21172 9192
rect 21196 9190 21252 9192
rect 15956 8700 16012 8702
rect 16036 8700 16092 8702
rect 16116 8700 16172 8702
rect 16196 8700 16252 8702
rect 15956 8648 15982 8700
rect 15982 8648 16012 8700
rect 16036 8648 16046 8700
rect 16046 8648 16092 8700
rect 16116 8648 16162 8700
rect 16162 8648 16172 8700
rect 16196 8648 16226 8700
rect 16226 8648 16252 8700
rect 15956 8646 16012 8648
rect 16036 8646 16092 8648
rect 16116 8646 16172 8648
rect 16196 8646 16252 8648
rect 20956 8156 21012 8158
rect 21036 8156 21092 8158
rect 21116 8156 21172 8158
rect 21196 8156 21252 8158
rect 20956 8104 20982 8156
rect 20982 8104 21012 8156
rect 21036 8104 21046 8156
rect 21046 8104 21092 8156
rect 21116 8104 21162 8156
rect 21162 8104 21172 8156
rect 21196 8104 21226 8156
rect 21226 8104 21252 8156
rect 20956 8102 21012 8104
rect 21036 8102 21092 8104
rect 21116 8102 21172 8104
rect 21196 8102 21252 8104
rect 15956 7612 16012 7614
rect 16036 7612 16092 7614
rect 16116 7612 16172 7614
rect 16196 7612 16252 7614
rect 15956 7560 15982 7612
rect 15982 7560 16012 7612
rect 16036 7560 16046 7612
rect 16046 7560 16092 7612
rect 16116 7560 16162 7612
rect 16162 7560 16172 7612
rect 16196 7560 16226 7612
rect 16226 7560 16252 7612
rect 15956 7558 16012 7560
rect 16036 7558 16092 7560
rect 16116 7558 16172 7560
rect 16196 7558 16252 7560
rect 20534 7490 20590 7546
rect 18418 7354 18474 7410
rect 18602 7390 18604 7410
rect 18604 7390 18656 7410
rect 18656 7390 18658 7410
rect 18602 7354 18658 7390
rect 20534 7218 20590 7274
rect 20956 7068 21012 7070
rect 21036 7068 21092 7070
rect 21116 7068 21172 7070
rect 21196 7068 21252 7070
rect 20956 7016 20982 7068
rect 20982 7016 21012 7068
rect 21036 7016 21046 7068
rect 21046 7016 21092 7068
rect 21116 7016 21162 7068
rect 21162 7016 21172 7068
rect 21196 7016 21226 7068
rect 21226 7016 21252 7068
rect 20956 7014 21012 7016
rect 21036 7014 21092 7016
rect 21116 7014 21172 7016
rect 21196 7014 21252 7016
rect 10956 5980 11012 5982
rect 11036 5980 11092 5982
rect 11116 5980 11172 5982
rect 11196 5980 11252 5982
rect 10956 5928 10982 5980
rect 10982 5928 11012 5980
rect 11036 5928 11046 5980
rect 11046 5928 11092 5980
rect 11116 5928 11162 5980
rect 11162 5928 11172 5980
rect 11196 5928 11226 5980
rect 11226 5928 11252 5980
rect 10956 5926 11012 5928
rect 11036 5926 11092 5928
rect 11116 5926 11172 5928
rect 11196 5926 11252 5928
rect 12622 5178 12678 5234
rect 10956 4892 11012 4894
rect 11036 4892 11092 4894
rect 11116 4892 11172 4894
rect 11196 4892 11252 4894
rect 10956 4840 10982 4892
rect 10982 4840 11012 4892
rect 11036 4840 11046 4892
rect 11046 4840 11092 4892
rect 11116 4840 11162 4892
rect 11162 4840 11172 4892
rect 11196 4840 11226 4892
rect 11226 4840 11252 4892
rect 10956 4838 11012 4840
rect 11036 4838 11092 4840
rect 11116 4838 11172 4840
rect 11196 4838 11252 4840
rect 10956 3804 11012 3806
rect 11036 3804 11092 3806
rect 11116 3804 11172 3806
rect 11196 3804 11252 3806
rect 10956 3752 10982 3804
rect 10982 3752 11012 3804
rect 11036 3752 11046 3804
rect 11046 3752 11092 3804
rect 11116 3752 11162 3804
rect 11162 3752 11172 3804
rect 11196 3752 11226 3804
rect 11226 3752 11252 3804
rect 10956 3750 11012 3752
rect 11036 3750 11092 3752
rect 11116 3750 11172 3752
rect 11196 3750 11252 3752
rect 8390 2458 8446 2514
rect 5956 2172 6012 2174
rect 6036 2172 6092 2174
rect 6116 2172 6172 2174
rect 6196 2172 6252 2174
rect 5956 2120 5982 2172
rect 5982 2120 6012 2172
rect 6036 2120 6046 2172
rect 6046 2120 6092 2172
rect 6116 2120 6162 2172
rect 6162 2120 6172 2172
rect 6196 2120 6226 2172
rect 6226 2120 6252 2172
rect 5956 2118 6012 2120
rect 6036 2118 6092 2120
rect 6116 2118 6172 2120
rect 6196 2118 6252 2120
rect 2134 1370 2190 1426
rect 1582 826 1638 882
rect 1398 282 1454 338
rect 10956 2716 11012 2718
rect 11036 2716 11092 2718
rect 11116 2716 11172 2718
rect 11196 2716 11252 2718
rect 10956 2664 10982 2716
rect 10982 2664 11012 2716
rect 11036 2664 11046 2716
rect 11046 2664 11092 2716
rect 11116 2664 11162 2716
rect 11162 2664 11172 2716
rect 11196 2664 11226 2716
rect 11226 2664 11252 2716
rect 10956 2662 11012 2664
rect 11036 2662 11092 2664
rect 11116 2662 11172 2664
rect 11196 2662 11252 2664
rect 14922 6810 14978 6866
rect 15956 6524 16012 6526
rect 16036 6524 16092 6526
rect 16116 6524 16172 6526
rect 16196 6524 16252 6526
rect 15956 6472 15982 6524
rect 15982 6472 16012 6524
rect 16036 6472 16046 6524
rect 16046 6472 16092 6524
rect 16116 6472 16162 6524
rect 16162 6472 16172 6524
rect 16196 6472 16226 6524
rect 16226 6472 16252 6524
rect 15956 6470 16012 6472
rect 16036 6470 16092 6472
rect 16116 6470 16172 6472
rect 16196 6470 16252 6472
rect 20956 5980 21012 5982
rect 21036 5980 21092 5982
rect 21116 5980 21172 5982
rect 21196 5980 21252 5982
rect 20956 5928 20982 5980
rect 20982 5928 21012 5980
rect 21036 5928 21046 5980
rect 21046 5928 21092 5980
rect 21116 5928 21162 5980
rect 21162 5928 21172 5980
rect 21196 5928 21226 5980
rect 21226 5928 21252 5980
rect 20956 5926 21012 5928
rect 21036 5926 21092 5928
rect 21116 5926 21172 5928
rect 21196 5926 21252 5928
rect 13082 5722 13138 5778
rect 13634 5742 13690 5778
rect 13634 5722 13636 5742
rect 13636 5722 13688 5742
rect 13688 5722 13690 5742
rect 15956 5436 16012 5438
rect 16036 5436 16092 5438
rect 16116 5436 16172 5438
rect 16196 5436 16252 5438
rect 15956 5384 15982 5436
rect 15982 5384 16012 5436
rect 16036 5384 16046 5436
rect 16046 5384 16092 5436
rect 16116 5384 16162 5436
rect 16162 5384 16172 5436
rect 16196 5384 16226 5436
rect 16226 5384 16252 5436
rect 15956 5382 16012 5384
rect 16036 5382 16092 5384
rect 16116 5382 16172 5384
rect 16196 5382 16252 5384
rect 15566 5178 15622 5234
rect 20956 4892 21012 4894
rect 21036 4892 21092 4894
rect 21116 4892 21172 4894
rect 21196 4892 21252 4894
rect 20956 4840 20982 4892
rect 20982 4840 21012 4892
rect 21036 4840 21046 4892
rect 21046 4840 21092 4892
rect 21116 4840 21162 4892
rect 21162 4840 21172 4892
rect 21196 4840 21226 4892
rect 21226 4840 21252 4892
rect 20956 4838 21012 4840
rect 21036 4838 21092 4840
rect 21116 4838 21172 4840
rect 21196 4838 21252 4840
rect 20442 4654 20498 4690
rect 20442 4634 20444 4654
rect 20444 4634 20496 4654
rect 20496 4634 20498 4654
rect 15750 4518 15806 4554
rect 15750 4498 15752 4518
rect 15752 4498 15804 4518
rect 15804 4498 15806 4518
rect 15956 4348 16012 4350
rect 16036 4348 16092 4350
rect 16116 4348 16172 4350
rect 16196 4348 16252 4350
rect 15956 4296 15982 4348
rect 15982 4296 16012 4348
rect 16036 4296 16046 4348
rect 16046 4296 16092 4348
rect 16116 4296 16162 4348
rect 16162 4296 16172 4348
rect 16196 4296 16226 4348
rect 16226 4296 16252 4348
rect 15956 4294 16012 4296
rect 16036 4294 16092 4296
rect 16116 4294 16172 4296
rect 16196 4294 16252 4296
rect 20626 4518 20682 4554
rect 20626 4498 20628 4518
rect 20628 4498 20680 4518
rect 20680 4498 20682 4518
rect 12806 4090 12862 4146
rect 22926 13746 22982 13802
rect 22466 7626 22522 7682
rect 23938 18798 23994 18834
rect 23938 18778 23940 18798
rect 23940 18778 23992 18798
rect 23992 18778 23994 18798
rect 23938 18234 23994 18290
rect 23754 17826 23810 17882
rect 23478 12250 23534 12306
rect 23662 9394 23718 9450
rect 23938 17710 23994 17746
rect 23938 17690 23940 17710
rect 23940 17690 23992 17710
rect 23992 17690 23994 17710
rect 23938 13338 23994 13394
rect 24030 12386 24086 12442
rect 23938 9530 23994 9586
rect 23938 9006 23994 9042
rect 23938 8986 23940 9006
rect 23940 8986 23992 9006
rect 23992 8986 23994 9006
rect 23570 8306 23626 8362
rect 23478 7898 23534 7954
rect 23938 7510 23994 7546
rect 23938 7490 23940 7510
rect 23940 7490 23992 7510
rect 23992 7490 23994 7510
rect 24122 11570 24178 11626
rect 24122 10618 24178 10674
rect 24490 21226 24546 21282
rect 25042 22994 25098 23050
rect 24858 21498 24914 21554
rect 24858 20002 24914 20058
rect 24950 18778 25006 18834
rect 25502 19322 25558 19378
rect 24858 17826 24914 17882
rect 24766 17010 24822 17066
rect 24674 15378 24730 15434
rect 24306 11026 24362 11082
rect 24214 10346 24270 10402
rect 24122 9294 24124 9314
rect 24124 9294 24176 9314
rect 24176 9294 24178 9314
rect 24122 9258 24178 9294
rect 24122 8442 24178 8498
rect 24122 8054 24178 8090
rect 24122 8034 24124 8054
rect 24124 8034 24176 8054
rect 24176 8034 24178 8054
rect 24122 6694 24178 6730
rect 24122 6674 24124 6694
rect 24124 6674 24176 6694
rect 24176 6674 24178 6694
rect 24122 5042 24178 5098
rect 24306 5042 24362 5098
rect 24306 4090 24362 4146
rect 23938 3990 23940 4010
rect 23940 3990 23992 4010
rect 23992 3990 23994 4010
rect 23938 3954 23994 3990
rect 24122 3854 24124 3874
rect 24124 3854 24176 3874
rect 24176 3854 24178 3874
rect 24122 3818 24178 3854
rect 20956 3804 21012 3806
rect 21036 3804 21092 3806
rect 21116 3804 21172 3806
rect 21196 3804 21252 3806
rect 20956 3752 20982 3804
rect 20982 3752 21012 3804
rect 21036 3752 21046 3804
rect 21046 3752 21092 3804
rect 21116 3752 21162 3804
rect 21162 3752 21172 3804
rect 21196 3752 21226 3804
rect 21226 3752 21252 3804
rect 20956 3750 21012 3752
rect 21036 3750 21092 3752
rect 21116 3750 21172 3752
rect 21196 3750 21252 3752
rect 20718 3546 20774 3602
rect 24858 13338 24914 13394
rect 25226 17962 25282 18018
rect 25134 14562 25190 14618
rect 25042 13882 25098 13938
rect 24950 12386 25006 12442
rect 24950 12250 25006 12306
rect 24858 11842 24914 11898
rect 25956 21756 26012 21758
rect 26036 21756 26092 21758
rect 26116 21756 26172 21758
rect 26196 21756 26252 21758
rect 25956 21704 25982 21756
rect 25982 21704 26012 21756
rect 26036 21704 26046 21756
rect 26046 21704 26092 21756
rect 26116 21704 26162 21756
rect 26162 21704 26172 21756
rect 26196 21704 26226 21756
rect 26226 21704 26252 21756
rect 25956 21702 26012 21704
rect 26036 21702 26092 21704
rect 26116 21702 26172 21704
rect 26196 21702 26252 21704
rect 25956 20668 26012 20670
rect 26036 20668 26092 20670
rect 26116 20668 26172 20670
rect 26196 20668 26252 20670
rect 25956 20616 25982 20668
rect 25982 20616 26012 20668
rect 26036 20616 26046 20668
rect 26046 20616 26092 20668
rect 26116 20616 26162 20668
rect 26162 20616 26172 20668
rect 26196 20616 26226 20668
rect 26226 20616 26252 20668
rect 25956 20614 26012 20616
rect 26036 20614 26092 20616
rect 26116 20614 26172 20616
rect 26196 20614 26252 20616
rect 25956 19580 26012 19582
rect 26036 19580 26092 19582
rect 26116 19580 26172 19582
rect 26196 19580 26252 19582
rect 25956 19528 25982 19580
rect 25982 19528 26012 19580
rect 26036 19528 26046 19580
rect 26046 19528 26092 19580
rect 26116 19528 26162 19580
rect 26162 19528 26172 19580
rect 26196 19528 26226 19580
rect 26226 19528 26252 19580
rect 25956 19526 26012 19528
rect 26036 19526 26092 19528
rect 26116 19526 26172 19528
rect 26196 19526 26252 19528
rect 25870 19186 25926 19242
rect 25956 18492 26012 18494
rect 26036 18492 26092 18494
rect 26116 18492 26172 18494
rect 26196 18492 26252 18494
rect 25956 18440 25982 18492
rect 25982 18440 26012 18492
rect 26036 18440 26046 18492
rect 26046 18440 26092 18492
rect 26116 18440 26162 18492
rect 26162 18440 26172 18492
rect 26196 18440 26226 18492
rect 26226 18440 26252 18492
rect 25956 18438 26012 18440
rect 26036 18438 26092 18440
rect 26116 18438 26172 18440
rect 26196 18438 26252 18440
rect 25594 17554 25650 17610
rect 25502 13746 25558 13802
rect 25502 12794 25558 12850
rect 25134 11706 25190 11762
rect 25042 11162 25098 11218
rect 24950 10482 25006 10538
rect 24858 9938 24914 9994
rect 15956 3260 16012 3262
rect 16036 3260 16092 3262
rect 16116 3260 16172 3262
rect 16196 3260 16252 3262
rect 15956 3208 15982 3260
rect 15982 3208 16012 3260
rect 16036 3208 16046 3260
rect 16046 3208 16092 3260
rect 16116 3208 16162 3260
rect 16162 3208 16172 3260
rect 16196 3208 16226 3260
rect 16226 3208 16252 3260
rect 15956 3206 16012 3208
rect 16036 3206 16092 3208
rect 16116 3206 16172 3208
rect 16196 3206 16252 3208
rect 24122 3430 24178 3466
rect 24122 3410 24124 3430
rect 24124 3410 24176 3430
rect 24176 3410 24178 3430
rect 23938 3002 23994 3058
rect 20956 2716 21012 2718
rect 21036 2716 21092 2718
rect 21116 2716 21172 2718
rect 21196 2716 21252 2718
rect 20956 2664 20982 2716
rect 20982 2664 21012 2716
rect 21036 2664 21046 2716
rect 21046 2664 21092 2716
rect 21116 2664 21162 2716
rect 21162 2664 21172 2716
rect 21196 2664 21226 2716
rect 21226 2664 21252 2716
rect 20956 2662 21012 2664
rect 21036 2662 21092 2664
rect 21116 2662 21172 2664
rect 21196 2662 21252 2664
rect 24214 2614 24270 2650
rect 24214 2594 24216 2614
rect 24216 2594 24268 2614
rect 24268 2594 24270 2614
rect 15956 2172 16012 2174
rect 16036 2172 16092 2174
rect 16116 2172 16172 2174
rect 16196 2172 16252 2174
rect 15956 2120 15982 2172
rect 15982 2120 16012 2172
rect 16036 2120 16046 2172
rect 16046 2120 16092 2172
rect 16116 2120 16162 2172
rect 16162 2120 16172 2172
rect 16196 2120 16226 2172
rect 16226 2120 16252 2172
rect 15956 2118 16012 2120
rect 16036 2118 16092 2120
rect 16116 2118 16172 2120
rect 16196 2118 16252 2120
rect 12714 1914 12770 1970
rect 24030 1914 24086 1970
rect 12346 1642 12402 1698
rect 12530 1642 12586 1698
rect 25134 2478 25190 2514
rect 25134 2458 25136 2478
rect 25136 2458 25188 2478
rect 25188 2458 25190 2478
rect 25956 17404 26012 17406
rect 26036 17404 26092 17406
rect 26116 17404 26172 17406
rect 26196 17404 26252 17406
rect 25956 17352 25982 17404
rect 25982 17352 26012 17404
rect 26036 17352 26046 17404
rect 26046 17352 26092 17404
rect 26116 17352 26162 17404
rect 26162 17352 26172 17404
rect 26196 17352 26226 17404
rect 26226 17352 26252 17404
rect 25956 17350 26012 17352
rect 26036 17350 26092 17352
rect 26116 17350 26172 17352
rect 26196 17350 26252 17352
rect 25956 16316 26012 16318
rect 26036 16316 26092 16318
rect 26116 16316 26172 16318
rect 26196 16316 26252 16318
rect 25956 16264 25982 16316
rect 25982 16264 26012 16316
rect 26036 16264 26046 16316
rect 26046 16264 26092 16316
rect 26116 16264 26162 16316
rect 26162 16264 26172 16316
rect 26196 16264 26226 16316
rect 26226 16264 26252 16316
rect 25956 16262 26012 16264
rect 26036 16262 26092 16264
rect 26116 16262 26172 16264
rect 26196 16262 26252 16264
rect 25686 16058 25742 16114
rect 25594 5722 25650 5778
rect 25956 15228 26012 15230
rect 26036 15228 26092 15230
rect 26116 15228 26172 15230
rect 26196 15228 26252 15230
rect 25956 15176 25982 15228
rect 25982 15176 26012 15228
rect 26036 15176 26046 15228
rect 26046 15176 26092 15228
rect 26116 15176 26162 15228
rect 26162 15176 26172 15228
rect 26196 15176 26226 15228
rect 26226 15176 26252 15228
rect 25956 15174 26012 15176
rect 26036 15174 26092 15176
rect 26116 15174 26172 15176
rect 26196 15174 26252 15176
rect 25956 14140 26012 14142
rect 26036 14140 26092 14142
rect 26116 14140 26172 14142
rect 26196 14140 26252 14142
rect 25956 14088 25982 14140
rect 25982 14088 26012 14140
rect 26036 14088 26046 14140
rect 26046 14088 26092 14140
rect 26116 14088 26162 14140
rect 26162 14088 26172 14140
rect 26196 14088 26226 14140
rect 26226 14088 26252 14140
rect 25956 14086 26012 14088
rect 26036 14086 26092 14088
rect 26116 14086 26172 14088
rect 26196 14086 26252 14088
rect 25956 13052 26012 13054
rect 26036 13052 26092 13054
rect 26116 13052 26172 13054
rect 26196 13052 26252 13054
rect 25956 13000 25982 13052
rect 25982 13000 26012 13052
rect 26036 13000 26046 13052
rect 26046 13000 26092 13052
rect 26116 13000 26162 13052
rect 26162 13000 26172 13052
rect 26196 13000 26226 13052
rect 26226 13000 26252 13052
rect 25956 12998 26012 13000
rect 26036 12998 26092 13000
rect 26116 12998 26172 13000
rect 26196 12998 26252 13000
rect 25956 11964 26012 11966
rect 26036 11964 26092 11966
rect 26116 11964 26172 11966
rect 26196 11964 26252 11966
rect 25956 11912 25982 11964
rect 25982 11912 26012 11964
rect 26036 11912 26046 11964
rect 26046 11912 26092 11964
rect 26116 11912 26162 11964
rect 26162 11912 26172 11964
rect 26196 11912 26226 11964
rect 26226 11912 26252 11964
rect 25956 11910 26012 11912
rect 26036 11910 26092 11912
rect 26116 11910 26172 11912
rect 26196 11910 26252 11912
rect 25956 10876 26012 10878
rect 26036 10876 26092 10878
rect 26116 10876 26172 10878
rect 26196 10876 26252 10878
rect 25956 10824 25982 10876
rect 25982 10824 26012 10876
rect 26036 10824 26046 10876
rect 26046 10824 26092 10876
rect 26116 10824 26162 10876
rect 26162 10824 26172 10876
rect 26196 10824 26226 10876
rect 26226 10824 26252 10876
rect 25956 10822 26012 10824
rect 26036 10822 26092 10824
rect 26116 10822 26172 10824
rect 26196 10822 26252 10824
rect 25956 9788 26012 9790
rect 26036 9788 26092 9790
rect 26116 9788 26172 9790
rect 26196 9788 26252 9790
rect 25956 9736 25982 9788
rect 25982 9736 26012 9788
rect 26036 9736 26046 9788
rect 26046 9736 26092 9788
rect 26116 9736 26162 9788
rect 26162 9736 26172 9788
rect 26196 9736 26226 9788
rect 26226 9736 26252 9788
rect 25956 9734 26012 9736
rect 26036 9734 26092 9736
rect 26116 9734 26172 9736
rect 26196 9734 26252 9736
rect 25956 8700 26012 8702
rect 26036 8700 26092 8702
rect 26116 8700 26172 8702
rect 26196 8700 26252 8702
rect 25956 8648 25982 8700
rect 25982 8648 26012 8700
rect 26036 8648 26046 8700
rect 26046 8648 26092 8700
rect 26116 8648 26162 8700
rect 26162 8648 26172 8700
rect 26196 8648 26226 8700
rect 26226 8648 26252 8700
rect 25956 8646 26012 8648
rect 26036 8646 26092 8648
rect 26116 8646 26172 8648
rect 26196 8646 26252 8648
rect 25956 7612 26012 7614
rect 26036 7612 26092 7614
rect 26116 7612 26172 7614
rect 26196 7612 26252 7614
rect 25956 7560 25982 7612
rect 25982 7560 26012 7612
rect 26036 7560 26046 7612
rect 26046 7560 26092 7612
rect 26116 7560 26162 7612
rect 26162 7560 26172 7612
rect 26196 7560 26226 7612
rect 26226 7560 26252 7612
rect 25956 7558 26012 7560
rect 26036 7558 26092 7560
rect 26116 7558 26172 7560
rect 26196 7558 26252 7560
rect 25956 6524 26012 6526
rect 26036 6524 26092 6526
rect 26116 6524 26172 6526
rect 26196 6524 26252 6526
rect 25956 6472 25982 6524
rect 25982 6472 26012 6524
rect 26036 6472 26046 6524
rect 26046 6472 26092 6524
rect 26116 6472 26162 6524
rect 26162 6472 26172 6524
rect 26196 6472 26226 6524
rect 26226 6472 26252 6524
rect 25956 6470 26012 6472
rect 26036 6470 26092 6472
rect 26116 6470 26172 6472
rect 26196 6470 26252 6472
rect 25956 5436 26012 5438
rect 26036 5436 26092 5438
rect 26116 5436 26172 5438
rect 26196 5436 26252 5438
rect 25956 5384 25982 5436
rect 25982 5384 26012 5436
rect 26036 5384 26046 5436
rect 26046 5384 26092 5436
rect 26116 5384 26162 5436
rect 26162 5384 26172 5436
rect 26196 5384 26226 5436
rect 26226 5384 26252 5436
rect 25956 5382 26012 5384
rect 26036 5382 26092 5384
rect 26116 5382 26172 5384
rect 26196 5382 26252 5384
rect 25686 5178 25742 5234
rect 25956 4348 26012 4350
rect 26036 4348 26092 4350
rect 26116 4348 26172 4350
rect 26196 4348 26252 4350
rect 25956 4296 25982 4348
rect 25982 4296 26012 4348
rect 26036 4296 26046 4348
rect 26046 4296 26092 4348
rect 26116 4296 26162 4348
rect 26162 4296 26172 4348
rect 26196 4296 26226 4348
rect 26226 4296 26252 4348
rect 25956 4294 26012 4296
rect 26036 4294 26092 4296
rect 26116 4294 26172 4296
rect 26196 4294 26252 4296
rect 25956 3260 26012 3262
rect 26036 3260 26092 3262
rect 26116 3260 26172 3262
rect 26196 3260 26252 3262
rect 25956 3208 25982 3260
rect 25982 3208 26012 3260
rect 26036 3208 26046 3260
rect 26046 3208 26092 3260
rect 26116 3208 26162 3260
rect 26162 3208 26172 3260
rect 26196 3208 26226 3260
rect 26226 3208 26252 3260
rect 25956 3206 26012 3208
rect 26036 3206 26092 3208
rect 26116 3206 26172 3208
rect 26196 3206 26252 3208
rect 25502 2322 25558 2378
rect 24858 1506 24914 1562
rect 25956 2172 26012 2174
rect 26036 2172 26092 2174
rect 26116 2172 26172 2174
rect 26196 2172 26252 2174
rect 25956 2120 25982 2172
rect 25982 2120 26012 2172
rect 26036 2120 26046 2172
rect 26046 2120 26092 2172
rect 26116 2120 26162 2172
rect 26162 2120 26172 2172
rect 26196 2120 26226 2172
rect 26226 2120 26252 2172
rect 25956 2118 26012 2120
rect 26036 2118 26092 2120
rect 26116 2118 26172 2120
rect 26196 2118 26252 2120
rect 12346 282 12402 338
rect 12530 282 12586 338
rect 25318 282 25374 338
rect 9494 10 9550 66
<< metal3 >>
rect 0 23596 480 23626
rect 3877 23596 3943 23599
rect 0 23594 3943 23596
rect 0 23538 3882 23594
rect 3938 23538 3943 23594
rect 0 23536 3943 23538
rect 0 23506 480 23536
rect 3877 23533 3943 23536
rect 24761 23596 24827 23599
rect 29520 23596 30000 23626
rect 24761 23594 30000 23596
rect 24761 23538 24766 23594
rect 24822 23538 30000 23594
rect 24761 23536 30000 23538
rect 24761 23533 24827 23536
rect 29520 23506 30000 23536
rect 0 23052 480 23082
rect 3325 23052 3391 23055
rect 0 23050 3391 23052
rect 0 22994 3330 23050
rect 3386 22994 3391 23050
rect 0 22992 3391 22994
rect 0 22962 480 22992
rect 3325 22989 3391 22992
rect 25037 23052 25103 23055
rect 29520 23052 30000 23082
rect 25037 23050 30000 23052
rect 25037 22994 25042 23050
rect 25098 22994 30000 23050
rect 25037 22992 30000 22994
rect 25037 22989 25103 22992
rect 29520 22962 30000 22992
rect 0 22372 480 22402
rect 3509 22372 3575 22375
rect 0 22370 3575 22372
rect 0 22314 3514 22370
rect 3570 22314 3575 22370
rect 0 22312 3575 22314
rect 0 22282 480 22312
rect 3509 22309 3575 22312
rect 24393 22372 24459 22375
rect 29520 22372 30000 22402
rect 24393 22370 30000 22372
rect 24393 22314 24398 22370
rect 24454 22314 30000 22370
rect 24393 22312 30000 22314
rect 24393 22309 24459 22312
rect 29520 22282 30000 22312
rect 0 21828 480 21858
rect 3417 21828 3483 21831
rect 29520 21828 30000 21858
rect 0 21826 3483 21828
rect 0 21770 3422 21826
rect 3478 21770 3483 21826
rect 0 21768 3483 21770
rect 0 21738 480 21768
rect 3417 21765 3483 21768
rect 27846 21768 30000 21828
rect 5944 21762 6264 21763
rect 5944 21698 5952 21762
rect 6016 21698 6032 21762
rect 6096 21698 6112 21762
rect 6176 21698 6192 21762
rect 6256 21698 6264 21762
rect 5944 21697 6264 21698
rect 15944 21762 16264 21763
rect 15944 21698 15952 21762
rect 16016 21698 16032 21762
rect 16096 21698 16112 21762
rect 16176 21698 16192 21762
rect 16256 21698 16264 21762
rect 15944 21697 16264 21698
rect 25944 21762 26264 21763
rect 25944 21698 25952 21762
rect 26016 21698 26032 21762
rect 26096 21698 26112 21762
rect 26176 21698 26192 21762
rect 26256 21698 26264 21762
rect 25944 21697 26264 21698
rect 24853 21556 24919 21559
rect 27846 21556 27906 21768
rect 29520 21738 30000 21768
rect 24853 21554 27906 21556
rect 24853 21498 24858 21554
rect 24914 21498 27906 21554
rect 24853 21496 27906 21498
rect 24853 21493 24919 21496
rect 0 21284 480 21314
rect 3141 21284 3207 21287
rect 0 21282 3207 21284
rect 0 21226 3146 21282
rect 3202 21226 3207 21282
rect 0 21224 3207 21226
rect 0 21194 480 21224
rect 3141 21221 3207 21224
rect 24485 21284 24551 21287
rect 29520 21284 30000 21314
rect 24485 21282 30000 21284
rect 24485 21226 24490 21282
rect 24546 21226 30000 21282
rect 24485 21224 30000 21226
rect 24485 21221 24551 21224
rect 10944 21218 11264 21219
rect 10944 21154 10952 21218
rect 11016 21154 11032 21218
rect 11096 21154 11112 21218
rect 11176 21154 11192 21218
rect 11256 21154 11264 21218
rect 10944 21153 11264 21154
rect 20944 21218 21264 21219
rect 20944 21154 20952 21218
rect 21016 21154 21032 21218
rect 21096 21154 21112 21218
rect 21176 21154 21192 21218
rect 21256 21154 21264 21218
rect 29520 21194 30000 21224
rect 20944 21153 21264 21154
rect 5944 20674 6264 20675
rect 0 20604 480 20634
rect 5944 20610 5952 20674
rect 6016 20610 6032 20674
rect 6096 20610 6112 20674
rect 6176 20610 6192 20674
rect 6256 20610 6264 20674
rect 5944 20609 6264 20610
rect 15944 20674 16264 20675
rect 15944 20610 15952 20674
rect 16016 20610 16032 20674
rect 16096 20610 16112 20674
rect 16176 20610 16192 20674
rect 16256 20610 16264 20674
rect 15944 20609 16264 20610
rect 25944 20674 26264 20675
rect 25944 20610 25952 20674
rect 26016 20610 26032 20674
rect 26096 20610 26112 20674
rect 26176 20610 26192 20674
rect 26256 20610 26264 20674
rect 25944 20609 26264 20610
rect 3969 20604 4035 20607
rect 29520 20604 30000 20634
rect 0 20602 4035 20604
rect 0 20546 3974 20602
rect 4030 20546 4035 20602
rect 0 20544 4035 20546
rect 0 20514 480 20544
rect 3969 20541 4035 20544
rect 27846 20544 30000 20604
rect 24025 20468 24091 20471
rect 27846 20468 27906 20544
rect 29520 20514 30000 20544
rect 24025 20466 27906 20468
rect 24025 20410 24030 20466
rect 24086 20410 27906 20466
rect 24025 20408 27906 20410
rect 24025 20405 24091 20408
rect 10944 20130 11264 20131
rect 0 20060 480 20090
rect 10944 20066 10952 20130
rect 11016 20066 11032 20130
rect 11096 20066 11112 20130
rect 11176 20066 11192 20130
rect 11256 20066 11264 20130
rect 10944 20065 11264 20066
rect 20944 20130 21264 20131
rect 20944 20066 20952 20130
rect 21016 20066 21032 20130
rect 21096 20066 21112 20130
rect 21176 20066 21192 20130
rect 21256 20066 21264 20130
rect 20944 20065 21264 20066
rect 3601 20060 3667 20063
rect 0 20058 3667 20060
rect 0 20002 3606 20058
rect 3662 20002 3667 20058
rect 0 20000 3667 20002
rect 0 19970 480 20000
rect 3601 19997 3667 20000
rect 24853 20060 24919 20063
rect 29520 20060 30000 20090
rect 24853 20058 30000 20060
rect 24853 20002 24858 20058
rect 24914 20002 30000 20058
rect 24853 20000 30000 20002
rect 24853 19997 24919 20000
rect 29520 19970 30000 20000
rect 5944 19586 6264 19587
rect 5944 19522 5952 19586
rect 6016 19522 6032 19586
rect 6096 19522 6112 19586
rect 6176 19522 6192 19586
rect 6256 19522 6264 19586
rect 5944 19521 6264 19522
rect 15944 19586 16264 19587
rect 15944 19522 15952 19586
rect 16016 19522 16032 19586
rect 16096 19522 16112 19586
rect 16176 19522 16192 19586
rect 16256 19522 16264 19586
rect 15944 19521 16264 19522
rect 25944 19586 26264 19587
rect 25944 19522 25952 19586
rect 26016 19522 26032 19586
rect 26096 19522 26112 19586
rect 26176 19522 26192 19586
rect 26256 19522 26264 19586
rect 25944 19521 26264 19522
rect 0 19380 480 19410
rect 3785 19380 3851 19383
rect 0 19378 3851 19380
rect 0 19322 3790 19378
rect 3846 19322 3851 19378
rect 0 19320 3851 19322
rect 0 19290 480 19320
rect 3785 19317 3851 19320
rect 8845 19380 8911 19383
rect 11329 19380 11395 19383
rect 8845 19378 11395 19380
rect 8845 19322 8850 19378
rect 8906 19322 11334 19378
rect 11390 19322 11395 19378
rect 8845 19320 11395 19322
rect 8845 19317 8911 19320
rect 11329 19317 11395 19320
rect 25497 19380 25563 19383
rect 29520 19380 30000 19410
rect 25497 19378 30000 19380
rect 25497 19322 25502 19378
rect 25558 19322 30000 19378
rect 25497 19320 30000 19322
rect 25497 19317 25563 19320
rect 29520 19290 30000 19320
rect 20805 19244 20871 19247
rect 25865 19244 25931 19247
rect 20805 19242 25931 19244
rect 20805 19186 20810 19242
rect 20866 19186 25870 19242
rect 25926 19186 25931 19242
rect 20805 19184 25931 19186
rect 20805 19181 20871 19184
rect 25865 19181 25931 19184
rect 10944 19042 11264 19043
rect 10944 18978 10952 19042
rect 11016 18978 11032 19042
rect 11096 18978 11112 19042
rect 11176 18978 11192 19042
rect 11256 18978 11264 19042
rect 10944 18977 11264 18978
rect 20944 19042 21264 19043
rect 20944 18978 20952 19042
rect 21016 18978 21032 19042
rect 21096 18978 21112 19042
rect 21176 18978 21192 19042
rect 21256 18978 21264 19042
rect 20944 18977 21264 18978
rect 3693 18972 3759 18975
rect 7005 18972 7071 18975
rect 8569 18972 8635 18975
rect 3693 18970 8635 18972
rect 3693 18914 3698 18970
rect 3754 18914 7010 18970
rect 7066 18914 8574 18970
rect 8630 18914 8635 18970
rect 3693 18912 8635 18914
rect 3693 18909 3759 18912
rect 7005 18909 7071 18912
rect 8569 18909 8635 18912
rect 16757 18972 16823 18975
rect 18689 18972 18755 18975
rect 16757 18970 18755 18972
rect 16757 18914 16762 18970
rect 16818 18914 18694 18970
rect 18750 18914 18755 18970
rect 16757 18912 18755 18914
rect 16757 18909 16823 18912
rect 18689 18909 18755 18912
rect 0 18836 480 18866
rect 3233 18836 3299 18839
rect 0 18834 3299 18836
rect 0 18778 3238 18834
rect 3294 18778 3299 18834
rect 0 18776 3299 18778
rect 0 18746 480 18776
rect 3233 18773 3299 18776
rect 3877 18836 3943 18839
rect 23933 18836 23999 18839
rect 3877 18834 23999 18836
rect 3877 18778 3882 18834
rect 3938 18778 23938 18834
rect 23994 18778 23999 18834
rect 3877 18776 23999 18778
rect 3877 18773 3943 18776
rect 23933 18773 23999 18776
rect 24945 18836 25011 18839
rect 29520 18836 30000 18866
rect 24945 18834 30000 18836
rect 24945 18778 24950 18834
rect 25006 18778 30000 18834
rect 24945 18776 30000 18778
rect 24945 18773 25011 18776
rect 29520 18746 30000 18776
rect 5944 18498 6264 18499
rect 5944 18434 5952 18498
rect 6016 18434 6032 18498
rect 6096 18434 6112 18498
rect 6176 18434 6192 18498
rect 6256 18434 6264 18498
rect 5944 18433 6264 18434
rect 15944 18498 16264 18499
rect 15944 18434 15952 18498
rect 16016 18434 16032 18498
rect 16096 18434 16112 18498
rect 16176 18434 16192 18498
rect 16256 18434 16264 18498
rect 15944 18433 16264 18434
rect 25944 18498 26264 18499
rect 25944 18434 25952 18498
rect 26016 18434 26032 18498
rect 26096 18434 26112 18498
rect 26176 18434 26192 18498
rect 26256 18434 26264 18498
rect 25944 18433 26264 18434
rect 19885 18428 19951 18431
rect 19885 18426 24226 18428
rect 19885 18370 19890 18426
rect 19946 18370 24226 18426
rect 19885 18368 24226 18370
rect 19885 18365 19951 18368
rect 0 18292 480 18322
rect 2865 18292 2931 18295
rect 0 18290 2931 18292
rect 0 18234 2870 18290
rect 2926 18234 2931 18290
rect 0 18232 2931 18234
rect 0 18202 480 18232
rect 2865 18229 2931 18232
rect 3325 18292 3391 18295
rect 23933 18292 23999 18295
rect 3325 18290 23999 18292
rect 3325 18234 3330 18290
rect 3386 18234 23938 18290
rect 23994 18234 23999 18290
rect 3325 18232 23999 18234
rect 24166 18292 24226 18368
rect 29520 18292 30000 18322
rect 24166 18232 30000 18292
rect 3325 18229 3391 18232
rect 23933 18229 23999 18232
rect 29520 18202 30000 18232
rect 8569 18156 8635 18159
rect 13077 18156 13143 18159
rect 15377 18156 15443 18159
rect 8569 18154 15443 18156
rect 8569 18098 8574 18154
rect 8630 18098 13082 18154
rect 13138 18098 15382 18154
rect 15438 18098 15443 18154
rect 8569 18096 15443 18098
rect 8569 18093 8635 18096
rect 13077 18093 13143 18096
rect 15377 18093 15443 18096
rect 24894 17958 24900 18022
rect 24964 18020 24970 18022
rect 25221 18020 25287 18023
rect 24964 18018 25287 18020
rect 24964 17962 25226 18018
rect 25282 17962 25287 18018
rect 24964 17960 25287 17962
rect 24964 17958 24970 17960
rect 25221 17957 25287 17960
rect 10944 17954 11264 17955
rect 10944 17890 10952 17954
rect 11016 17890 11032 17954
rect 11096 17890 11112 17954
rect 11176 17890 11192 17954
rect 11256 17890 11264 17954
rect 10944 17889 11264 17890
rect 20944 17954 21264 17955
rect 20944 17890 20952 17954
rect 21016 17890 21032 17954
rect 21096 17890 21112 17954
rect 21176 17890 21192 17954
rect 21256 17890 21264 17954
rect 20944 17889 21264 17890
rect 23749 17884 23815 17887
rect 24853 17884 24919 17887
rect 23749 17882 24919 17884
rect 23749 17826 23754 17882
rect 23810 17826 24858 17882
rect 24914 17826 24919 17882
rect 23749 17824 24919 17826
rect 23749 17821 23815 17824
rect 24853 17821 24919 17824
rect 3509 17748 3575 17751
rect 23933 17748 23999 17751
rect 3509 17746 23999 17748
rect 3509 17690 3514 17746
rect 3570 17690 23938 17746
rect 23994 17690 23999 17746
rect 3509 17688 23999 17690
rect 3509 17685 3575 17688
rect 23933 17685 23999 17688
rect 0 17612 480 17642
rect 3325 17612 3391 17615
rect 0 17610 3391 17612
rect 0 17554 3330 17610
rect 3386 17554 3391 17610
rect 0 17552 3391 17554
rect 0 17522 480 17552
rect 3325 17549 3391 17552
rect 25589 17612 25655 17615
rect 29520 17612 30000 17642
rect 25589 17610 30000 17612
rect 25589 17554 25594 17610
rect 25650 17554 30000 17610
rect 25589 17552 30000 17554
rect 25589 17549 25655 17552
rect 29520 17522 30000 17552
rect 5944 17410 6264 17411
rect 5944 17346 5952 17410
rect 6016 17346 6032 17410
rect 6096 17346 6112 17410
rect 6176 17346 6192 17410
rect 6256 17346 6264 17410
rect 5944 17345 6264 17346
rect 15944 17410 16264 17411
rect 15944 17346 15952 17410
rect 16016 17346 16032 17410
rect 16096 17346 16112 17410
rect 16176 17346 16192 17410
rect 16256 17346 16264 17410
rect 15944 17345 16264 17346
rect 25944 17410 26264 17411
rect 25944 17346 25952 17410
rect 26016 17346 26032 17410
rect 26096 17346 26112 17410
rect 26176 17346 26192 17410
rect 26256 17346 26264 17410
rect 25944 17345 26264 17346
rect 0 17068 480 17098
rect 3509 17068 3575 17071
rect 0 17066 3575 17068
rect 0 17010 3514 17066
rect 3570 17010 3575 17066
rect 0 17008 3575 17010
rect 0 16978 480 17008
rect 3509 17005 3575 17008
rect 24761 17068 24827 17071
rect 29520 17068 30000 17098
rect 24761 17066 30000 17068
rect 24761 17010 24766 17066
rect 24822 17010 30000 17066
rect 24761 17008 30000 17010
rect 24761 17005 24827 17008
rect 29520 16978 30000 17008
rect 13537 16932 13603 16935
rect 17493 16932 17559 16935
rect 13537 16930 17559 16932
rect 13537 16874 13542 16930
rect 13598 16874 17498 16930
rect 17554 16874 17559 16930
rect 13537 16872 17559 16874
rect 13537 16869 13603 16872
rect 17493 16869 17559 16872
rect 10944 16866 11264 16867
rect 10944 16802 10952 16866
rect 11016 16802 11032 16866
rect 11096 16802 11112 16866
rect 11176 16802 11192 16866
rect 11256 16802 11264 16866
rect 10944 16801 11264 16802
rect 20944 16866 21264 16867
rect 20944 16802 20952 16866
rect 21016 16802 21032 16866
rect 21096 16802 21112 16866
rect 21176 16802 21192 16866
rect 21256 16802 21264 16866
rect 20944 16801 21264 16802
rect 0 16388 480 16418
rect 4061 16388 4127 16391
rect 29520 16388 30000 16418
rect 0 16386 4127 16388
rect 0 16330 4066 16386
rect 4122 16330 4127 16386
rect 0 16328 4127 16330
rect 0 16298 480 16328
rect 4061 16325 4127 16328
rect 27846 16328 30000 16388
rect 5944 16322 6264 16323
rect 5944 16258 5952 16322
rect 6016 16258 6032 16322
rect 6096 16258 6112 16322
rect 6176 16258 6192 16322
rect 6256 16258 6264 16322
rect 5944 16257 6264 16258
rect 15944 16322 16264 16323
rect 15944 16258 15952 16322
rect 16016 16258 16032 16322
rect 16096 16258 16112 16322
rect 16176 16258 16192 16322
rect 16256 16258 16264 16322
rect 15944 16257 16264 16258
rect 25944 16322 26264 16323
rect 25944 16258 25952 16322
rect 26016 16258 26032 16322
rect 26096 16258 26112 16322
rect 26176 16258 26192 16322
rect 26256 16258 26264 16322
rect 25944 16257 26264 16258
rect 25681 16116 25747 16119
rect 27846 16116 27906 16328
rect 29520 16298 30000 16328
rect 25681 16114 27906 16116
rect 25681 16058 25686 16114
rect 25742 16058 27906 16114
rect 25681 16056 27906 16058
rect 25681 16053 25747 16056
rect 7189 15980 7255 15983
rect 9949 15980 10015 15983
rect 7189 15978 10015 15980
rect 7189 15922 7194 15978
rect 7250 15922 9954 15978
rect 10010 15922 10015 15978
rect 7189 15920 10015 15922
rect 7189 15917 7255 15920
rect 9949 15917 10015 15920
rect 0 15844 480 15874
rect 3049 15844 3115 15847
rect 0 15842 3115 15844
rect 0 15786 3054 15842
rect 3110 15786 3115 15842
rect 0 15784 3115 15786
rect 0 15754 480 15784
rect 3049 15781 3115 15784
rect 21449 15844 21515 15847
rect 29520 15844 30000 15874
rect 21449 15842 30000 15844
rect 21449 15786 21454 15842
rect 21510 15786 30000 15842
rect 21449 15784 30000 15786
rect 21449 15781 21515 15784
rect 10944 15778 11264 15779
rect 10944 15714 10952 15778
rect 11016 15714 11032 15778
rect 11096 15714 11112 15778
rect 11176 15714 11192 15778
rect 11256 15714 11264 15778
rect 10944 15713 11264 15714
rect 20944 15778 21264 15779
rect 20944 15714 20952 15778
rect 21016 15714 21032 15778
rect 21096 15714 21112 15778
rect 21176 15714 21192 15778
rect 21256 15714 21264 15778
rect 29520 15754 30000 15784
rect 20944 15713 21264 15714
rect 24669 15436 24735 15439
rect 24669 15434 27906 15436
rect 24669 15378 24674 15434
rect 24730 15378 27906 15434
rect 24669 15376 27906 15378
rect 24669 15373 24735 15376
rect 0 15300 480 15330
rect 1393 15300 1459 15303
rect 0 15298 1459 15300
rect 0 15242 1398 15298
rect 1454 15242 1459 15298
rect 0 15240 1459 15242
rect 27846 15300 27906 15376
rect 29520 15300 30000 15330
rect 27846 15240 30000 15300
rect 0 15210 480 15240
rect 1393 15237 1459 15240
rect 5944 15234 6264 15235
rect 5944 15170 5952 15234
rect 6016 15170 6032 15234
rect 6096 15170 6112 15234
rect 6176 15170 6192 15234
rect 6256 15170 6264 15234
rect 5944 15169 6264 15170
rect 15944 15234 16264 15235
rect 15944 15170 15952 15234
rect 16016 15170 16032 15234
rect 16096 15170 16112 15234
rect 16176 15170 16192 15234
rect 16256 15170 16264 15234
rect 15944 15169 16264 15170
rect 25944 15234 26264 15235
rect 25944 15170 25952 15234
rect 26016 15170 26032 15234
rect 26096 15170 26112 15234
rect 26176 15170 26192 15234
rect 26256 15170 26264 15234
rect 29520 15210 30000 15240
rect 25944 15169 26264 15170
rect 8477 15164 8543 15167
rect 13445 15164 13511 15167
rect 8477 15162 13511 15164
rect 8477 15106 8482 15162
rect 8538 15106 13450 15162
rect 13506 15106 13511 15162
rect 8477 15104 13511 15106
rect 8477 15101 8543 15104
rect 13445 15101 13511 15104
rect 14089 15028 14155 15031
rect 18781 15028 18847 15031
rect 14089 15026 18847 15028
rect 14089 14970 14094 15026
rect 14150 14970 18786 15026
rect 18842 14970 18847 15026
rect 14089 14968 18847 14970
rect 14089 14965 14155 14968
rect 18781 14965 18847 14968
rect 10944 14690 11264 14691
rect 0 14620 480 14650
rect 10944 14626 10952 14690
rect 11016 14626 11032 14690
rect 11096 14626 11112 14690
rect 11176 14626 11192 14690
rect 11256 14626 11264 14690
rect 10944 14625 11264 14626
rect 20944 14690 21264 14691
rect 20944 14626 20952 14690
rect 21016 14626 21032 14690
rect 21096 14626 21112 14690
rect 21176 14626 21192 14690
rect 21256 14626 21264 14690
rect 20944 14625 21264 14626
rect 3417 14620 3483 14623
rect 0 14618 3483 14620
rect 0 14562 3422 14618
rect 3478 14562 3483 14618
rect 0 14560 3483 14562
rect 0 14530 480 14560
rect 3417 14557 3483 14560
rect 25129 14620 25195 14623
rect 29520 14620 30000 14650
rect 25129 14618 30000 14620
rect 25129 14562 25134 14618
rect 25190 14562 30000 14618
rect 25129 14560 30000 14562
rect 25129 14557 25195 14560
rect 29520 14530 30000 14560
rect 13445 14484 13511 14487
rect 19977 14484 20043 14487
rect 13445 14482 20043 14484
rect 13445 14426 13450 14482
rect 13506 14426 19982 14482
rect 20038 14426 20043 14482
rect 13445 14424 20043 14426
rect 13445 14421 13511 14424
rect 19977 14421 20043 14424
rect 5944 14146 6264 14147
rect 0 14076 480 14106
rect 5944 14082 5952 14146
rect 6016 14082 6032 14146
rect 6096 14082 6112 14146
rect 6176 14082 6192 14146
rect 6256 14082 6264 14146
rect 5944 14081 6264 14082
rect 15944 14146 16264 14147
rect 15944 14082 15952 14146
rect 16016 14082 16032 14146
rect 16096 14082 16112 14146
rect 16176 14082 16192 14146
rect 16256 14082 16264 14146
rect 15944 14081 16264 14082
rect 25944 14146 26264 14147
rect 25944 14082 25952 14146
rect 26016 14082 26032 14146
rect 26096 14082 26112 14146
rect 26176 14082 26192 14146
rect 26256 14082 26264 14146
rect 25944 14081 26264 14082
rect 1577 14076 1643 14079
rect 29520 14076 30000 14106
rect 0 14074 1643 14076
rect 0 14018 1582 14074
rect 1638 14018 1643 14074
rect 0 14016 1643 14018
rect 0 13986 480 14016
rect 1577 14013 1643 14016
rect 27846 14016 30000 14076
rect 25037 13940 25103 13943
rect 27846 13940 27906 14016
rect 29520 13986 30000 14016
rect 25037 13938 27906 13940
rect 25037 13882 25042 13938
rect 25098 13882 27906 13938
rect 25037 13880 27906 13882
rect 25037 13877 25103 13880
rect 22921 13804 22987 13807
rect 25497 13804 25563 13807
rect 22921 13802 25563 13804
rect 22921 13746 22926 13802
rect 22982 13746 25502 13802
rect 25558 13746 25563 13802
rect 22921 13744 25563 13746
rect 22921 13741 22987 13744
rect 25497 13741 25563 13744
rect 10944 13602 11264 13603
rect 10944 13538 10952 13602
rect 11016 13538 11032 13602
rect 11096 13538 11112 13602
rect 11176 13538 11192 13602
rect 11256 13538 11264 13602
rect 10944 13537 11264 13538
rect 20944 13602 21264 13603
rect 20944 13538 20952 13602
rect 21016 13538 21032 13602
rect 21096 13538 21112 13602
rect 21176 13538 21192 13602
rect 21256 13538 21264 13602
rect 20944 13537 21264 13538
rect 19517 13532 19583 13535
rect 19517 13530 20730 13532
rect 19517 13474 19522 13530
rect 19578 13474 20730 13530
rect 19517 13472 20730 13474
rect 19517 13469 19583 13472
rect 0 13396 480 13426
rect 1485 13396 1551 13399
rect 19701 13396 19767 13399
rect 0 13336 1410 13396
rect 0 13306 480 13336
rect 1350 13260 1410 13336
rect 1485 13394 19767 13396
rect 1485 13338 1490 13394
rect 1546 13338 19706 13394
rect 19762 13338 19767 13394
rect 1485 13336 19767 13338
rect 20670 13396 20730 13472
rect 23933 13396 23999 13399
rect 20670 13394 23999 13396
rect 20670 13338 23938 13394
rect 23994 13338 23999 13394
rect 20670 13336 23999 13338
rect 1485 13333 1551 13336
rect 19701 13333 19767 13336
rect 23933 13333 23999 13336
rect 24853 13396 24919 13399
rect 29520 13396 30000 13426
rect 24853 13394 30000 13396
rect 24853 13338 24858 13394
rect 24914 13338 30000 13394
rect 24853 13336 30000 13338
rect 24853 13333 24919 13336
rect 29520 13306 30000 13336
rect 3233 13260 3299 13263
rect 1350 13258 3299 13260
rect 1350 13202 3238 13258
rect 3294 13202 3299 13258
rect 1350 13200 3299 13202
rect 3233 13197 3299 13200
rect 3417 13260 3483 13263
rect 11973 13260 12039 13263
rect 3417 13258 12039 13260
rect 3417 13202 3422 13258
rect 3478 13202 11978 13258
rect 12034 13202 12039 13258
rect 3417 13200 12039 13202
rect 3417 13197 3483 13200
rect 11973 13197 12039 13200
rect 5944 13058 6264 13059
rect 5944 12994 5952 13058
rect 6016 12994 6032 13058
rect 6096 12994 6112 13058
rect 6176 12994 6192 13058
rect 6256 12994 6264 13058
rect 5944 12993 6264 12994
rect 15944 13058 16264 13059
rect 15944 12994 15952 13058
rect 16016 12994 16032 13058
rect 16096 12994 16112 13058
rect 16176 12994 16192 13058
rect 16256 12994 16264 13058
rect 15944 12993 16264 12994
rect 25944 13058 26264 13059
rect 25944 12994 25952 13058
rect 26016 12994 26032 13058
rect 26096 12994 26112 13058
rect 26176 12994 26192 13058
rect 26256 12994 26264 13058
rect 25944 12993 26264 12994
rect 0 12852 480 12882
rect 2773 12852 2839 12855
rect 0 12850 2839 12852
rect 0 12794 2778 12850
rect 2834 12794 2839 12850
rect 0 12792 2839 12794
rect 0 12762 480 12792
rect 2773 12789 2839 12792
rect 25497 12852 25563 12855
rect 29520 12852 30000 12882
rect 25497 12850 30000 12852
rect 25497 12794 25502 12850
rect 25558 12794 30000 12850
rect 25497 12792 30000 12794
rect 25497 12789 25563 12792
rect 29520 12762 30000 12792
rect 2221 12716 2287 12719
rect 19149 12716 19215 12719
rect 2221 12714 19215 12716
rect 2221 12658 2226 12714
rect 2282 12658 19154 12714
rect 19210 12658 19215 12714
rect 2221 12656 19215 12658
rect 2221 12653 2287 12656
rect 19149 12653 19215 12656
rect 10944 12514 11264 12515
rect 10944 12450 10952 12514
rect 11016 12450 11032 12514
rect 11096 12450 11112 12514
rect 11176 12450 11192 12514
rect 11256 12450 11264 12514
rect 10944 12449 11264 12450
rect 20944 12514 21264 12515
rect 20944 12450 20952 12514
rect 21016 12450 21032 12514
rect 21096 12450 21112 12514
rect 21176 12450 21192 12514
rect 21256 12450 21264 12514
rect 20944 12449 21264 12450
rect 24025 12444 24091 12447
rect 24945 12444 25011 12447
rect 24025 12442 25011 12444
rect 24025 12386 24030 12442
rect 24086 12386 24950 12442
rect 25006 12386 25011 12442
rect 24025 12384 25011 12386
rect 24025 12381 24091 12384
rect 24945 12381 25011 12384
rect 0 12308 480 12338
rect 3141 12308 3207 12311
rect 0 12306 3207 12308
rect 0 12250 3146 12306
rect 3202 12250 3207 12306
rect 0 12248 3207 12250
rect 0 12218 480 12248
rect 3141 12245 3207 12248
rect 3325 12308 3391 12311
rect 23473 12308 23539 12311
rect 3325 12306 23539 12308
rect 3325 12250 3330 12306
rect 3386 12250 23478 12306
rect 23534 12250 23539 12306
rect 3325 12248 23539 12250
rect 3325 12245 3391 12248
rect 23473 12245 23539 12248
rect 24945 12308 25011 12311
rect 29520 12308 30000 12338
rect 24945 12306 30000 12308
rect 24945 12250 24950 12306
rect 25006 12250 30000 12306
rect 24945 12248 30000 12250
rect 24945 12245 25011 12248
rect 29520 12218 30000 12248
rect 3233 12172 3299 12175
rect 7373 12172 7439 12175
rect 3233 12170 7439 12172
rect 3233 12114 3238 12170
rect 3294 12114 7378 12170
rect 7434 12114 7439 12170
rect 3233 12112 7439 12114
rect 3233 12109 3299 12112
rect 7373 12109 7439 12112
rect 7925 12172 7991 12175
rect 13905 12172 13971 12175
rect 7925 12170 13971 12172
rect 7925 12114 7930 12170
rect 7986 12114 13910 12170
rect 13966 12114 13971 12170
rect 7925 12112 13971 12114
rect 7925 12109 7991 12112
rect 13905 12109 13971 12112
rect 5944 11970 6264 11971
rect 5944 11906 5952 11970
rect 6016 11906 6032 11970
rect 6096 11906 6112 11970
rect 6176 11906 6192 11970
rect 6256 11906 6264 11970
rect 5944 11905 6264 11906
rect 15944 11970 16264 11971
rect 15944 11906 15952 11970
rect 16016 11906 16032 11970
rect 16096 11906 16112 11970
rect 16176 11906 16192 11970
rect 16256 11906 16264 11970
rect 15944 11905 16264 11906
rect 25944 11970 26264 11971
rect 25944 11906 25952 11970
rect 26016 11906 26032 11970
rect 26096 11906 26112 11970
rect 26176 11906 26192 11970
rect 26256 11906 26264 11970
rect 25944 11905 26264 11906
rect 13077 11900 13143 11903
rect 14733 11900 14799 11903
rect 24853 11900 24919 11903
rect 7974 11898 14799 11900
rect 7974 11842 13082 11898
rect 13138 11842 14738 11898
rect 14794 11842 14799 11898
rect 7974 11840 14799 11842
rect 2865 11764 2931 11767
rect 7974 11764 8034 11840
rect 13077 11837 13143 11840
rect 14733 11837 14799 11840
rect 16438 11898 24919 11900
rect 16438 11842 24858 11898
rect 24914 11842 24919 11898
rect 16438 11840 24919 11842
rect 2865 11762 8034 11764
rect 2865 11706 2870 11762
rect 2926 11706 8034 11762
rect 2865 11704 8034 11706
rect 8109 11764 8175 11767
rect 16438 11764 16498 11840
rect 24853 11837 24919 11840
rect 25129 11764 25195 11767
rect 8109 11762 16498 11764
rect 8109 11706 8114 11762
rect 8170 11706 16498 11762
rect 8109 11704 16498 11706
rect 21406 11762 25195 11764
rect 21406 11706 25134 11762
rect 25190 11706 25195 11762
rect 21406 11704 25195 11706
rect 2865 11701 2931 11704
rect 8109 11701 8175 11704
rect 0 11628 480 11658
rect 3325 11628 3391 11631
rect 12157 11628 12223 11631
rect 21406 11628 21466 11704
rect 25129 11701 25195 11704
rect 0 11626 3391 11628
rect 0 11570 3330 11626
rect 3386 11570 3391 11626
rect 0 11568 3391 11570
rect 0 11538 480 11568
rect 3325 11565 3391 11568
rect 3558 11626 21466 11628
rect 3558 11570 12162 11626
rect 12218 11570 21466 11626
rect 3558 11568 21466 11570
rect 24117 11628 24183 11631
rect 29520 11628 30000 11658
rect 24117 11626 30000 11628
rect 24117 11570 24122 11626
rect 24178 11570 30000 11626
rect 24117 11568 30000 11570
rect 2405 11492 2471 11495
rect 3558 11492 3618 11568
rect 12157 11565 12223 11568
rect 24117 11565 24183 11568
rect 29520 11538 30000 11568
rect 2405 11490 3618 11492
rect 2405 11434 2410 11490
rect 2466 11434 3618 11490
rect 2405 11432 3618 11434
rect 2405 11429 2471 11432
rect 10944 11426 11264 11427
rect 10944 11362 10952 11426
rect 11016 11362 11032 11426
rect 11096 11362 11112 11426
rect 11176 11362 11192 11426
rect 11256 11362 11264 11426
rect 10944 11361 11264 11362
rect 20944 11426 21264 11427
rect 20944 11362 20952 11426
rect 21016 11362 21032 11426
rect 21096 11362 21112 11426
rect 21176 11362 21192 11426
rect 21256 11362 21264 11426
rect 20944 11361 21264 11362
rect 2497 11356 2563 11359
rect 7097 11356 7163 11359
rect 8109 11356 8175 11359
rect 2497 11354 8175 11356
rect 2497 11298 2502 11354
rect 2558 11298 7102 11354
rect 7158 11298 8114 11354
rect 8170 11298 8175 11354
rect 2497 11296 8175 11298
rect 2497 11293 2563 11296
rect 7097 11293 7163 11296
rect 8109 11293 8175 11296
rect 2037 11220 2103 11223
rect 25037 11220 25103 11223
rect 2037 11218 25103 11220
rect 2037 11162 2042 11218
rect 2098 11162 25042 11218
rect 25098 11162 25103 11218
rect 2037 11160 25103 11162
rect 2037 11157 2103 11160
rect 25037 11157 25103 11160
rect 0 11084 480 11114
rect 3366 11084 3372 11086
rect 0 11024 3372 11084
rect 0 10994 480 11024
rect 3366 11022 3372 11024
rect 3436 11022 3442 11086
rect 8293 11084 8359 11087
rect 12065 11084 12131 11087
rect 8293 11082 12131 11084
rect 8293 11026 8298 11082
rect 8354 11026 12070 11082
rect 12126 11026 12131 11082
rect 8293 11024 12131 11026
rect 8293 11021 8359 11024
rect 12065 11021 12131 11024
rect 24301 11084 24367 11087
rect 29520 11084 30000 11114
rect 24301 11082 30000 11084
rect 24301 11026 24306 11082
rect 24362 11026 30000 11082
rect 24301 11024 30000 11026
rect 24301 11021 24367 11024
rect 29520 10994 30000 11024
rect 5944 10882 6264 10883
rect 5944 10818 5952 10882
rect 6016 10818 6032 10882
rect 6096 10818 6112 10882
rect 6176 10818 6192 10882
rect 6256 10818 6264 10882
rect 5944 10817 6264 10818
rect 15944 10882 16264 10883
rect 15944 10818 15952 10882
rect 16016 10818 16032 10882
rect 16096 10818 16112 10882
rect 16176 10818 16192 10882
rect 16256 10818 16264 10882
rect 15944 10817 16264 10818
rect 25944 10882 26264 10883
rect 25944 10818 25952 10882
rect 26016 10818 26032 10882
rect 26096 10818 26112 10882
rect 26176 10818 26192 10882
rect 26256 10818 26264 10882
rect 25944 10817 26264 10818
rect 24117 10676 24183 10679
rect 3374 10674 24183 10676
rect 3374 10618 24122 10674
rect 24178 10618 24183 10674
rect 3374 10616 24183 10618
rect 0 10404 480 10434
rect 3374 10404 3434 10616
rect 24117 10613 24183 10616
rect 8293 10540 8359 10543
rect 24945 10540 25011 10543
rect 8293 10538 25011 10540
rect 8293 10482 8298 10538
rect 8354 10482 24950 10538
rect 25006 10482 25011 10538
rect 8293 10480 25011 10482
rect 8293 10477 8359 10480
rect 24945 10477 25011 10480
rect 0 10344 3434 10404
rect 24209 10404 24275 10407
rect 29520 10404 30000 10434
rect 24209 10402 30000 10404
rect 24209 10346 24214 10402
rect 24270 10346 30000 10402
rect 24209 10344 30000 10346
rect 0 10314 480 10344
rect 24209 10341 24275 10344
rect 10944 10338 11264 10339
rect 10944 10274 10952 10338
rect 11016 10274 11032 10338
rect 11096 10274 11112 10338
rect 11176 10274 11192 10338
rect 11256 10274 11264 10338
rect 10944 10273 11264 10274
rect 20944 10338 21264 10339
rect 20944 10274 20952 10338
rect 21016 10274 21032 10338
rect 21096 10274 21112 10338
rect 21176 10274 21192 10338
rect 21256 10274 21264 10338
rect 29520 10314 30000 10344
rect 20944 10273 21264 10274
rect 3141 10268 3207 10271
rect 7833 10268 7899 10271
rect 3141 10266 7899 10268
rect 3141 10210 3146 10266
rect 3202 10210 7838 10266
rect 7894 10210 7899 10266
rect 3141 10208 7899 10210
rect 3141 10205 3207 10208
rect 7833 10205 7899 10208
rect 1393 9996 1459 9999
rect 8293 9996 8359 9999
rect 1393 9994 8359 9996
rect 1393 9938 1398 9994
rect 1454 9938 8298 9994
rect 8354 9938 8359 9994
rect 1393 9936 8359 9938
rect 1393 9933 1459 9936
rect 8293 9933 8359 9936
rect 24853 9996 24919 9999
rect 24853 9994 27906 9996
rect 24853 9938 24858 9994
rect 24914 9938 27906 9994
rect 24853 9936 27906 9938
rect 24853 9933 24919 9936
rect 0 9860 480 9890
rect 1577 9860 1643 9863
rect 0 9858 1643 9860
rect 0 9802 1582 9858
rect 1638 9802 1643 9858
rect 0 9800 1643 9802
rect 27846 9860 27906 9936
rect 29520 9860 30000 9890
rect 27846 9800 30000 9860
rect 0 9770 480 9800
rect 1577 9797 1643 9800
rect 5944 9794 6264 9795
rect 5944 9730 5952 9794
rect 6016 9730 6032 9794
rect 6096 9730 6112 9794
rect 6176 9730 6192 9794
rect 6256 9730 6264 9794
rect 5944 9729 6264 9730
rect 15944 9794 16264 9795
rect 15944 9730 15952 9794
rect 16016 9730 16032 9794
rect 16096 9730 16112 9794
rect 16176 9730 16192 9794
rect 16256 9730 16264 9794
rect 15944 9729 16264 9730
rect 25944 9794 26264 9795
rect 25944 9730 25952 9794
rect 26016 9730 26032 9794
rect 26096 9730 26112 9794
rect 26176 9730 26192 9794
rect 26256 9730 26264 9794
rect 29520 9770 30000 9800
rect 25944 9729 26264 9730
rect 3417 9588 3483 9591
rect 4153 9588 4219 9591
rect 23933 9588 23999 9591
rect 3417 9586 4219 9588
rect 3417 9530 3422 9586
rect 3478 9530 4158 9586
rect 4214 9530 4219 9586
rect 3417 9528 4219 9530
rect 3417 9525 3483 9528
rect 4153 9525 4219 9528
rect 4294 9586 23999 9588
rect 4294 9530 23938 9586
rect 23994 9530 23999 9586
rect 4294 9528 23999 9530
rect 3693 9452 3759 9455
rect 4294 9452 4354 9528
rect 23933 9525 23999 9528
rect 23657 9452 23723 9455
rect 3693 9450 4354 9452
rect 3693 9394 3698 9450
rect 3754 9394 4354 9450
rect 3693 9392 4354 9394
rect 4478 9450 23723 9452
rect 4478 9394 23662 9450
rect 23718 9394 23723 9450
rect 4478 9392 23723 9394
rect 3693 9389 3759 9392
rect 0 9316 480 9346
rect 4478 9316 4538 9392
rect 23657 9389 23723 9392
rect 0 9256 4538 9316
rect 24117 9316 24183 9319
rect 29520 9316 30000 9346
rect 24117 9314 30000 9316
rect 24117 9258 24122 9314
rect 24178 9258 30000 9314
rect 24117 9256 30000 9258
rect 0 9226 480 9256
rect 24117 9253 24183 9256
rect 10944 9250 11264 9251
rect 10944 9186 10952 9250
rect 11016 9186 11032 9250
rect 11096 9186 11112 9250
rect 11176 9186 11192 9250
rect 11256 9186 11264 9250
rect 10944 9185 11264 9186
rect 20944 9250 21264 9251
rect 20944 9186 20952 9250
rect 21016 9186 21032 9250
rect 21096 9186 21112 9250
rect 21176 9186 21192 9250
rect 21256 9186 21264 9250
rect 29520 9226 30000 9256
rect 20944 9185 21264 9186
rect 3969 9044 4035 9047
rect 23933 9044 23999 9047
rect 3969 9042 23999 9044
rect 3969 8986 3974 9042
rect 4030 8986 23938 9042
rect 23994 8986 23999 9042
rect 3969 8984 23999 8986
rect 3969 8981 4035 8984
rect 23933 8981 23999 8984
rect 5944 8706 6264 8707
rect 0 8636 480 8666
rect 5944 8642 5952 8706
rect 6016 8642 6032 8706
rect 6096 8642 6112 8706
rect 6176 8642 6192 8706
rect 6256 8642 6264 8706
rect 5944 8641 6264 8642
rect 15944 8706 16264 8707
rect 15944 8642 15952 8706
rect 16016 8642 16032 8706
rect 16096 8642 16112 8706
rect 16176 8642 16192 8706
rect 16256 8642 16264 8706
rect 15944 8641 16264 8642
rect 25944 8706 26264 8707
rect 25944 8642 25952 8706
rect 26016 8642 26032 8706
rect 26096 8642 26112 8706
rect 26176 8642 26192 8706
rect 26256 8642 26264 8706
rect 25944 8641 26264 8642
rect 29520 8636 30000 8666
rect 0 8576 3618 8636
rect 0 8546 480 8576
rect 3558 8364 3618 8576
rect 10550 8576 11714 8636
rect 10550 8364 10610 8576
rect 11654 8364 11714 8576
rect 27846 8576 30000 8636
rect 24117 8500 24183 8503
rect 27846 8500 27906 8576
rect 29520 8546 30000 8576
rect 24117 8498 27906 8500
rect 24117 8442 24122 8498
rect 24178 8442 27906 8498
rect 24117 8440 27906 8442
rect 24117 8437 24183 8440
rect 23565 8364 23631 8367
rect 3558 8304 10610 8364
rect 10734 8304 11530 8364
rect 11654 8362 23631 8364
rect 11654 8306 23570 8362
rect 23626 8306 23631 8362
rect 11654 8304 23631 8306
rect 10734 8228 10794 8304
rect 3374 8168 10794 8228
rect 11470 8228 11530 8304
rect 23565 8301 23631 8304
rect 11470 8168 20362 8228
rect 0 8092 480 8122
rect 3374 8092 3434 8168
rect 10944 8162 11264 8163
rect 10944 8098 10952 8162
rect 11016 8098 11032 8162
rect 11096 8098 11112 8162
rect 11176 8098 11192 8162
rect 11256 8098 11264 8162
rect 10944 8097 11264 8098
rect 0 8032 3434 8092
rect 0 8002 480 8032
rect 20302 7956 20362 8168
rect 20944 8162 21264 8163
rect 20944 8098 20952 8162
rect 21016 8098 21032 8162
rect 21096 8098 21112 8162
rect 21176 8098 21192 8162
rect 21256 8098 21264 8162
rect 20944 8097 21264 8098
rect 24117 8092 24183 8095
rect 29520 8092 30000 8122
rect 24117 8090 30000 8092
rect 24117 8034 24122 8090
rect 24178 8034 30000 8090
rect 24117 8032 30000 8034
rect 24117 8029 24183 8032
rect 29520 8002 30000 8032
rect 23473 7956 23539 7959
rect 3558 7896 19626 7956
rect 20302 7954 23539 7956
rect 20302 7898 23478 7954
rect 23534 7898 23539 7954
rect 20302 7896 23539 7898
rect 0 7412 480 7442
rect 3558 7412 3618 7896
rect 3877 7820 3943 7823
rect 13077 7820 13143 7823
rect 3877 7818 13143 7820
rect 3877 7762 3882 7818
rect 3938 7762 13082 7818
rect 13138 7762 13143 7818
rect 3877 7760 13143 7762
rect 3877 7757 3943 7760
rect 13077 7757 13143 7760
rect 19566 7684 19626 7896
rect 23473 7893 23539 7896
rect 22461 7684 22527 7687
rect 19566 7682 22527 7684
rect 19566 7626 22466 7682
rect 22522 7626 22527 7682
rect 19566 7624 22527 7626
rect 22461 7621 22527 7624
rect 5944 7618 6264 7619
rect 5944 7554 5952 7618
rect 6016 7554 6032 7618
rect 6096 7554 6112 7618
rect 6176 7554 6192 7618
rect 6256 7554 6264 7618
rect 5944 7553 6264 7554
rect 15944 7618 16264 7619
rect 15944 7554 15952 7618
rect 16016 7554 16032 7618
rect 16096 7554 16112 7618
rect 16176 7554 16192 7618
rect 16256 7554 16264 7618
rect 15944 7553 16264 7554
rect 25944 7618 26264 7619
rect 25944 7554 25952 7618
rect 26016 7554 26032 7618
rect 26096 7554 26112 7618
rect 26176 7554 26192 7618
rect 26256 7554 26264 7618
rect 25944 7553 26264 7554
rect 20529 7548 20595 7551
rect 23933 7548 23999 7551
rect 20529 7546 23999 7548
rect 20529 7490 20534 7546
rect 20590 7490 23938 7546
rect 23994 7490 23999 7546
rect 20529 7488 23999 7490
rect 20529 7485 20595 7488
rect 23933 7485 23999 7488
rect 0 7352 3618 7412
rect 3785 7412 3851 7415
rect 18413 7412 18479 7415
rect 3785 7410 18479 7412
rect 3785 7354 3790 7410
rect 3846 7354 18418 7410
rect 18474 7354 18479 7410
rect 3785 7352 18479 7354
rect 0 7322 480 7352
rect 3785 7349 3851 7352
rect 18413 7349 18479 7352
rect 18597 7412 18663 7415
rect 29520 7412 30000 7442
rect 18597 7410 30000 7412
rect 18597 7354 18602 7410
rect 18658 7354 30000 7410
rect 18597 7352 30000 7354
rect 18597 7349 18663 7352
rect 29520 7322 30000 7352
rect 3601 7276 3667 7279
rect 20529 7276 20595 7279
rect 3601 7274 20595 7276
rect 3601 7218 3606 7274
rect 3662 7218 20534 7274
rect 20590 7218 20595 7274
rect 3601 7216 20595 7218
rect 3601 7213 3667 7216
rect 20529 7213 20595 7216
rect 20670 7216 24962 7276
rect 13261 7140 13327 7143
rect 20670 7140 20730 7216
rect 13261 7138 20730 7140
rect 13261 7082 13266 7138
rect 13322 7082 20730 7138
rect 13261 7080 20730 7082
rect 13261 7077 13327 7080
rect 10944 7074 11264 7075
rect 10944 7010 10952 7074
rect 11016 7010 11032 7074
rect 11096 7010 11112 7074
rect 11176 7010 11192 7074
rect 11256 7010 11264 7074
rect 10944 7009 11264 7010
rect 20944 7074 21264 7075
rect 20944 7010 20952 7074
rect 21016 7010 21032 7074
rect 21096 7010 21112 7074
rect 21176 7010 21192 7074
rect 21256 7010 21264 7074
rect 20944 7009 21264 7010
rect 0 6868 480 6898
rect 14917 6868 14983 6871
rect 24902 6868 24962 7216
rect 29520 6868 30000 6898
rect 0 6808 674 6868
rect 0 6778 480 6808
rect 614 6732 674 6808
rect 14917 6866 24410 6868
rect 14917 6810 14922 6866
rect 14978 6810 24410 6866
rect 14917 6808 24410 6810
rect 24902 6808 30000 6868
rect 14917 6805 14983 6808
rect 24117 6732 24183 6735
rect 614 6730 24183 6732
rect 614 6674 24122 6730
rect 24178 6674 24183 6730
rect 614 6672 24183 6674
rect 24117 6669 24183 6672
rect 5944 6530 6264 6531
rect 5944 6466 5952 6530
rect 6016 6466 6032 6530
rect 6096 6466 6112 6530
rect 6176 6466 6192 6530
rect 6256 6466 6264 6530
rect 5944 6465 6264 6466
rect 15944 6530 16264 6531
rect 15944 6466 15952 6530
rect 16016 6466 16032 6530
rect 16096 6466 16112 6530
rect 16176 6466 16192 6530
rect 16256 6466 16264 6530
rect 15944 6465 16264 6466
rect 0 6324 480 6354
rect 1301 6324 1367 6327
rect 0 6322 1367 6324
rect 0 6266 1306 6322
rect 1362 6266 1367 6322
rect 0 6264 1367 6266
rect 24350 6324 24410 6808
rect 29520 6778 30000 6808
rect 25944 6530 26264 6531
rect 25944 6466 25952 6530
rect 26016 6466 26032 6530
rect 26096 6466 26112 6530
rect 26176 6466 26192 6530
rect 26256 6466 26264 6530
rect 25944 6465 26264 6466
rect 29520 6324 30000 6354
rect 24350 6264 30000 6324
rect 0 6234 480 6264
rect 1301 6261 1367 6264
rect 29520 6234 30000 6264
rect 10944 5986 11264 5987
rect 10944 5922 10952 5986
rect 11016 5922 11032 5986
rect 11096 5922 11112 5986
rect 11176 5922 11192 5986
rect 11256 5922 11264 5986
rect 10944 5921 11264 5922
rect 20944 5986 21264 5987
rect 20944 5922 20952 5986
rect 21016 5922 21032 5986
rect 21096 5922 21112 5986
rect 21176 5922 21192 5986
rect 21256 5922 21264 5986
rect 20944 5921 21264 5922
rect 13077 5780 13143 5783
rect 3374 5778 13143 5780
rect 3374 5722 13082 5778
rect 13138 5722 13143 5778
rect 3374 5720 13143 5722
rect 0 5644 480 5674
rect 3374 5644 3434 5720
rect 13077 5717 13143 5720
rect 13629 5780 13695 5783
rect 25589 5780 25655 5783
rect 13629 5778 25655 5780
rect 13629 5722 13634 5778
rect 13690 5722 25594 5778
rect 25650 5722 25655 5778
rect 13629 5720 25655 5722
rect 13629 5717 13695 5720
rect 25589 5717 25655 5720
rect 0 5584 3434 5644
rect 4337 5644 4403 5647
rect 29520 5644 30000 5674
rect 4337 5642 30000 5644
rect 4337 5586 4342 5642
rect 4398 5586 30000 5642
rect 4337 5584 30000 5586
rect 0 5554 480 5584
rect 4337 5581 4403 5584
rect 29520 5554 30000 5584
rect 5944 5442 6264 5443
rect 5944 5378 5952 5442
rect 6016 5378 6032 5442
rect 6096 5378 6112 5442
rect 6176 5378 6192 5442
rect 6256 5378 6264 5442
rect 5944 5377 6264 5378
rect 15944 5442 16264 5443
rect 15944 5378 15952 5442
rect 16016 5378 16032 5442
rect 16096 5378 16112 5442
rect 16176 5378 16192 5442
rect 16256 5378 16264 5442
rect 15944 5377 16264 5378
rect 25944 5442 26264 5443
rect 25944 5378 25952 5442
rect 26016 5378 26032 5442
rect 26096 5378 26112 5442
rect 26176 5378 26192 5442
rect 26256 5378 26264 5442
rect 25944 5377 26264 5378
rect 3509 5236 3575 5239
rect 12617 5236 12683 5239
rect 3509 5234 12683 5236
rect 3509 5178 3514 5234
rect 3570 5178 12622 5234
rect 12678 5178 12683 5234
rect 3509 5176 12683 5178
rect 3509 5173 3575 5176
rect 12617 5173 12683 5176
rect 15561 5236 15627 5239
rect 25681 5236 25747 5239
rect 15561 5234 25747 5236
rect 15561 5178 15566 5234
rect 15622 5178 25686 5234
rect 25742 5178 25747 5234
rect 15561 5176 25747 5178
rect 15561 5173 15627 5176
rect 25681 5173 25747 5176
rect 0 5100 480 5130
rect 24117 5100 24183 5103
rect 0 5098 24183 5100
rect 0 5042 24122 5098
rect 24178 5042 24183 5098
rect 0 5040 24183 5042
rect 0 5010 480 5040
rect 24117 5037 24183 5040
rect 24301 5100 24367 5103
rect 29520 5100 30000 5130
rect 24301 5098 30000 5100
rect 24301 5042 24306 5098
rect 24362 5042 30000 5098
rect 24301 5040 30000 5042
rect 24301 5037 24367 5040
rect 29520 5010 30000 5040
rect 10944 4898 11264 4899
rect 10944 4834 10952 4898
rect 11016 4834 11032 4898
rect 11096 4834 11112 4898
rect 11176 4834 11192 4898
rect 11256 4834 11264 4898
rect 10944 4833 11264 4834
rect 20944 4898 21264 4899
rect 20944 4834 20952 4898
rect 21016 4834 21032 4898
rect 21096 4834 21112 4898
rect 21176 4834 21192 4898
rect 21256 4834 21264 4898
rect 20944 4833 21264 4834
rect 3877 4692 3943 4695
rect 20437 4692 20503 4695
rect 3877 4690 20503 4692
rect 3877 4634 3882 4690
rect 3938 4634 20442 4690
rect 20498 4634 20503 4690
rect 3877 4632 20503 4634
rect 3877 4629 3943 4632
rect 20437 4629 20503 4632
rect 15745 4556 15811 4559
rect 3374 4554 15811 4556
rect 3374 4498 15750 4554
rect 15806 4498 15811 4554
rect 3374 4496 15811 4498
rect 0 4420 480 4450
rect 3374 4420 3434 4496
rect 15745 4493 15811 4496
rect 20621 4556 20687 4559
rect 20621 4554 27906 4556
rect 20621 4498 20626 4554
rect 20682 4498 27906 4554
rect 20621 4496 27906 4498
rect 20621 4493 20687 4496
rect 0 4360 3434 4420
rect 27846 4420 27906 4496
rect 29520 4420 30000 4450
rect 27846 4360 30000 4420
rect 0 4330 480 4360
rect 5944 4354 6264 4355
rect 5944 4290 5952 4354
rect 6016 4290 6032 4354
rect 6096 4290 6112 4354
rect 6176 4290 6192 4354
rect 6256 4290 6264 4354
rect 5944 4289 6264 4290
rect 15944 4354 16264 4355
rect 15944 4290 15952 4354
rect 16016 4290 16032 4354
rect 16096 4290 16112 4354
rect 16176 4290 16192 4354
rect 16256 4290 16264 4354
rect 15944 4289 16264 4290
rect 25944 4354 26264 4355
rect 25944 4290 25952 4354
rect 26016 4290 26032 4354
rect 26096 4290 26112 4354
rect 26176 4290 26192 4354
rect 26256 4290 26264 4354
rect 29520 4330 30000 4360
rect 25944 4289 26264 4290
rect 12801 4148 12867 4151
rect 24301 4148 24367 4151
rect 12801 4146 24367 4148
rect 12801 4090 12806 4146
rect 12862 4090 24306 4146
rect 24362 4090 24367 4146
rect 12801 4088 24367 4090
rect 12801 4085 12867 4088
rect 24301 4085 24367 4088
rect 3417 4012 3483 4015
rect 23933 4012 23999 4015
rect 3417 4010 23999 4012
rect 3417 3954 3422 4010
rect 3478 3954 23938 4010
rect 23994 3954 23999 4010
rect 3417 3952 23999 3954
rect 3417 3949 3483 3952
rect 23933 3949 23999 3952
rect 0 3876 480 3906
rect 24117 3876 24183 3879
rect 29520 3876 30000 3906
rect 0 3816 674 3876
rect 0 3786 480 3816
rect 614 3604 674 3816
rect 24117 3874 30000 3876
rect 24117 3818 24122 3874
rect 24178 3818 30000 3874
rect 24117 3816 30000 3818
rect 24117 3813 24183 3816
rect 10944 3810 11264 3811
rect 10944 3746 10952 3810
rect 11016 3746 11032 3810
rect 11096 3746 11112 3810
rect 11176 3746 11192 3810
rect 11256 3746 11264 3810
rect 10944 3745 11264 3746
rect 20944 3810 21264 3811
rect 20944 3746 20952 3810
rect 21016 3746 21032 3810
rect 21096 3746 21112 3810
rect 21176 3746 21192 3810
rect 21256 3746 21264 3810
rect 29520 3786 30000 3816
rect 20944 3745 21264 3746
rect 20713 3604 20779 3607
rect 614 3602 20779 3604
rect 614 3546 20718 3602
rect 20774 3546 20779 3602
rect 614 3544 20779 3546
rect 20713 3541 20779 3544
rect 24117 3468 24183 3471
rect 3374 3466 24183 3468
rect 3374 3410 24122 3466
rect 24178 3410 24183 3466
rect 3374 3408 24183 3410
rect 0 3332 480 3362
rect 3374 3332 3434 3408
rect 24117 3405 24183 3408
rect 29520 3332 30000 3362
rect 0 3272 3434 3332
rect 27846 3272 30000 3332
rect 0 3242 480 3272
rect 5944 3266 6264 3267
rect 5944 3202 5952 3266
rect 6016 3202 6032 3266
rect 6096 3202 6112 3266
rect 6176 3202 6192 3266
rect 6256 3202 6264 3266
rect 5944 3201 6264 3202
rect 15944 3266 16264 3267
rect 15944 3202 15952 3266
rect 16016 3202 16032 3266
rect 16096 3202 16112 3266
rect 16176 3202 16192 3266
rect 16256 3202 16264 3266
rect 15944 3201 16264 3202
rect 25944 3266 26264 3267
rect 25944 3202 25952 3266
rect 26016 3202 26032 3266
rect 26096 3202 26112 3266
rect 26176 3202 26192 3266
rect 26256 3202 26264 3266
rect 25944 3201 26264 3202
rect 7373 3060 7439 3063
rect 23933 3060 23999 3063
rect 7373 3058 23999 3060
rect 7373 3002 7378 3058
rect 7434 3002 23938 3058
rect 23994 3002 23999 3058
rect 7373 3000 23999 3002
rect 7373 2997 7439 3000
rect 23933 2997 23999 3000
rect 1669 2924 1735 2927
rect 27846 2924 27906 3272
rect 29520 3242 30000 3272
rect 1669 2922 27906 2924
rect 1669 2866 1674 2922
rect 1730 2866 27906 2922
rect 1669 2864 27906 2866
rect 1669 2861 1735 2864
rect 10944 2722 11264 2723
rect 0 2652 480 2682
rect 10944 2658 10952 2722
rect 11016 2658 11032 2722
rect 11096 2658 11112 2722
rect 11176 2658 11192 2722
rect 11256 2658 11264 2722
rect 10944 2657 11264 2658
rect 20944 2722 21264 2723
rect 20944 2658 20952 2722
rect 21016 2658 21032 2722
rect 21096 2658 21112 2722
rect 21176 2658 21192 2722
rect 21256 2658 21264 2722
rect 20944 2657 21264 2658
rect 1761 2652 1827 2655
rect 0 2650 1827 2652
rect 0 2594 1766 2650
rect 1822 2594 1827 2650
rect 0 2592 1827 2594
rect 0 2562 480 2592
rect 1761 2589 1827 2592
rect 24209 2652 24275 2655
rect 29520 2652 30000 2682
rect 24209 2650 30000 2652
rect 24209 2594 24214 2650
rect 24270 2594 30000 2650
rect 24209 2592 30000 2594
rect 24209 2589 24275 2592
rect 29520 2562 30000 2592
rect 2037 2516 2103 2519
rect 982 2514 2103 2516
rect 982 2458 2042 2514
rect 2098 2458 2103 2514
rect 982 2456 2103 2458
rect 0 2108 480 2138
rect 982 2108 1042 2456
rect 2037 2453 2103 2456
rect 8385 2516 8451 2519
rect 25129 2516 25195 2519
rect 8385 2514 25195 2516
rect 8385 2458 8390 2514
rect 8446 2458 25134 2514
rect 25190 2458 25195 2514
rect 8385 2456 25195 2458
rect 8385 2453 8451 2456
rect 25129 2453 25195 2456
rect 2037 2380 2103 2383
rect 25497 2380 25563 2383
rect 2037 2378 25563 2380
rect 2037 2322 2042 2378
rect 2098 2322 25502 2378
rect 25558 2322 25563 2378
rect 2037 2320 25563 2322
rect 2037 2317 2103 2320
rect 25497 2317 25563 2320
rect 5944 2178 6264 2179
rect 5944 2114 5952 2178
rect 6016 2114 6032 2178
rect 6096 2114 6112 2178
rect 6176 2114 6192 2178
rect 6256 2114 6264 2178
rect 5944 2113 6264 2114
rect 15944 2178 16264 2179
rect 15944 2114 15952 2178
rect 16016 2114 16032 2178
rect 16096 2114 16112 2178
rect 16176 2114 16192 2178
rect 16256 2114 16264 2178
rect 15944 2113 16264 2114
rect 25944 2178 26264 2179
rect 25944 2114 25952 2178
rect 26016 2114 26032 2178
rect 26096 2114 26112 2178
rect 26176 2114 26192 2178
rect 26256 2114 26264 2178
rect 25944 2113 26264 2114
rect 29520 2108 30000 2138
rect 0 2048 1042 2108
rect 26926 2048 30000 2108
rect 0 2018 480 2048
rect 12709 1972 12775 1975
rect 24025 1972 24091 1975
rect 12709 1970 24091 1972
rect 12709 1914 12714 1970
rect 12770 1914 24030 1970
rect 24086 1914 24091 1970
rect 12709 1912 24091 1914
rect 12709 1909 12775 1912
rect 24025 1909 24091 1912
rect 26926 1836 26986 2048
rect 29520 2018 30000 2048
rect 21958 1776 26986 1836
rect 9622 1638 9628 1702
rect 9692 1700 9698 1702
rect 12341 1700 12407 1703
rect 9692 1698 12407 1700
rect 9692 1642 12346 1698
rect 12402 1642 12407 1698
rect 9692 1640 12407 1642
rect 9692 1638 9698 1640
rect 12341 1637 12407 1640
rect 12525 1700 12591 1703
rect 21958 1700 22018 1776
rect 12525 1698 22018 1700
rect 12525 1642 12530 1698
rect 12586 1642 22018 1698
rect 12525 1640 22018 1642
rect 12525 1637 12591 1640
rect 24853 1564 24919 1567
rect 24853 1562 29378 1564
rect 24853 1506 24858 1562
rect 24914 1506 29378 1562
rect 24853 1504 29378 1506
rect 24853 1501 24919 1504
rect 0 1428 480 1458
rect 1485 1428 1551 1431
rect 0 1426 1551 1428
rect 0 1370 1490 1426
rect 1546 1370 1551 1426
rect 0 1368 1551 1370
rect 0 1338 480 1368
rect 1485 1365 1551 1368
rect 2129 1428 2195 1431
rect 9622 1428 9628 1430
rect 2129 1426 9628 1428
rect 2129 1370 2134 1426
rect 2190 1370 9628 1426
rect 2129 1368 9628 1370
rect 2129 1365 2195 1368
rect 9622 1366 9628 1368
rect 9692 1366 9698 1430
rect 29318 1428 29378 1504
rect 29520 1428 30000 1458
rect 29318 1368 30000 1428
rect 29520 1338 30000 1368
rect 0 884 480 914
rect 1577 884 1643 887
rect 29520 884 30000 914
rect 0 882 1643 884
rect 0 826 1582 882
rect 1638 826 1643 882
rect 0 824 1643 826
rect 0 794 480 824
rect 1577 821 1643 824
rect 29318 824 30000 884
rect 29318 476 29378 824
rect 29520 794 30000 824
rect 21958 416 29378 476
rect 0 340 480 370
rect 1393 340 1459 343
rect 0 338 1459 340
rect 0 282 1398 338
rect 1454 282 1459 338
rect 0 280 1459 282
rect 0 250 480 280
rect 1393 277 1459 280
rect 9622 278 9628 342
rect 9692 340 9698 342
rect 12341 340 12407 343
rect 9692 338 12407 340
rect 9692 282 12346 338
rect 12402 282 12407 338
rect 9692 280 12407 282
rect 9692 278 9698 280
rect 12341 277 12407 280
rect 12525 340 12591 343
rect 21958 340 22018 416
rect 12525 338 22018 340
rect 12525 282 12530 338
rect 12586 282 22018 338
rect 12525 280 22018 282
rect 25313 340 25379 343
rect 29520 340 30000 370
rect 25313 338 30000 340
rect 25313 282 25318 338
rect 25374 282 30000 338
rect 25313 280 30000 282
rect 12525 277 12591 280
rect 25313 277 25379 280
rect 29520 250 30000 280
rect 9489 68 9555 71
rect 9622 68 9628 70
rect 9489 66 9628 68
rect 9489 10 9494 66
rect 9550 10 9628 66
rect 9489 8 9628 10
rect 9489 5 9555 8
rect 9622 6 9628 8
rect 9692 6 9698 70
<< via3 >>
rect 5952 21758 6016 21762
rect 5952 21702 5956 21758
rect 5956 21702 6012 21758
rect 6012 21702 6016 21758
rect 5952 21698 6016 21702
rect 6032 21758 6096 21762
rect 6032 21702 6036 21758
rect 6036 21702 6092 21758
rect 6092 21702 6096 21758
rect 6032 21698 6096 21702
rect 6112 21758 6176 21762
rect 6112 21702 6116 21758
rect 6116 21702 6172 21758
rect 6172 21702 6176 21758
rect 6112 21698 6176 21702
rect 6192 21758 6256 21762
rect 6192 21702 6196 21758
rect 6196 21702 6252 21758
rect 6252 21702 6256 21758
rect 6192 21698 6256 21702
rect 15952 21758 16016 21762
rect 15952 21702 15956 21758
rect 15956 21702 16012 21758
rect 16012 21702 16016 21758
rect 15952 21698 16016 21702
rect 16032 21758 16096 21762
rect 16032 21702 16036 21758
rect 16036 21702 16092 21758
rect 16092 21702 16096 21758
rect 16032 21698 16096 21702
rect 16112 21758 16176 21762
rect 16112 21702 16116 21758
rect 16116 21702 16172 21758
rect 16172 21702 16176 21758
rect 16112 21698 16176 21702
rect 16192 21758 16256 21762
rect 16192 21702 16196 21758
rect 16196 21702 16252 21758
rect 16252 21702 16256 21758
rect 16192 21698 16256 21702
rect 25952 21758 26016 21762
rect 25952 21702 25956 21758
rect 25956 21702 26012 21758
rect 26012 21702 26016 21758
rect 25952 21698 26016 21702
rect 26032 21758 26096 21762
rect 26032 21702 26036 21758
rect 26036 21702 26092 21758
rect 26092 21702 26096 21758
rect 26032 21698 26096 21702
rect 26112 21758 26176 21762
rect 26112 21702 26116 21758
rect 26116 21702 26172 21758
rect 26172 21702 26176 21758
rect 26112 21698 26176 21702
rect 26192 21758 26256 21762
rect 26192 21702 26196 21758
rect 26196 21702 26252 21758
rect 26252 21702 26256 21758
rect 26192 21698 26256 21702
rect 10952 21214 11016 21218
rect 10952 21158 10956 21214
rect 10956 21158 11012 21214
rect 11012 21158 11016 21214
rect 10952 21154 11016 21158
rect 11032 21214 11096 21218
rect 11032 21158 11036 21214
rect 11036 21158 11092 21214
rect 11092 21158 11096 21214
rect 11032 21154 11096 21158
rect 11112 21214 11176 21218
rect 11112 21158 11116 21214
rect 11116 21158 11172 21214
rect 11172 21158 11176 21214
rect 11112 21154 11176 21158
rect 11192 21214 11256 21218
rect 11192 21158 11196 21214
rect 11196 21158 11252 21214
rect 11252 21158 11256 21214
rect 11192 21154 11256 21158
rect 20952 21214 21016 21218
rect 20952 21158 20956 21214
rect 20956 21158 21012 21214
rect 21012 21158 21016 21214
rect 20952 21154 21016 21158
rect 21032 21214 21096 21218
rect 21032 21158 21036 21214
rect 21036 21158 21092 21214
rect 21092 21158 21096 21214
rect 21032 21154 21096 21158
rect 21112 21214 21176 21218
rect 21112 21158 21116 21214
rect 21116 21158 21172 21214
rect 21172 21158 21176 21214
rect 21112 21154 21176 21158
rect 21192 21214 21256 21218
rect 21192 21158 21196 21214
rect 21196 21158 21252 21214
rect 21252 21158 21256 21214
rect 21192 21154 21256 21158
rect 5952 20670 6016 20674
rect 5952 20614 5956 20670
rect 5956 20614 6012 20670
rect 6012 20614 6016 20670
rect 5952 20610 6016 20614
rect 6032 20670 6096 20674
rect 6032 20614 6036 20670
rect 6036 20614 6092 20670
rect 6092 20614 6096 20670
rect 6032 20610 6096 20614
rect 6112 20670 6176 20674
rect 6112 20614 6116 20670
rect 6116 20614 6172 20670
rect 6172 20614 6176 20670
rect 6112 20610 6176 20614
rect 6192 20670 6256 20674
rect 6192 20614 6196 20670
rect 6196 20614 6252 20670
rect 6252 20614 6256 20670
rect 6192 20610 6256 20614
rect 15952 20670 16016 20674
rect 15952 20614 15956 20670
rect 15956 20614 16012 20670
rect 16012 20614 16016 20670
rect 15952 20610 16016 20614
rect 16032 20670 16096 20674
rect 16032 20614 16036 20670
rect 16036 20614 16092 20670
rect 16092 20614 16096 20670
rect 16032 20610 16096 20614
rect 16112 20670 16176 20674
rect 16112 20614 16116 20670
rect 16116 20614 16172 20670
rect 16172 20614 16176 20670
rect 16112 20610 16176 20614
rect 16192 20670 16256 20674
rect 16192 20614 16196 20670
rect 16196 20614 16252 20670
rect 16252 20614 16256 20670
rect 16192 20610 16256 20614
rect 25952 20670 26016 20674
rect 25952 20614 25956 20670
rect 25956 20614 26012 20670
rect 26012 20614 26016 20670
rect 25952 20610 26016 20614
rect 26032 20670 26096 20674
rect 26032 20614 26036 20670
rect 26036 20614 26092 20670
rect 26092 20614 26096 20670
rect 26032 20610 26096 20614
rect 26112 20670 26176 20674
rect 26112 20614 26116 20670
rect 26116 20614 26172 20670
rect 26172 20614 26176 20670
rect 26112 20610 26176 20614
rect 26192 20670 26256 20674
rect 26192 20614 26196 20670
rect 26196 20614 26252 20670
rect 26252 20614 26256 20670
rect 26192 20610 26256 20614
rect 10952 20126 11016 20130
rect 10952 20070 10956 20126
rect 10956 20070 11012 20126
rect 11012 20070 11016 20126
rect 10952 20066 11016 20070
rect 11032 20126 11096 20130
rect 11032 20070 11036 20126
rect 11036 20070 11092 20126
rect 11092 20070 11096 20126
rect 11032 20066 11096 20070
rect 11112 20126 11176 20130
rect 11112 20070 11116 20126
rect 11116 20070 11172 20126
rect 11172 20070 11176 20126
rect 11112 20066 11176 20070
rect 11192 20126 11256 20130
rect 11192 20070 11196 20126
rect 11196 20070 11252 20126
rect 11252 20070 11256 20126
rect 11192 20066 11256 20070
rect 20952 20126 21016 20130
rect 20952 20070 20956 20126
rect 20956 20070 21012 20126
rect 21012 20070 21016 20126
rect 20952 20066 21016 20070
rect 21032 20126 21096 20130
rect 21032 20070 21036 20126
rect 21036 20070 21092 20126
rect 21092 20070 21096 20126
rect 21032 20066 21096 20070
rect 21112 20126 21176 20130
rect 21112 20070 21116 20126
rect 21116 20070 21172 20126
rect 21172 20070 21176 20126
rect 21112 20066 21176 20070
rect 21192 20126 21256 20130
rect 21192 20070 21196 20126
rect 21196 20070 21252 20126
rect 21252 20070 21256 20126
rect 21192 20066 21256 20070
rect 5952 19582 6016 19586
rect 5952 19526 5956 19582
rect 5956 19526 6012 19582
rect 6012 19526 6016 19582
rect 5952 19522 6016 19526
rect 6032 19582 6096 19586
rect 6032 19526 6036 19582
rect 6036 19526 6092 19582
rect 6092 19526 6096 19582
rect 6032 19522 6096 19526
rect 6112 19582 6176 19586
rect 6112 19526 6116 19582
rect 6116 19526 6172 19582
rect 6172 19526 6176 19582
rect 6112 19522 6176 19526
rect 6192 19582 6256 19586
rect 6192 19526 6196 19582
rect 6196 19526 6252 19582
rect 6252 19526 6256 19582
rect 6192 19522 6256 19526
rect 15952 19582 16016 19586
rect 15952 19526 15956 19582
rect 15956 19526 16012 19582
rect 16012 19526 16016 19582
rect 15952 19522 16016 19526
rect 16032 19582 16096 19586
rect 16032 19526 16036 19582
rect 16036 19526 16092 19582
rect 16092 19526 16096 19582
rect 16032 19522 16096 19526
rect 16112 19582 16176 19586
rect 16112 19526 16116 19582
rect 16116 19526 16172 19582
rect 16172 19526 16176 19582
rect 16112 19522 16176 19526
rect 16192 19582 16256 19586
rect 16192 19526 16196 19582
rect 16196 19526 16252 19582
rect 16252 19526 16256 19582
rect 16192 19522 16256 19526
rect 25952 19582 26016 19586
rect 25952 19526 25956 19582
rect 25956 19526 26012 19582
rect 26012 19526 26016 19582
rect 25952 19522 26016 19526
rect 26032 19582 26096 19586
rect 26032 19526 26036 19582
rect 26036 19526 26092 19582
rect 26092 19526 26096 19582
rect 26032 19522 26096 19526
rect 26112 19582 26176 19586
rect 26112 19526 26116 19582
rect 26116 19526 26172 19582
rect 26172 19526 26176 19582
rect 26112 19522 26176 19526
rect 26192 19582 26256 19586
rect 26192 19526 26196 19582
rect 26196 19526 26252 19582
rect 26252 19526 26256 19582
rect 26192 19522 26256 19526
rect 10952 19038 11016 19042
rect 10952 18982 10956 19038
rect 10956 18982 11012 19038
rect 11012 18982 11016 19038
rect 10952 18978 11016 18982
rect 11032 19038 11096 19042
rect 11032 18982 11036 19038
rect 11036 18982 11092 19038
rect 11092 18982 11096 19038
rect 11032 18978 11096 18982
rect 11112 19038 11176 19042
rect 11112 18982 11116 19038
rect 11116 18982 11172 19038
rect 11172 18982 11176 19038
rect 11112 18978 11176 18982
rect 11192 19038 11256 19042
rect 11192 18982 11196 19038
rect 11196 18982 11252 19038
rect 11252 18982 11256 19038
rect 11192 18978 11256 18982
rect 20952 19038 21016 19042
rect 20952 18982 20956 19038
rect 20956 18982 21012 19038
rect 21012 18982 21016 19038
rect 20952 18978 21016 18982
rect 21032 19038 21096 19042
rect 21032 18982 21036 19038
rect 21036 18982 21092 19038
rect 21092 18982 21096 19038
rect 21032 18978 21096 18982
rect 21112 19038 21176 19042
rect 21112 18982 21116 19038
rect 21116 18982 21172 19038
rect 21172 18982 21176 19038
rect 21112 18978 21176 18982
rect 21192 19038 21256 19042
rect 21192 18982 21196 19038
rect 21196 18982 21252 19038
rect 21252 18982 21256 19038
rect 21192 18978 21256 18982
rect 5952 18494 6016 18498
rect 5952 18438 5956 18494
rect 5956 18438 6012 18494
rect 6012 18438 6016 18494
rect 5952 18434 6016 18438
rect 6032 18494 6096 18498
rect 6032 18438 6036 18494
rect 6036 18438 6092 18494
rect 6092 18438 6096 18494
rect 6032 18434 6096 18438
rect 6112 18494 6176 18498
rect 6112 18438 6116 18494
rect 6116 18438 6172 18494
rect 6172 18438 6176 18494
rect 6112 18434 6176 18438
rect 6192 18494 6256 18498
rect 6192 18438 6196 18494
rect 6196 18438 6252 18494
rect 6252 18438 6256 18494
rect 6192 18434 6256 18438
rect 15952 18494 16016 18498
rect 15952 18438 15956 18494
rect 15956 18438 16012 18494
rect 16012 18438 16016 18494
rect 15952 18434 16016 18438
rect 16032 18494 16096 18498
rect 16032 18438 16036 18494
rect 16036 18438 16092 18494
rect 16092 18438 16096 18494
rect 16032 18434 16096 18438
rect 16112 18494 16176 18498
rect 16112 18438 16116 18494
rect 16116 18438 16172 18494
rect 16172 18438 16176 18494
rect 16112 18434 16176 18438
rect 16192 18494 16256 18498
rect 16192 18438 16196 18494
rect 16196 18438 16252 18494
rect 16252 18438 16256 18494
rect 16192 18434 16256 18438
rect 25952 18494 26016 18498
rect 25952 18438 25956 18494
rect 25956 18438 26012 18494
rect 26012 18438 26016 18494
rect 25952 18434 26016 18438
rect 26032 18494 26096 18498
rect 26032 18438 26036 18494
rect 26036 18438 26092 18494
rect 26092 18438 26096 18494
rect 26032 18434 26096 18438
rect 26112 18494 26176 18498
rect 26112 18438 26116 18494
rect 26116 18438 26172 18494
rect 26172 18438 26176 18494
rect 26112 18434 26176 18438
rect 26192 18494 26256 18498
rect 26192 18438 26196 18494
rect 26196 18438 26252 18494
rect 26252 18438 26256 18494
rect 26192 18434 26256 18438
rect 24900 17958 24964 18022
rect 10952 17950 11016 17954
rect 10952 17894 10956 17950
rect 10956 17894 11012 17950
rect 11012 17894 11016 17950
rect 10952 17890 11016 17894
rect 11032 17950 11096 17954
rect 11032 17894 11036 17950
rect 11036 17894 11092 17950
rect 11092 17894 11096 17950
rect 11032 17890 11096 17894
rect 11112 17950 11176 17954
rect 11112 17894 11116 17950
rect 11116 17894 11172 17950
rect 11172 17894 11176 17950
rect 11112 17890 11176 17894
rect 11192 17950 11256 17954
rect 11192 17894 11196 17950
rect 11196 17894 11252 17950
rect 11252 17894 11256 17950
rect 11192 17890 11256 17894
rect 20952 17950 21016 17954
rect 20952 17894 20956 17950
rect 20956 17894 21012 17950
rect 21012 17894 21016 17950
rect 20952 17890 21016 17894
rect 21032 17950 21096 17954
rect 21032 17894 21036 17950
rect 21036 17894 21092 17950
rect 21092 17894 21096 17950
rect 21032 17890 21096 17894
rect 21112 17950 21176 17954
rect 21112 17894 21116 17950
rect 21116 17894 21172 17950
rect 21172 17894 21176 17950
rect 21112 17890 21176 17894
rect 21192 17950 21256 17954
rect 21192 17894 21196 17950
rect 21196 17894 21252 17950
rect 21252 17894 21256 17950
rect 21192 17890 21256 17894
rect 5952 17406 6016 17410
rect 5952 17350 5956 17406
rect 5956 17350 6012 17406
rect 6012 17350 6016 17406
rect 5952 17346 6016 17350
rect 6032 17406 6096 17410
rect 6032 17350 6036 17406
rect 6036 17350 6092 17406
rect 6092 17350 6096 17406
rect 6032 17346 6096 17350
rect 6112 17406 6176 17410
rect 6112 17350 6116 17406
rect 6116 17350 6172 17406
rect 6172 17350 6176 17406
rect 6112 17346 6176 17350
rect 6192 17406 6256 17410
rect 6192 17350 6196 17406
rect 6196 17350 6252 17406
rect 6252 17350 6256 17406
rect 6192 17346 6256 17350
rect 15952 17406 16016 17410
rect 15952 17350 15956 17406
rect 15956 17350 16012 17406
rect 16012 17350 16016 17406
rect 15952 17346 16016 17350
rect 16032 17406 16096 17410
rect 16032 17350 16036 17406
rect 16036 17350 16092 17406
rect 16092 17350 16096 17406
rect 16032 17346 16096 17350
rect 16112 17406 16176 17410
rect 16112 17350 16116 17406
rect 16116 17350 16172 17406
rect 16172 17350 16176 17406
rect 16112 17346 16176 17350
rect 16192 17406 16256 17410
rect 16192 17350 16196 17406
rect 16196 17350 16252 17406
rect 16252 17350 16256 17406
rect 16192 17346 16256 17350
rect 25952 17406 26016 17410
rect 25952 17350 25956 17406
rect 25956 17350 26012 17406
rect 26012 17350 26016 17406
rect 25952 17346 26016 17350
rect 26032 17406 26096 17410
rect 26032 17350 26036 17406
rect 26036 17350 26092 17406
rect 26092 17350 26096 17406
rect 26032 17346 26096 17350
rect 26112 17406 26176 17410
rect 26112 17350 26116 17406
rect 26116 17350 26172 17406
rect 26172 17350 26176 17406
rect 26112 17346 26176 17350
rect 26192 17406 26256 17410
rect 26192 17350 26196 17406
rect 26196 17350 26252 17406
rect 26252 17350 26256 17406
rect 26192 17346 26256 17350
rect 10952 16862 11016 16866
rect 10952 16806 10956 16862
rect 10956 16806 11012 16862
rect 11012 16806 11016 16862
rect 10952 16802 11016 16806
rect 11032 16862 11096 16866
rect 11032 16806 11036 16862
rect 11036 16806 11092 16862
rect 11092 16806 11096 16862
rect 11032 16802 11096 16806
rect 11112 16862 11176 16866
rect 11112 16806 11116 16862
rect 11116 16806 11172 16862
rect 11172 16806 11176 16862
rect 11112 16802 11176 16806
rect 11192 16862 11256 16866
rect 11192 16806 11196 16862
rect 11196 16806 11252 16862
rect 11252 16806 11256 16862
rect 11192 16802 11256 16806
rect 20952 16862 21016 16866
rect 20952 16806 20956 16862
rect 20956 16806 21012 16862
rect 21012 16806 21016 16862
rect 20952 16802 21016 16806
rect 21032 16862 21096 16866
rect 21032 16806 21036 16862
rect 21036 16806 21092 16862
rect 21092 16806 21096 16862
rect 21032 16802 21096 16806
rect 21112 16862 21176 16866
rect 21112 16806 21116 16862
rect 21116 16806 21172 16862
rect 21172 16806 21176 16862
rect 21112 16802 21176 16806
rect 21192 16862 21256 16866
rect 21192 16806 21196 16862
rect 21196 16806 21252 16862
rect 21252 16806 21256 16862
rect 21192 16802 21256 16806
rect 5952 16318 6016 16322
rect 5952 16262 5956 16318
rect 5956 16262 6012 16318
rect 6012 16262 6016 16318
rect 5952 16258 6016 16262
rect 6032 16318 6096 16322
rect 6032 16262 6036 16318
rect 6036 16262 6092 16318
rect 6092 16262 6096 16318
rect 6032 16258 6096 16262
rect 6112 16318 6176 16322
rect 6112 16262 6116 16318
rect 6116 16262 6172 16318
rect 6172 16262 6176 16318
rect 6112 16258 6176 16262
rect 6192 16318 6256 16322
rect 6192 16262 6196 16318
rect 6196 16262 6252 16318
rect 6252 16262 6256 16318
rect 6192 16258 6256 16262
rect 15952 16318 16016 16322
rect 15952 16262 15956 16318
rect 15956 16262 16012 16318
rect 16012 16262 16016 16318
rect 15952 16258 16016 16262
rect 16032 16318 16096 16322
rect 16032 16262 16036 16318
rect 16036 16262 16092 16318
rect 16092 16262 16096 16318
rect 16032 16258 16096 16262
rect 16112 16318 16176 16322
rect 16112 16262 16116 16318
rect 16116 16262 16172 16318
rect 16172 16262 16176 16318
rect 16112 16258 16176 16262
rect 16192 16318 16256 16322
rect 16192 16262 16196 16318
rect 16196 16262 16252 16318
rect 16252 16262 16256 16318
rect 16192 16258 16256 16262
rect 25952 16318 26016 16322
rect 25952 16262 25956 16318
rect 25956 16262 26012 16318
rect 26012 16262 26016 16318
rect 25952 16258 26016 16262
rect 26032 16318 26096 16322
rect 26032 16262 26036 16318
rect 26036 16262 26092 16318
rect 26092 16262 26096 16318
rect 26032 16258 26096 16262
rect 26112 16318 26176 16322
rect 26112 16262 26116 16318
rect 26116 16262 26172 16318
rect 26172 16262 26176 16318
rect 26112 16258 26176 16262
rect 26192 16318 26256 16322
rect 26192 16262 26196 16318
rect 26196 16262 26252 16318
rect 26252 16262 26256 16318
rect 26192 16258 26256 16262
rect 10952 15774 11016 15778
rect 10952 15718 10956 15774
rect 10956 15718 11012 15774
rect 11012 15718 11016 15774
rect 10952 15714 11016 15718
rect 11032 15774 11096 15778
rect 11032 15718 11036 15774
rect 11036 15718 11092 15774
rect 11092 15718 11096 15774
rect 11032 15714 11096 15718
rect 11112 15774 11176 15778
rect 11112 15718 11116 15774
rect 11116 15718 11172 15774
rect 11172 15718 11176 15774
rect 11112 15714 11176 15718
rect 11192 15774 11256 15778
rect 11192 15718 11196 15774
rect 11196 15718 11252 15774
rect 11252 15718 11256 15774
rect 11192 15714 11256 15718
rect 20952 15774 21016 15778
rect 20952 15718 20956 15774
rect 20956 15718 21012 15774
rect 21012 15718 21016 15774
rect 20952 15714 21016 15718
rect 21032 15774 21096 15778
rect 21032 15718 21036 15774
rect 21036 15718 21092 15774
rect 21092 15718 21096 15774
rect 21032 15714 21096 15718
rect 21112 15774 21176 15778
rect 21112 15718 21116 15774
rect 21116 15718 21172 15774
rect 21172 15718 21176 15774
rect 21112 15714 21176 15718
rect 21192 15774 21256 15778
rect 21192 15718 21196 15774
rect 21196 15718 21252 15774
rect 21252 15718 21256 15774
rect 21192 15714 21256 15718
rect 5952 15230 6016 15234
rect 5952 15174 5956 15230
rect 5956 15174 6012 15230
rect 6012 15174 6016 15230
rect 5952 15170 6016 15174
rect 6032 15230 6096 15234
rect 6032 15174 6036 15230
rect 6036 15174 6092 15230
rect 6092 15174 6096 15230
rect 6032 15170 6096 15174
rect 6112 15230 6176 15234
rect 6112 15174 6116 15230
rect 6116 15174 6172 15230
rect 6172 15174 6176 15230
rect 6112 15170 6176 15174
rect 6192 15230 6256 15234
rect 6192 15174 6196 15230
rect 6196 15174 6252 15230
rect 6252 15174 6256 15230
rect 6192 15170 6256 15174
rect 15952 15230 16016 15234
rect 15952 15174 15956 15230
rect 15956 15174 16012 15230
rect 16012 15174 16016 15230
rect 15952 15170 16016 15174
rect 16032 15230 16096 15234
rect 16032 15174 16036 15230
rect 16036 15174 16092 15230
rect 16092 15174 16096 15230
rect 16032 15170 16096 15174
rect 16112 15230 16176 15234
rect 16112 15174 16116 15230
rect 16116 15174 16172 15230
rect 16172 15174 16176 15230
rect 16112 15170 16176 15174
rect 16192 15230 16256 15234
rect 16192 15174 16196 15230
rect 16196 15174 16252 15230
rect 16252 15174 16256 15230
rect 16192 15170 16256 15174
rect 25952 15230 26016 15234
rect 25952 15174 25956 15230
rect 25956 15174 26012 15230
rect 26012 15174 26016 15230
rect 25952 15170 26016 15174
rect 26032 15230 26096 15234
rect 26032 15174 26036 15230
rect 26036 15174 26092 15230
rect 26092 15174 26096 15230
rect 26032 15170 26096 15174
rect 26112 15230 26176 15234
rect 26112 15174 26116 15230
rect 26116 15174 26172 15230
rect 26172 15174 26176 15230
rect 26112 15170 26176 15174
rect 26192 15230 26256 15234
rect 26192 15174 26196 15230
rect 26196 15174 26252 15230
rect 26252 15174 26256 15230
rect 26192 15170 26256 15174
rect 10952 14686 11016 14690
rect 10952 14630 10956 14686
rect 10956 14630 11012 14686
rect 11012 14630 11016 14686
rect 10952 14626 11016 14630
rect 11032 14686 11096 14690
rect 11032 14630 11036 14686
rect 11036 14630 11092 14686
rect 11092 14630 11096 14686
rect 11032 14626 11096 14630
rect 11112 14686 11176 14690
rect 11112 14630 11116 14686
rect 11116 14630 11172 14686
rect 11172 14630 11176 14686
rect 11112 14626 11176 14630
rect 11192 14686 11256 14690
rect 11192 14630 11196 14686
rect 11196 14630 11252 14686
rect 11252 14630 11256 14686
rect 11192 14626 11256 14630
rect 20952 14686 21016 14690
rect 20952 14630 20956 14686
rect 20956 14630 21012 14686
rect 21012 14630 21016 14686
rect 20952 14626 21016 14630
rect 21032 14686 21096 14690
rect 21032 14630 21036 14686
rect 21036 14630 21092 14686
rect 21092 14630 21096 14686
rect 21032 14626 21096 14630
rect 21112 14686 21176 14690
rect 21112 14630 21116 14686
rect 21116 14630 21172 14686
rect 21172 14630 21176 14686
rect 21112 14626 21176 14630
rect 21192 14686 21256 14690
rect 21192 14630 21196 14686
rect 21196 14630 21252 14686
rect 21252 14630 21256 14686
rect 21192 14626 21256 14630
rect 5952 14142 6016 14146
rect 5952 14086 5956 14142
rect 5956 14086 6012 14142
rect 6012 14086 6016 14142
rect 5952 14082 6016 14086
rect 6032 14142 6096 14146
rect 6032 14086 6036 14142
rect 6036 14086 6092 14142
rect 6092 14086 6096 14142
rect 6032 14082 6096 14086
rect 6112 14142 6176 14146
rect 6112 14086 6116 14142
rect 6116 14086 6172 14142
rect 6172 14086 6176 14142
rect 6112 14082 6176 14086
rect 6192 14142 6256 14146
rect 6192 14086 6196 14142
rect 6196 14086 6252 14142
rect 6252 14086 6256 14142
rect 6192 14082 6256 14086
rect 15952 14142 16016 14146
rect 15952 14086 15956 14142
rect 15956 14086 16012 14142
rect 16012 14086 16016 14142
rect 15952 14082 16016 14086
rect 16032 14142 16096 14146
rect 16032 14086 16036 14142
rect 16036 14086 16092 14142
rect 16092 14086 16096 14142
rect 16032 14082 16096 14086
rect 16112 14142 16176 14146
rect 16112 14086 16116 14142
rect 16116 14086 16172 14142
rect 16172 14086 16176 14142
rect 16112 14082 16176 14086
rect 16192 14142 16256 14146
rect 16192 14086 16196 14142
rect 16196 14086 16252 14142
rect 16252 14086 16256 14142
rect 16192 14082 16256 14086
rect 25952 14142 26016 14146
rect 25952 14086 25956 14142
rect 25956 14086 26012 14142
rect 26012 14086 26016 14142
rect 25952 14082 26016 14086
rect 26032 14142 26096 14146
rect 26032 14086 26036 14142
rect 26036 14086 26092 14142
rect 26092 14086 26096 14142
rect 26032 14082 26096 14086
rect 26112 14142 26176 14146
rect 26112 14086 26116 14142
rect 26116 14086 26172 14142
rect 26172 14086 26176 14142
rect 26112 14082 26176 14086
rect 26192 14142 26256 14146
rect 26192 14086 26196 14142
rect 26196 14086 26252 14142
rect 26252 14086 26256 14142
rect 26192 14082 26256 14086
rect 10952 13598 11016 13602
rect 10952 13542 10956 13598
rect 10956 13542 11012 13598
rect 11012 13542 11016 13598
rect 10952 13538 11016 13542
rect 11032 13598 11096 13602
rect 11032 13542 11036 13598
rect 11036 13542 11092 13598
rect 11092 13542 11096 13598
rect 11032 13538 11096 13542
rect 11112 13598 11176 13602
rect 11112 13542 11116 13598
rect 11116 13542 11172 13598
rect 11172 13542 11176 13598
rect 11112 13538 11176 13542
rect 11192 13598 11256 13602
rect 11192 13542 11196 13598
rect 11196 13542 11252 13598
rect 11252 13542 11256 13598
rect 11192 13538 11256 13542
rect 20952 13598 21016 13602
rect 20952 13542 20956 13598
rect 20956 13542 21012 13598
rect 21012 13542 21016 13598
rect 20952 13538 21016 13542
rect 21032 13598 21096 13602
rect 21032 13542 21036 13598
rect 21036 13542 21092 13598
rect 21092 13542 21096 13598
rect 21032 13538 21096 13542
rect 21112 13598 21176 13602
rect 21112 13542 21116 13598
rect 21116 13542 21172 13598
rect 21172 13542 21176 13598
rect 21112 13538 21176 13542
rect 21192 13598 21256 13602
rect 21192 13542 21196 13598
rect 21196 13542 21252 13598
rect 21252 13542 21256 13598
rect 21192 13538 21256 13542
rect 5952 13054 6016 13058
rect 5952 12998 5956 13054
rect 5956 12998 6012 13054
rect 6012 12998 6016 13054
rect 5952 12994 6016 12998
rect 6032 13054 6096 13058
rect 6032 12998 6036 13054
rect 6036 12998 6092 13054
rect 6092 12998 6096 13054
rect 6032 12994 6096 12998
rect 6112 13054 6176 13058
rect 6112 12998 6116 13054
rect 6116 12998 6172 13054
rect 6172 12998 6176 13054
rect 6112 12994 6176 12998
rect 6192 13054 6256 13058
rect 6192 12998 6196 13054
rect 6196 12998 6252 13054
rect 6252 12998 6256 13054
rect 6192 12994 6256 12998
rect 15952 13054 16016 13058
rect 15952 12998 15956 13054
rect 15956 12998 16012 13054
rect 16012 12998 16016 13054
rect 15952 12994 16016 12998
rect 16032 13054 16096 13058
rect 16032 12998 16036 13054
rect 16036 12998 16092 13054
rect 16092 12998 16096 13054
rect 16032 12994 16096 12998
rect 16112 13054 16176 13058
rect 16112 12998 16116 13054
rect 16116 12998 16172 13054
rect 16172 12998 16176 13054
rect 16112 12994 16176 12998
rect 16192 13054 16256 13058
rect 16192 12998 16196 13054
rect 16196 12998 16252 13054
rect 16252 12998 16256 13054
rect 16192 12994 16256 12998
rect 25952 13054 26016 13058
rect 25952 12998 25956 13054
rect 25956 12998 26012 13054
rect 26012 12998 26016 13054
rect 25952 12994 26016 12998
rect 26032 13054 26096 13058
rect 26032 12998 26036 13054
rect 26036 12998 26092 13054
rect 26092 12998 26096 13054
rect 26032 12994 26096 12998
rect 26112 13054 26176 13058
rect 26112 12998 26116 13054
rect 26116 12998 26172 13054
rect 26172 12998 26176 13054
rect 26112 12994 26176 12998
rect 26192 13054 26256 13058
rect 26192 12998 26196 13054
rect 26196 12998 26252 13054
rect 26252 12998 26256 13054
rect 26192 12994 26256 12998
rect 10952 12510 11016 12514
rect 10952 12454 10956 12510
rect 10956 12454 11012 12510
rect 11012 12454 11016 12510
rect 10952 12450 11016 12454
rect 11032 12510 11096 12514
rect 11032 12454 11036 12510
rect 11036 12454 11092 12510
rect 11092 12454 11096 12510
rect 11032 12450 11096 12454
rect 11112 12510 11176 12514
rect 11112 12454 11116 12510
rect 11116 12454 11172 12510
rect 11172 12454 11176 12510
rect 11112 12450 11176 12454
rect 11192 12510 11256 12514
rect 11192 12454 11196 12510
rect 11196 12454 11252 12510
rect 11252 12454 11256 12510
rect 11192 12450 11256 12454
rect 20952 12510 21016 12514
rect 20952 12454 20956 12510
rect 20956 12454 21012 12510
rect 21012 12454 21016 12510
rect 20952 12450 21016 12454
rect 21032 12510 21096 12514
rect 21032 12454 21036 12510
rect 21036 12454 21092 12510
rect 21092 12454 21096 12510
rect 21032 12450 21096 12454
rect 21112 12510 21176 12514
rect 21112 12454 21116 12510
rect 21116 12454 21172 12510
rect 21172 12454 21176 12510
rect 21112 12450 21176 12454
rect 21192 12510 21256 12514
rect 21192 12454 21196 12510
rect 21196 12454 21252 12510
rect 21252 12454 21256 12510
rect 21192 12450 21256 12454
rect 5952 11966 6016 11970
rect 5952 11910 5956 11966
rect 5956 11910 6012 11966
rect 6012 11910 6016 11966
rect 5952 11906 6016 11910
rect 6032 11966 6096 11970
rect 6032 11910 6036 11966
rect 6036 11910 6092 11966
rect 6092 11910 6096 11966
rect 6032 11906 6096 11910
rect 6112 11966 6176 11970
rect 6112 11910 6116 11966
rect 6116 11910 6172 11966
rect 6172 11910 6176 11966
rect 6112 11906 6176 11910
rect 6192 11966 6256 11970
rect 6192 11910 6196 11966
rect 6196 11910 6252 11966
rect 6252 11910 6256 11966
rect 6192 11906 6256 11910
rect 15952 11966 16016 11970
rect 15952 11910 15956 11966
rect 15956 11910 16012 11966
rect 16012 11910 16016 11966
rect 15952 11906 16016 11910
rect 16032 11966 16096 11970
rect 16032 11910 16036 11966
rect 16036 11910 16092 11966
rect 16092 11910 16096 11966
rect 16032 11906 16096 11910
rect 16112 11966 16176 11970
rect 16112 11910 16116 11966
rect 16116 11910 16172 11966
rect 16172 11910 16176 11966
rect 16112 11906 16176 11910
rect 16192 11966 16256 11970
rect 16192 11910 16196 11966
rect 16196 11910 16252 11966
rect 16252 11910 16256 11966
rect 16192 11906 16256 11910
rect 25952 11966 26016 11970
rect 25952 11910 25956 11966
rect 25956 11910 26012 11966
rect 26012 11910 26016 11966
rect 25952 11906 26016 11910
rect 26032 11966 26096 11970
rect 26032 11910 26036 11966
rect 26036 11910 26092 11966
rect 26092 11910 26096 11966
rect 26032 11906 26096 11910
rect 26112 11966 26176 11970
rect 26112 11910 26116 11966
rect 26116 11910 26172 11966
rect 26172 11910 26176 11966
rect 26112 11906 26176 11910
rect 26192 11966 26256 11970
rect 26192 11910 26196 11966
rect 26196 11910 26252 11966
rect 26252 11910 26256 11966
rect 26192 11906 26256 11910
rect 10952 11422 11016 11426
rect 10952 11366 10956 11422
rect 10956 11366 11012 11422
rect 11012 11366 11016 11422
rect 10952 11362 11016 11366
rect 11032 11422 11096 11426
rect 11032 11366 11036 11422
rect 11036 11366 11092 11422
rect 11092 11366 11096 11422
rect 11032 11362 11096 11366
rect 11112 11422 11176 11426
rect 11112 11366 11116 11422
rect 11116 11366 11172 11422
rect 11172 11366 11176 11422
rect 11112 11362 11176 11366
rect 11192 11422 11256 11426
rect 11192 11366 11196 11422
rect 11196 11366 11252 11422
rect 11252 11366 11256 11422
rect 11192 11362 11256 11366
rect 20952 11422 21016 11426
rect 20952 11366 20956 11422
rect 20956 11366 21012 11422
rect 21012 11366 21016 11422
rect 20952 11362 21016 11366
rect 21032 11422 21096 11426
rect 21032 11366 21036 11422
rect 21036 11366 21092 11422
rect 21092 11366 21096 11422
rect 21032 11362 21096 11366
rect 21112 11422 21176 11426
rect 21112 11366 21116 11422
rect 21116 11366 21172 11422
rect 21172 11366 21176 11422
rect 21112 11362 21176 11366
rect 21192 11422 21256 11426
rect 21192 11366 21196 11422
rect 21196 11366 21252 11422
rect 21252 11366 21256 11422
rect 21192 11362 21256 11366
rect 3372 11022 3436 11086
rect 5952 10878 6016 10882
rect 5952 10822 5956 10878
rect 5956 10822 6012 10878
rect 6012 10822 6016 10878
rect 5952 10818 6016 10822
rect 6032 10878 6096 10882
rect 6032 10822 6036 10878
rect 6036 10822 6092 10878
rect 6092 10822 6096 10878
rect 6032 10818 6096 10822
rect 6112 10878 6176 10882
rect 6112 10822 6116 10878
rect 6116 10822 6172 10878
rect 6172 10822 6176 10878
rect 6112 10818 6176 10822
rect 6192 10878 6256 10882
rect 6192 10822 6196 10878
rect 6196 10822 6252 10878
rect 6252 10822 6256 10878
rect 6192 10818 6256 10822
rect 15952 10878 16016 10882
rect 15952 10822 15956 10878
rect 15956 10822 16012 10878
rect 16012 10822 16016 10878
rect 15952 10818 16016 10822
rect 16032 10878 16096 10882
rect 16032 10822 16036 10878
rect 16036 10822 16092 10878
rect 16092 10822 16096 10878
rect 16032 10818 16096 10822
rect 16112 10878 16176 10882
rect 16112 10822 16116 10878
rect 16116 10822 16172 10878
rect 16172 10822 16176 10878
rect 16112 10818 16176 10822
rect 16192 10878 16256 10882
rect 16192 10822 16196 10878
rect 16196 10822 16252 10878
rect 16252 10822 16256 10878
rect 16192 10818 16256 10822
rect 25952 10878 26016 10882
rect 25952 10822 25956 10878
rect 25956 10822 26012 10878
rect 26012 10822 26016 10878
rect 25952 10818 26016 10822
rect 26032 10878 26096 10882
rect 26032 10822 26036 10878
rect 26036 10822 26092 10878
rect 26092 10822 26096 10878
rect 26032 10818 26096 10822
rect 26112 10878 26176 10882
rect 26112 10822 26116 10878
rect 26116 10822 26172 10878
rect 26172 10822 26176 10878
rect 26112 10818 26176 10822
rect 26192 10878 26256 10882
rect 26192 10822 26196 10878
rect 26196 10822 26252 10878
rect 26252 10822 26256 10878
rect 26192 10818 26256 10822
rect 10952 10334 11016 10338
rect 10952 10278 10956 10334
rect 10956 10278 11012 10334
rect 11012 10278 11016 10334
rect 10952 10274 11016 10278
rect 11032 10334 11096 10338
rect 11032 10278 11036 10334
rect 11036 10278 11092 10334
rect 11092 10278 11096 10334
rect 11032 10274 11096 10278
rect 11112 10334 11176 10338
rect 11112 10278 11116 10334
rect 11116 10278 11172 10334
rect 11172 10278 11176 10334
rect 11112 10274 11176 10278
rect 11192 10334 11256 10338
rect 11192 10278 11196 10334
rect 11196 10278 11252 10334
rect 11252 10278 11256 10334
rect 11192 10274 11256 10278
rect 20952 10334 21016 10338
rect 20952 10278 20956 10334
rect 20956 10278 21012 10334
rect 21012 10278 21016 10334
rect 20952 10274 21016 10278
rect 21032 10334 21096 10338
rect 21032 10278 21036 10334
rect 21036 10278 21092 10334
rect 21092 10278 21096 10334
rect 21032 10274 21096 10278
rect 21112 10334 21176 10338
rect 21112 10278 21116 10334
rect 21116 10278 21172 10334
rect 21172 10278 21176 10334
rect 21112 10274 21176 10278
rect 21192 10334 21256 10338
rect 21192 10278 21196 10334
rect 21196 10278 21252 10334
rect 21252 10278 21256 10334
rect 21192 10274 21256 10278
rect 5952 9790 6016 9794
rect 5952 9734 5956 9790
rect 5956 9734 6012 9790
rect 6012 9734 6016 9790
rect 5952 9730 6016 9734
rect 6032 9790 6096 9794
rect 6032 9734 6036 9790
rect 6036 9734 6092 9790
rect 6092 9734 6096 9790
rect 6032 9730 6096 9734
rect 6112 9790 6176 9794
rect 6112 9734 6116 9790
rect 6116 9734 6172 9790
rect 6172 9734 6176 9790
rect 6112 9730 6176 9734
rect 6192 9790 6256 9794
rect 6192 9734 6196 9790
rect 6196 9734 6252 9790
rect 6252 9734 6256 9790
rect 6192 9730 6256 9734
rect 15952 9790 16016 9794
rect 15952 9734 15956 9790
rect 15956 9734 16012 9790
rect 16012 9734 16016 9790
rect 15952 9730 16016 9734
rect 16032 9790 16096 9794
rect 16032 9734 16036 9790
rect 16036 9734 16092 9790
rect 16092 9734 16096 9790
rect 16032 9730 16096 9734
rect 16112 9790 16176 9794
rect 16112 9734 16116 9790
rect 16116 9734 16172 9790
rect 16172 9734 16176 9790
rect 16112 9730 16176 9734
rect 16192 9790 16256 9794
rect 16192 9734 16196 9790
rect 16196 9734 16252 9790
rect 16252 9734 16256 9790
rect 16192 9730 16256 9734
rect 25952 9790 26016 9794
rect 25952 9734 25956 9790
rect 25956 9734 26012 9790
rect 26012 9734 26016 9790
rect 25952 9730 26016 9734
rect 26032 9790 26096 9794
rect 26032 9734 26036 9790
rect 26036 9734 26092 9790
rect 26092 9734 26096 9790
rect 26032 9730 26096 9734
rect 26112 9790 26176 9794
rect 26112 9734 26116 9790
rect 26116 9734 26172 9790
rect 26172 9734 26176 9790
rect 26112 9730 26176 9734
rect 26192 9790 26256 9794
rect 26192 9734 26196 9790
rect 26196 9734 26252 9790
rect 26252 9734 26256 9790
rect 26192 9730 26256 9734
rect 10952 9246 11016 9250
rect 10952 9190 10956 9246
rect 10956 9190 11012 9246
rect 11012 9190 11016 9246
rect 10952 9186 11016 9190
rect 11032 9246 11096 9250
rect 11032 9190 11036 9246
rect 11036 9190 11092 9246
rect 11092 9190 11096 9246
rect 11032 9186 11096 9190
rect 11112 9246 11176 9250
rect 11112 9190 11116 9246
rect 11116 9190 11172 9246
rect 11172 9190 11176 9246
rect 11112 9186 11176 9190
rect 11192 9246 11256 9250
rect 11192 9190 11196 9246
rect 11196 9190 11252 9246
rect 11252 9190 11256 9246
rect 11192 9186 11256 9190
rect 20952 9246 21016 9250
rect 20952 9190 20956 9246
rect 20956 9190 21012 9246
rect 21012 9190 21016 9246
rect 20952 9186 21016 9190
rect 21032 9246 21096 9250
rect 21032 9190 21036 9246
rect 21036 9190 21092 9246
rect 21092 9190 21096 9246
rect 21032 9186 21096 9190
rect 21112 9246 21176 9250
rect 21112 9190 21116 9246
rect 21116 9190 21172 9246
rect 21172 9190 21176 9246
rect 21112 9186 21176 9190
rect 21192 9246 21256 9250
rect 21192 9190 21196 9246
rect 21196 9190 21252 9246
rect 21252 9190 21256 9246
rect 21192 9186 21256 9190
rect 5952 8702 6016 8706
rect 5952 8646 5956 8702
rect 5956 8646 6012 8702
rect 6012 8646 6016 8702
rect 5952 8642 6016 8646
rect 6032 8702 6096 8706
rect 6032 8646 6036 8702
rect 6036 8646 6092 8702
rect 6092 8646 6096 8702
rect 6032 8642 6096 8646
rect 6112 8702 6176 8706
rect 6112 8646 6116 8702
rect 6116 8646 6172 8702
rect 6172 8646 6176 8702
rect 6112 8642 6176 8646
rect 6192 8702 6256 8706
rect 6192 8646 6196 8702
rect 6196 8646 6252 8702
rect 6252 8646 6256 8702
rect 6192 8642 6256 8646
rect 15952 8702 16016 8706
rect 15952 8646 15956 8702
rect 15956 8646 16012 8702
rect 16012 8646 16016 8702
rect 15952 8642 16016 8646
rect 16032 8702 16096 8706
rect 16032 8646 16036 8702
rect 16036 8646 16092 8702
rect 16092 8646 16096 8702
rect 16032 8642 16096 8646
rect 16112 8702 16176 8706
rect 16112 8646 16116 8702
rect 16116 8646 16172 8702
rect 16172 8646 16176 8702
rect 16112 8642 16176 8646
rect 16192 8702 16256 8706
rect 16192 8646 16196 8702
rect 16196 8646 16252 8702
rect 16252 8646 16256 8702
rect 16192 8642 16256 8646
rect 25952 8702 26016 8706
rect 25952 8646 25956 8702
rect 25956 8646 26012 8702
rect 26012 8646 26016 8702
rect 25952 8642 26016 8646
rect 26032 8702 26096 8706
rect 26032 8646 26036 8702
rect 26036 8646 26092 8702
rect 26092 8646 26096 8702
rect 26032 8642 26096 8646
rect 26112 8702 26176 8706
rect 26112 8646 26116 8702
rect 26116 8646 26172 8702
rect 26172 8646 26176 8702
rect 26112 8642 26176 8646
rect 26192 8702 26256 8706
rect 26192 8646 26196 8702
rect 26196 8646 26252 8702
rect 26252 8646 26256 8702
rect 26192 8642 26256 8646
rect 10952 8158 11016 8162
rect 10952 8102 10956 8158
rect 10956 8102 11012 8158
rect 11012 8102 11016 8158
rect 10952 8098 11016 8102
rect 11032 8158 11096 8162
rect 11032 8102 11036 8158
rect 11036 8102 11092 8158
rect 11092 8102 11096 8158
rect 11032 8098 11096 8102
rect 11112 8158 11176 8162
rect 11112 8102 11116 8158
rect 11116 8102 11172 8158
rect 11172 8102 11176 8158
rect 11112 8098 11176 8102
rect 11192 8158 11256 8162
rect 11192 8102 11196 8158
rect 11196 8102 11252 8158
rect 11252 8102 11256 8158
rect 11192 8098 11256 8102
rect 20952 8158 21016 8162
rect 20952 8102 20956 8158
rect 20956 8102 21012 8158
rect 21012 8102 21016 8158
rect 20952 8098 21016 8102
rect 21032 8158 21096 8162
rect 21032 8102 21036 8158
rect 21036 8102 21092 8158
rect 21092 8102 21096 8158
rect 21032 8098 21096 8102
rect 21112 8158 21176 8162
rect 21112 8102 21116 8158
rect 21116 8102 21172 8158
rect 21172 8102 21176 8158
rect 21112 8098 21176 8102
rect 21192 8158 21256 8162
rect 21192 8102 21196 8158
rect 21196 8102 21252 8158
rect 21252 8102 21256 8158
rect 21192 8098 21256 8102
rect 5952 7614 6016 7618
rect 5952 7558 5956 7614
rect 5956 7558 6012 7614
rect 6012 7558 6016 7614
rect 5952 7554 6016 7558
rect 6032 7614 6096 7618
rect 6032 7558 6036 7614
rect 6036 7558 6092 7614
rect 6092 7558 6096 7614
rect 6032 7554 6096 7558
rect 6112 7614 6176 7618
rect 6112 7558 6116 7614
rect 6116 7558 6172 7614
rect 6172 7558 6176 7614
rect 6112 7554 6176 7558
rect 6192 7614 6256 7618
rect 6192 7558 6196 7614
rect 6196 7558 6252 7614
rect 6252 7558 6256 7614
rect 6192 7554 6256 7558
rect 15952 7614 16016 7618
rect 15952 7558 15956 7614
rect 15956 7558 16012 7614
rect 16012 7558 16016 7614
rect 15952 7554 16016 7558
rect 16032 7614 16096 7618
rect 16032 7558 16036 7614
rect 16036 7558 16092 7614
rect 16092 7558 16096 7614
rect 16032 7554 16096 7558
rect 16112 7614 16176 7618
rect 16112 7558 16116 7614
rect 16116 7558 16172 7614
rect 16172 7558 16176 7614
rect 16112 7554 16176 7558
rect 16192 7614 16256 7618
rect 16192 7558 16196 7614
rect 16196 7558 16252 7614
rect 16252 7558 16256 7614
rect 16192 7554 16256 7558
rect 25952 7614 26016 7618
rect 25952 7558 25956 7614
rect 25956 7558 26012 7614
rect 26012 7558 26016 7614
rect 25952 7554 26016 7558
rect 26032 7614 26096 7618
rect 26032 7558 26036 7614
rect 26036 7558 26092 7614
rect 26092 7558 26096 7614
rect 26032 7554 26096 7558
rect 26112 7614 26176 7618
rect 26112 7558 26116 7614
rect 26116 7558 26172 7614
rect 26172 7558 26176 7614
rect 26112 7554 26176 7558
rect 26192 7614 26256 7618
rect 26192 7558 26196 7614
rect 26196 7558 26252 7614
rect 26252 7558 26256 7614
rect 26192 7554 26256 7558
rect 10952 7070 11016 7074
rect 10952 7014 10956 7070
rect 10956 7014 11012 7070
rect 11012 7014 11016 7070
rect 10952 7010 11016 7014
rect 11032 7070 11096 7074
rect 11032 7014 11036 7070
rect 11036 7014 11092 7070
rect 11092 7014 11096 7070
rect 11032 7010 11096 7014
rect 11112 7070 11176 7074
rect 11112 7014 11116 7070
rect 11116 7014 11172 7070
rect 11172 7014 11176 7070
rect 11112 7010 11176 7014
rect 11192 7070 11256 7074
rect 11192 7014 11196 7070
rect 11196 7014 11252 7070
rect 11252 7014 11256 7070
rect 11192 7010 11256 7014
rect 20952 7070 21016 7074
rect 20952 7014 20956 7070
rect 20956 7014 21012 7070
rect 21012 7014 21016 7070
rect 20952 7010 21016 7014
rect 21032 7070 21096 7074
rect 21032 7014 21036 7070
rect 21036 7014 21092 7070
rect 21092 7014 21096 7070
rect 21032 7010 21096 7014
rect 21112 7070 21176 7074
rect 21112 7014 21116 7070
rect 21116 7014 21172 7070
rect 21172 7014 21176 7070
rect 21112 7010 21176 7014
rect 21192 7070 21256 7074
rect 21192 7014 21196 7070
rect 21196 7014 21252 7070
rect 21252 7014 21256 7070
rect 21192 7010 21256 7014
rect 5952 6526 6016 6530
rect 5952 6470 5956 6526
rect 5956 6470 6012 6526
rect 6012 6470 6016 6526
rect 5952 6466 6016 6470
rect 6032 6526 6096 6530
rect 6032 6470 6036 6526
rect 6036 6470 6092 6526
rect 6092 6470 6096 6526
rect 6032 6466 6096 6470
rect 6112 6526 6176 6530
rect 6112 6470 6116 6526
rect 6116 6470 6172 6526
rect 6172 6470 6176 6526
rect 6112 6466 6176 6470
rect 6192 6526 6256 6530
rect 6192 6470 6196 6526
rect 6196 6470 6252 6526
rect 6252 6470 6256 6526
rect 6192 6466 6256 6470
rect 15952 6526 16016 6530
rect 15952 6470 15956 6526
rect 15956 6470 16012 6526
rect 16012 6470 16016 6526
rect 15952 6466 16016 6470
rect 16032 6526 16096 6530
rect 16032 6470 16036 6526
rect 16036 6470 16092 6526
rect 16092 6470 16096 6526
rect 16032 6466 16096 6470
rect 16112 6526 16176 6530
rect 16112 6470 16116 6526
rect 16116 6470 16172 6526
rect 16172 6470 16176 6526
rect 16112 6466 16176 6470
rect 16192 6526 16256 6530
rect 16192 6470 16196 6526
rect 16196 6470 16252 6526
rect 16252 6470 16256 6526
rect 16192 6466 16256 6470
rect 25952 6526 26016 6530
rect 25952 6470 25956 6526
rect 25956 6470 26012 6526
rect 26012 6470 26016 6526
rect 25952 6466 26016 6470
rect 26032 6526 26096 6530
rect 26032 6470 26036 6526
rect 26036 6470 26092 6526
rect 26092 6470 26096 6526
rect 26032 6466 26096 6470
rect 26112 6526 26176 6530
rect 26112 6470 26116 6526
rect 26116 6470 26172 6526
rect 26172 6470 26176 6526
rect 26112 6466 26176 6470
rect 26192 6526 26256 6530
rect 26192 6470 26196 6526
rect 26196 6470 26252 6526
rect 26252 6470 26256 6526
rect 26192 6466 26256 6470
rect 10952 5982 11016 5986
rect 10952 5926 10956 5982
rect 10956 5926 11012 5982
rect 11012 5926 11016 5982
rect 10952 5922 11016 5926
rect 11032 5982 11096 5986
rect 11032 5926 11036 5982
rect 11036 5926 11092 5982
rect 11092 5926 11096 5982
rect 11032 5922 11096 5926
rect 11112 5982 11176 5986
rect 11112 5926 11116 5982
rect 11116 5926 11172 5982
rect 11172 5926 11176 5982
rect 11112 5922 11176 5926
rect 11192 5982 11256 5986
rect 11192 5926 11196 5982
rect 11196 5926 11252 5982
rect 11252 5926 11256 5982
rect 11192 5922 11256 5926
rect 20952 5982 21016 5986
rect 20952 5926 20956 5982
rect 20956 5926 21012 5982
rect 21012 5926 21016 5982
rect 20952 5922 21016 5926
rect 21032 5982 21096 5986
rect 21032 5926 21036 5982
rect 21036 5926 21092 5982
rect 21092 5926 21096 5982
rect 21032 5922 21096 5926
rect 21112 5982 21176 5986
rect 21112 5926 21116 5982
rect 21116 5926 21172 5982
rect 21172 5926 21176 5982
rect 21112 5922 21176 5926
rect 21192 5982 21256 5986
rect 21192 5926 21196 5982
rect 21196 5926 21252 5982
rect 21252 5926 21256 5982
rect 21192 5922 21256 5926
rect 5952 5438 6016 5442
rect 5952 5382 5956 5438
rect 5956 5382 6012 5438
rect 6012 5382 6016 5438
rect 5952 5378 6016 5382
rect 6032 5438 6096 5442
rect 6032 5382 6036 5438
rect 6036 5382 6092 5438
rect 6092 5382 6096 5438
rect 6032 5378 6096 5382
rect 6112 5438 6176 5442
rect 6112 5382 6116 5438
rect 6116 5382 6172 5438
rect 6172 5382 6176 5438
rect 6112 5378 6176 5382
rect 6192 5438 6256 5442
rect 6192 5382 6196 5438
rect 6196 5382 6252 5438
rect 6252 5382 6256 5438
rect 6192 5378 6256 5382
rect 15952 5438 16016 5442
rect 15952 5382 15956 5438
rect 15956 5382 16012 5438
rect 16012 5382 16016 5438
rect 15952 5378 16016 5382
rect 16032 5438 16096 5442
rect 16032 5382 16036 5438
rect 16036 5382 16092 5438
rect 16092 5382 16096 5438
rect 16032 5378 16096 5382
rect 16112 5438 16176 5442
rect 16112 5382 16116 5438
rect 16116 5382 16172 5438
rect 16172 5382 16176 5438
rect 16112 5378 16176 5382
rect 16192 5438 16256 5442
rect 16192 5382 16196 5438
rect 16196 5382 16252 5438
rect 16252 5382 16256 5438
rect 16192 5378 16256 5382
rect 25952 5438 26016 5442
rect 25952 5382 25956 5438
rect 25956 5382 26012 5438
rect 26012 5382 26016 5438
rect 25952 5378 26016 5382
rect 26032 5438 26096 5442
rect 26032 5382 26036 5438
rect 26036 5382 26092 5438
rect 26092 5382 26096 5438
rect 26032 5378 26096 5382
rect 26112 5438 26176 5442
rect 26112 5382 26116 5438
rect 26116 5382 26172 5438
rect 26172 5382 26176 5438
rect 26112 5378 26176 5382
rect 26192 5438 26256 5442
rect 26192 5382 26196 5438
rect 26196 5382 26252 5438
rect 26252 5382 26256 5438
rect 26192 5378 26256 5382
rect 10952 4894 11016 4898
rect 10952 4838 10956 4894
rect 10956 4838 11012 4894
rect 11012 4838 11016 4894
rect 10952 4834 11016 4838
rect 11032 4894 11096 4898
rect 11032 4838 11036 4894
rect 11036 4838 11092 4894
rect 11092 4838 11096 4894
rect 11032 4834 11096 4838
rect 11112 4894 11176 4898
rect 11112 4838 11116 4894
rect 11116 4838 11172 4894
rect 11172 4838 11176 4894
rect 11112 4834 11176 4838
rect 11192 4894 11256 4898
rect 11192 4838 11196 4894
rect 11196 4838 11252 4894
rect 11252 4838 11256 4894
rect 11192 4834 11256 4838
rect 20952 4894 21016 4898
rect 20952 4838 20956 4894
rect 20956 4838 21012 4894
rect 21012 4838 21016 4894
rect 20952 4834 21016 4838
rect 21032 4894 21096 4898
rect 21032 4838 21036 4894
rect 21036 4838 21092 4894
rect 21092 4838 21096 4894
rect 21032 4834 21096 4838
rect 21112 4894 21176 4898
rect 21112 4838 21116 4894
rect 21116 4838 21172 4894
rect 21172 4838 21176 4894
rect 21112 4834 21176 4838
rect 21192 4894 21256 4898
rect 21192 4838 21196 4894
rect 21196 4838 21252 4894
rect 21252 4838 21256 4894
rect 21192 4834 21256 4838
rect 5952 4350 6016 4354
rect 5952 4294 5956 4350
rect 5956 4294 6012 4350
rect 6012 4294 6016 4350
rect 5952 4290 6016 4294
rect 6032 4350 6096 4354
rect 6032 4294 6036 4350
rect 6036 4294 6092 4350
rect 6092 4294 6096 4350
rect 6032 4290 6096 4294
rect 6112 4350 6176 4354
rect 6112 4294 6116 4350
rect 6116 4294 6172 4350
rect 6172 4294 6176 4350
rect 6112 4290 6176 4294
rect 6192 4350 6256 4354
rect 6192 4294 6196 4350
rect 6196 4294 6252 4350
rect 6252 4294 6256 4350
rect 6192 4290 6256 4294
rect 15952 4350 16016 4354
rect 15952 4294 15956 4350
rect 15956 4294 16012 4350
rect 16012 4294 16016 4350
rect 15952 4290 16016 4294
rect 16032 4350 16096 4354
rect 16032 4294 16036 4350
rect 16036 4294 16092 4350
rect 16092 4294 16096 4350
rect 16032 4290 16096 4294
rect 16112 4350 16176 4354
rect 16112 4294 16116 4350
rect 16116 4294 16172 4350
rect 16172 4294 16176 4350
rect 16112 4290 16176 4294
rect 16192 4350 16256 4354
rect 16192 4294 16196 4350
rect 16196 4294 16252 4350
rect 16252 4294 16256 4350
rect 16192 4290 16256 4294
rect 25952 4350 26016 4354
rect 25952 4294 25956 4350
rect 25956 4294 26012 4350
rect 26012 4294 26016 4350
rect 25952 4290 26016 4294
rect 26032 4350 26096 4354
rect 26032 4294 26036 4350
rect 26036 4294 26092 4350
rect 26092 4294 26096 4350
rect 26032 4290 26096 4294
rect 26112 4350 26176 4354
rect 26112 4294 26116 4350
rect 26116 4294 26172 4350
rect 26172 4294 26176 4350
rect 26112 4290 26176 4294
rect 26192 4350 26256 4354
rect 26192 4294 26196 4350
rect 26196 4294 26252 4350
rect 26252 4294 26256 4350
rect 26192 4290 26256 4294
rect 10952 3806 11016 3810
rect 10952 3750 10956 3806
rect 10956 3750 11012 3806
rect 11012 3750 11016 3806
rect 10952 3746 11016 3750
rect 11032 3806 11096 3810
rect 11032 3750 11036 3806
rect 11036 3750 11092 3806
rect 11092 3750 11096 3806
rect 11032 3746 11096 3750
rect 11112 3806 11176 3810
rect 11112 3750 11116 3806
rect 11116 3750 11172 3806
rect 11172 3750 11176 3806
rect 11112 3746 11176 3750
rect 11192 3806 11256 3810
rect 11192 3750 11196 3806
rect 11196 3750 11252 3806
rect 11252 3750 11256 3806
rect 11192 3746 11256 3750
rect 20952 3806 21016 3810
rect 20952 3750 20956 3806
rect 20956 3750 21012 3806
rect 21012 3750 21016 3806
rect 20952 3746 21016 3750
rect 21032 3806 21096 3810
rect 21032 3750 21036 3806
rect 21036 3750 21092 3806
rect 21092 3750 21096 3806
rect 21032 3746 21096 3750
rect 21112 3806 21176 3810
rect 21112 3750 21116 3806
rect 21116 3750 21172 3806
rect 21172 3750 21176 3806
rect 21112 3746 21176 3750
rect 21192 3806 21256 3810
rect 21192 3750 21196 3806
rect 21196 3750 21252 3806
rect 21252 3750 21256 3806
rect 21192 3746 21256 3750
rect 5952 3262 6016 3266
rect 5952 3206 5956 3262
rect 5956 3206 6012 3262
rect 6012 3206 6016 3262
rect 5952 3202 6016 3206
rect 6032 3262 6096 3266
rect 6032 3206 6036 3262
rect 6036 3206 6092 3262
rect 6092 3206 6096 3262
rect 6032 3202 6096 3206
rect 6112 3262 6176 3266
rect 6112 3206 6116 3262
rect 6116 3206 6172 3262
rect 6172 3206 6176 3262
rect 6112 3202 6176 3206
rect 6192 3262 6256 3266
rect 6192 3206 6196 3262
rect 6196 3206 6252 3262
rect 6252 3206 6256 3262
rect 6192 3202 6256 3206
rect 15952 3262 16016 3266
rect 15952 3206 15956 3262
rect 15956 3206 16012 3262
rect 16012 3206 16016 3262
rect 15952 3202 16016 3206
rect 16032 3262 16096 3266
rect 16032 3206 16036 3262
rect 16036 3206 16092 3262
rect 16092 3206 16096 3262
rect 16032 3202 16096 3206
rect 16112 3262 16176 3266
rect 16112 3206 16116 3262
rect 16116 3206 16172 3262
rect 16172 3206 16176 3262
rect 16112 3202 16176 3206
rect 16192 3262 16256 3266
rect 16192 3206 16196 3262
rect 16196 3206 16252 3262
rect 16252 3206 16256 3262
rect 16192 3202 16256 3206
rect 25952 3262 26016 3266
rect 25952 3206 25956 3262
rect 25956 3206 26012 3262
rect 26012 3206 26016 3262
rect 25952 3202 26016 3206
rect 26032 3262 26096 3266
rect 26032 3206 26036 3262
rect 26036 3206 26092 3262
rect 26092 3206 26096 3262
rect 26032 3202 26096 3206
rect 26112 3262 26176 3266
rect 26112 3206 26116 3262
rect 26116 3206 26172 3262
rect 26172 3206 26176 3262
rect 26112 3202 26176 3206
rect 26192 3262 26256 3266
rect 26192 3206 26196 3262
rect 26196 3206 26252 3262
rect 26252 3206 26256 3262
rect 26192 3202 26256 3206
rect 10952 2718 11016 2722
rect 10952 2662 10956 2718
rect 10956 2662 11012 2718
rect 11012 2662 11016 2718
rect 10952 2658 11016 2662
rect 11032 2718 11096 2722
rect 11032 2662 11036 2718
rect 11036 2662 11092 2718
rect 11092 2662 11096 2718
rect 11032 2658 11096 2662
rect 11112 2718 11176 2722
rect 11112 2662 11116 2718
rect 11116 2662 11172 2718
rect 11172 2662 11176 2718
rect 11112 2658 11176 2662
rect 11192 2718 11256 2722
rect 11192 2662 11196 2718
rect 11196 2662 11252 2718
rect 11252 2662 11256 2718
rect 11192 2658 11256 2662
rect 20952 2718 21016 2722
rect 20952 2662 20956 2718
rect 20956 2662 21012 2718
rect 21012 2662 21016 2718
rect 20952 2658 21016 2662
rect 21032 2718 21096 2722
rect 21032 2662 21036 2718
rect 21036 2662 21092 2718
rect 21092 2662 21096 2718
rect 21032 2658 21096 2662
rect 21112 2718 21176 2722
rect 21112 2662 21116 2718
rect 21116 2662 21172 2718
rect 21172 2662 21176 2718
rect 21112 2658 21176 2662
rect 21192 2718 21256 2722
rect 21192 2662 21196 2718
rect 21196 2662 21252 2718
rect 21252 2662 21256 2718
rect 21192 2658 21256 2662
rect 5952 2174 6016 2178
rect 5952 2118 5956 2174
rect 5956 2118 6012 2174
rect 6012 2118 6016 2174
rect 5952 2114 6016 2118
rect 6032 2174 6096 2178
rect 6032 2118 6036 2174
rect 6036 2118 6092 2174
rect 6092 2118 6096 2174
rect 6032 2114 6096 2118
rect 6112 2174 6176 2178
rect 6112 2118 6116 2174
rect 6116 2118 6172 2174
rect 6172 2118 6176 2174
rect 6112 2114 6176 2118
rect 6192 2174 6256 2178
rect 6192 2118 6196 2174
rect 6196 2118 6252 2174
rect 6252 2118 6256 2174
rect 6192 2114 6256 2118
rect 15952 2174 16016 2178
rect 15952 2118 15956 2174
rect 15956 2118 16012 2174
rect 16012 2118 16016 2174
rect 15952 2114 16016 2118
rect 16032 2174 16096 2178
rect 16032 2118 16036 2174
rect 16036 2118 16092 2174
rect 16092 2118 16096 2174
rect 16032 2114 16096 2118
rect 16112 2174 16176 2178
rect 16112 2118 16116 2174
rect 16116 2118 16172 2174
rect 16172 2118 16176 2174
rect 16112 2114 16176 2118
rect 16192 2174 16256 2178
rect 16192 2118 16196 2174
rect 16196 2118 16252 2174
rect 16252 2118 16256 2174
rect 16192 2114 16256 2118
rect 25952 2174 26016 2178
rect 25952 2118 25956 2174
rect 25956 2118 26012 2174
rect 26012 2118 26016 2174
rect 25952 2114 26016 2118
rect 26032 2174 26096 2178
rect 26032 2118 26036 2174
rect 26036 2118 26092 2174
rect 26092 2118 26096 2174
rect 26032 2114 26096 2118
rect 26112 2174 26176 2178
rect 26112 2118 26116 2174
rect 26116 2118 26172 2174
rect 26172 2118 26176 2174
rect 26112 2114 26176 2118
rect 26192 2174 26256 2178
rect 26192 2118 26196 2174
rect 26196 2118 26252 2174
rect 26252 2118 26256 2174
rect 26192 2114 26256 2118
rect 9628 1638 9692 1702
rect 9628 1366 9692 1430
rect 9628 278 9692 342
rect 9628 6 9692 70
<< metal4 >>
rect 5944 21762 6264 21778
rect 5944 21698 5952 21762
rect 6016 21698 6032 21762
rect 6096 21698 6112 21762
rect 6176 21698 6192 21762
rect 6256 21698 6264 21762
rect 5944 20674 6264 21698
rect 5944 20610 5952 20674
rect 6016 20610 6032 20674
rect 6096 20610 6112 20674
rect 6176 20610 6192 20674
rect 6256 20610 6264 20674
rect 5944 19586 6264 20610
rect 5944 19522 5952 19586
rect 6016 19522 6032 19586
rect 6096 19522 6112 19586
rect 6176 19522 6192 19586
rect 6256 19522 6264 19586
rect 5944 18498 6264 19522
rect 5944 18434 5952 18498
rect 6016 18434 6032 18498
rect 6096 18434 6112 18498
rect 6176 18434 6192 18498
rect 6256 18434 6264 18498
rect 5944 17410 6264 18434
rect 5944 17346 5952 17410
rect 6016 17346 6032 17410
rect 6096 17346 6112 17410
rect 6176 17346 6192 17410
rect 6256 17346 6264 17410
rect 5944 16322 6264 17346
rect 5944 16258 5952 16322
rect 6016 16258 6032 16322
rect 6096 16258 6112 16322
rect 6176 16258 6192 16322
rect 6256 16258 6264 16322
rect 5944 15234 6264 16258
rect 5944 15170 5952 15234
rect 6016 15170 6032 15234
rect 6096 15170 6112 15234
rect 6176 15170 6192 15234
rect 6256 15170 6264 15234
rect 5944 14146 6264 15170
rect 5944 14082 5952 14146
rect 6016 14082 6032 14146
rect 6096 14082 6112 14146
rect 6176 14082 6192 14146
rect 6256 14082 6264 14146
rect 5944 13058 6264 14082
rect 5944 12994 5952 13058
rect 6016 12994 6032 13058
rect 6096 12994 6112 13058
rect 6176 12994 6192 13058
rect 6256 12994 6264 13058
rect 5944 11970 6264 12994
rect 5944 11906 5952 11970
rect 6016 11906 6032 11970
rect 6096 11906 6112 11970
rect 6176 11906 6192 11970
rect 6256 11906 6264 11970
rect 3374 11087 3434 11752
rect 3371 11086 3437 11087
rect 3371 11022 3372 11086
rect 3436 11022 3437 11086
rect 3371 11021 3437 11022
rect 5944 10882 6264 11906
rect 5944 10818 5952 10882
rect 6016 10818 6032 10882
rect 6096 10818 6112 10882
rect 6176 10818 6192 10882
rect 6256 10818 6264 10882
rect 5944 9794 6264 10818
rect 5944 9730 5952 9794
rect 6016 9730 6032 9794
rect 6096 9730 6112 9794
rect 6176 9730 6192 9794
rect 6256 9730 6264 9794
rect 5944 8706 6264 9730
rect 5944 8642 5952 8706
rect 6016 8642 6032 8706
rect 6096 8642 6112 8706
rect 6176 8642 6192 8706
rect 6256 8642 6264 8706
rect 5944 7618 6264 8642
rect 5944 7554 5952 7618
rect 6016 7554 6032 7618
rect 6096 7554 6112 7618
rect 6176 7554 6192 7618
rect 6256 7554 6264 7618
rect 5944 6530 6264 7554
rect 5944 6466 5952 6530
rect 6016 6466 6032 6530
rect 6096 6466 6112 6530
rect 6176 6466 6192 6530
rect 6256 6466 6264 6530
rect 5944 5442 6264 6466
rect 5944 5378 5952 5442
rect 6016 5378 6032 5442
rect 6096 5378 6112 5442
rect 6176 5378 6192 5442
rect 6256 5378 6264 5442
rect 5944 4354 6264 5378
rect 5944 4290 5952 4354
rect 6016 4290 6032 4354
rect 6096 4290 6112 4354
rect 6176 4290 6192 4354
rect 6256 4290 6264 4354
rect 5944 3266 6264 4290
rect 5944 3202 5952 3266
rect 6016 3202 6032 3266
rect 6096 3202 6112 3266
rect 6176 3202 6192 3266
rect 6256 3202 6264 3266
rect 5944 2178 6264 3202
rect 5944 2114 5952 2178
rect 6016 2114 6032 2178
rect 6096 2114 6112 2178
rect 6176 2114 6192 2178
rect 6256 2114 6264 2178
rect 5944 2098 6264 2114
rect 10944 21218 11264 21778
rect 10944 21154 10952 21218
rect 11016 21154 11032 21218
rect 11096 21154 11112 21218
rect 11176 21154 11192 21218
rect 11256 21154 11264 21218
rect 10944 20130 11264 21154
rect 10944 20066 10952 20130
rect 11016 20066 11032 20130
rect 11096 20066 11112 20130
rect 11176 20066 11192 20130
rect 11256 20066 11264 20130
rect 10944 19042 11264 20066
rect 10944 18978 10952 19042
rect 11016 18978 11032 19042
rect 11096 18978 11112 19042
rect 11176 18978 11192 19042
rect 11256 18978 11264 19042
rect 10944 17954 11264 18978
rect 10944 17890 10952 17954
rect 11016 17890 11032 17954
rect 11096 17890 11112 17954
rect 11176 17890 11192 17954
rect 11256 17890 11264 17954
rect 10944 16866 11264 17890
rect 10944 16802 10952 16866
rect 11016 16802 11032 16866
rect 11096 16802 11112 16866
rect 11176 16802 11192 16866
rect 11256 16802 11264 16866
rect 10944 15778 11264 16802
rect 10944 15714 10952 15778
rect 11016 15714 11032 15778
rect 11096 15714 11112 15778
rect 11176 15714 11192 15778
rect 11256 15714 11264 15778
rect 10944 14690 11264 15714
rect 10944 14626 10952 14690
rect 11016 14626 11032 14690
rect 11096 14626 11112 14690
rect 11176 14626 11192 14690
rect 11256 14626 11264 14690
rect 10944 13602 11264 14626
rect 10944 13538 10952 13602
rect 11016 13538 11032 13602
rect 11096 13538 11112 13602
rect 11176 13538 11192 13602
rect 11256 13538 11264 13602
rect 10944 12514 11264 13538
rect 10944 12450 10952 12514
rect 11016 12450 11032 12514
rect 11096 12450 11112 12514
rect 11176 12450 11192 12514
rect 11256 12450 11264 12514
rect 10944 11426 11264 12450
rect 10944 11362 10952 11426
rect 11016 11362 11032 11426
rect 11096 11362 11112 11426
rect 11176 11362 11192 11426
rect 11256 11362 11264 11426
rect 10944 10338 11264 11362
rect 10944 10274 10952 10338
rect 11016 10274 11032 10338
rect 11096 10274 11112 10338
rect 11176 10274 11192 10338
rect 11256 10274 11264 10338
rect 10944 9250 11264 10274
rect 10944 9186 10952 9250
rect 11016 9186 11032 9250
rect 11096 9186 11112 9250
rect 11176 9186 11192 9250
rect 11256 9186 11264 9250
rect 10944 8162 11264 9186
rect 10944 8098 10952 8162
rect 11016 8098 11032 8162
rect 11096 8098 11112 8162
rect 11176 8098 11192 8162
rect 11256 8098 11264 8162
rect 10944 7074 11264 8098
rect 10944 7010 10952 7074
rect 11016 7010 11032 7074
rect 11096 7010 11112 7074
rect 11176 7010 11192 7074
rect 11256 7010 11264 7074
rect 10944 5986 11264 7010
rect 10944 5922 10952 5986
rect 11016 5922 11032 5986
rect 11096 5922 11112 5986
rect 11176 5922 11192 5986
rect 11256 5922 11264 5986
rect 10944 4898 11264 5922
rect 10944 4834 10952 4898
rect 11016 4834 11032 4898
rect 11096 4834 11112 4898
rect 11176 4834 11192 4898
rect 11256 4834 11264 4898
rect 10944 3810 11264 4834
rect 10944 3746 10952 3810
rect 11016 3746 11032 3810
rect 11096 3746 11112 3810
rect 11176 3746 11192 3810
rect 11256 3746 11264 3810
rect 10944 2722 11264 3746
rect 10944 2658 10952 2722
rect 11016 2658 11032 2722
rect 11096 2658 11112 2722
rect 11176 2658 11192 2722
rect 11256 2658 11264 2722
rect 10944 2098 11264 2658
rect 15944 21762 16264 21778
rect 15944 21698 15952 21762
rect 16016 21698 16032 21762
rect 16096 21698 16112 21762
rect 16176 21698 16192 21762
rect 16256 21698 16264 21762
rect 15944 20674 16264 21698
rect 15944 20610 15952 20674
rect 16016 20610 16032 20674
rect 16096 20610 16112 20674
rect 16176 20610 16192 20674
rect 16256 20610 16264 20674
rect 15944 19586 16264 20610
rect 15944 19522 15952 19586
rect 16016 19522 16032 19586
rect 16096 19522 16112 19586
rect 16176 19522 16192 19586
rect 16256 19522 16264 19586
rect 15944 18498 16264 19522
rect 15944 18434 15952 18498
rect 16016 18434 16032 18498
rect 16096 18434 16112 18498
rect 16176 18434 16192 18498
rect 16256 18434 16264 18498
rect 15944 17410 16264 18434
rect 15944 17346 15952 17410
rect 16016 17346 16032 17410
rect 16096 17346 16112 17410
rect 16176 17346 16192 17410
rect 16256 17346 16264 17410
rect 15944 16322 16264 17346
rect 15944 16258 15952 16322
rect 16016 16258 16032 16322
rect 16096 16258 16112 16322
rect 16176 16258 16192 16322
rect 16256 16258 16264 16322
rect 15944 15234 16264 16258
rect 15944 15170 15952 15234
rect 16016 15170 16032 15234
rect 16096 15170 16112 15234
rect 16176 15170 16192 15234
rect 16256 15170 16264 15234
rect 15944 14146 16264 15170
rect 15944 14082 15952 14146
rect 16016 14082 16032 14146
rect 16096 14082 16112 14146
rect 16176 14082 16192 14146
rect 16256 14082 16264 14146
rect 15944 13058 16264 14082
rect 15944 12994 15952 13058
rect 16016 12994 16032 13058
rect 16096 12994 16112 13058
rect 16176 12994 16192 13058
rect 16256 12994 16264 13058
rect 15944 11970 16264 12994
rect 15944 11906 15952 11970
rect 16016 11906 16032 11970
rect 16096 11906 16112 11970
rect 16176 11906 16192 11970
rect 16256 11906 16264 11970
rect 15944 10882 16264 11906
rect 15944 10818 15952 10882
rect 16016 10818 16032 10882
rect 16096 10818 16112 10882
rect 16176 10818 16192 10882
rect 16256 10818 16264 10882
rect 15944 9794 16264 10818
rect 15944 9730 15952 9794
rect 16016 9730 16032 9794
rect 16096 9730 16112 9794
rect 16176 9730 16192 9794
rect 16256 9730 16264 9794
rect 15944 8706 16264 9730
rect 15944 8642 15952 8706
rect 16016 8642 16032 8706
rect 16096 8642 16112 8706
rect 16176 8642 16192 8706
rect 16256 8642 16264 8706
rect 15944 7618 16264 8642
rect 15944 7554 15952 7618
rect 16016 7554 16032 7618
rect 16096 7554 16112 7618
rect 16176 7554 16192 7618
rect 16256 7554 16264 7618
rect 15944 6530 16264 7554
rect 15944 6466 15952 6530
rect 16016 6466 16032 6530
rect 16096 6466 16112 6530
rect 16176 6466 16192 6530
rect 16256 6466 16264 6530
rect 15944 5442 16264 6466
rect 15944 5378 15952 5442
rect 16016 5378 16032 5442
rect 16096 5378 16112 5442
rect 16176 5378 16192 5442
rect 16256 5378 16264 5442
rect 15944 4354 16264 5378
rect 15944 4290 15952 4354
rect 16016 4290 16032 4354
rect 16096 4290 16112 4354
rect 16176 4290 16192 4354
rect 16256 4290 16264 4354
rect 15944 3266 16264 4290
rect 15944 3202 15952 3266
rect 16016 3202 16032 3266
rect 16096 3202 16112 3266
rect 16176 3202 16192 3266
rect 16256 3202 16264 3266
rect 15944 2178 16264 3202
rect 15944 2114 15952 2178
rect 16016 2114 16032 2178
rect 16096 2114 16112 2178
rect 16176 2114 16192 2178
rect 16256 2114 16264 2178
rect 15944 2098 16264 2114
rect 20944 21218 21264 21778
rect 20944 21154 20952 21218
rect 21016 21154 21032 21218
rect 21096 21154 21112 21218
rect 21176 21154 21192 21218
rect 21256 21154 21264 21218
rect 20944 20130 21264 21154
rect 20944 20066 20952 20130
rect 21016 20066 21032 20130
rect 21096 20066 21112 20130
rect 21176 20066 21192 20130
rect 21256 20066 21264 20130
rect 20944 19042 21264 20066
rect 20944 18978 20952 19042
rect 21016 18978 21032 19042
rect 21096 18978 21112 19042
rect 21176 18978 21192 19042
rect 21256 18978 21264 19042
rect 20944 17954 21264 18978
rect 25944 21762 26264 21778
rect 25944 21698 25952 21762
rect 26016 21698 26032 21762
rect 26096 21698 26112 21762
rect 26176 21698 26192 21762
rect 26256 21698 26264 21762
rect 25944 20674 26264 21698
rect 25944 20610 25952 20674
rect 26016 20610 26032 20674
rect 26096 20610 26112 20674
rect 26176 20610 26192 20674
rect 26256 20610 26264 20674
rect 25944 19586 26264 20610
rect 25944 19522 25952 19586
rect 26016 19522 26032 19586
rect 26096 19522 26112 19586
rect 26176 19522 26192 19586
rect 26256 19522 26264 19586
rect 25944 18498 26264 19522
rect 25944 18434 25952 18498
rect 26016 18434 26032 18498
rect 26096 18434 26112 18498
rect 26176 18434 26192 18498
rect 26256 18434 26264 18498
rect 24899 18022 24965 18023
rect 24899 17958 24900 18022
rect 24964 17958 24965 18022
rect 24899 17957 24965 17958
rect 20944 17890 20952 17954
rect 21016 17890 21032 17954
rect 21096 17890 21112 17954
rect 21176 17890 21192 17954
rect 21256 17890 21264 17954
rect 20944 16866 21264 17890
rect 20944 16802 20952 16866
rect 21016 16802 21032 16866
rect 21096 16802 21112 16866
rect 21176 16802 21192 16866
rect 21256 16802 21264 16866
rect 20944 15778 21264 16802
rect 20944 15714 20952 15778
rect 21016 15714 21032 15778
rect 21096 15714 21112 15778
rect 21176 15714 21192 15778
rect 21256 15714 21264 15778
rect 20944 14690 21264 15714
rect 20944 14626 20952 14690
rect 21016 14626 21032 14690
rect 21096 14626 21112 14690
rect 21176 14626 21192 14690
rect 21256 14626 21264 14690
rect 20944 13602 21264 14626
rect 20944 13538 20952 13602
rect 21016 13538 21032 13602
rect 21096 13538 21112 13602
rect 21176 13538 21192 13602
rect 21256 13538 21264 13602
rect 20944 12514 21264 13538
rect 20944 12450 20952 12514
rect 21016 12450 21032 12514
rect 21096 12450 21112 12514
rect 21176 12450 21192 12514
rect 21256 12450 21264 12514
rect 20944 11426 21264 12450
rect 24902 11988 24962 17957
rect 25944 17410 26264 18434
rect 25944 17346 25952 17410
rect 26016 17346 26032 17410
rect 26096 17346 26112 17410
rect 26176 17346 26192 17410
rect 26256 17346 26264 17410
rect 25944 16322 26264 17346
rect 25944 16258 25952 16322
rect 26016 16258 26032 16322
rect 26096 16258 26112 16322
rect 26176 16258 26192 16322
rect 26256 16258 26264 16322
rect 25944 15234 26264 16258
rect 25944 15170 25952 15234
rect 26016 15170 26032 15234
rect 26096 15170 26112 15234
rect 26176 15170 26192 15234
rect 26256 15170 26264 15234
rect 25944 14146 26264 15170
rect 25944 14082 25952 14146
rect 26016 14082 26032 14146
rect 26096 14082 26112 14146
rect 26176 14082 26192 14146
rect 26256 14082 26264 14146
rect 25944 13058 26264 14082
rect 25944 12994 25952 13058
rect 26016 12994 26032 13058
rect 26096 12994 26112 13058
rect 26176 12994 26192 13058
rect 26256 12994 26264 13058
rect 25944 11970 26264 12994
rect 25944 11906 25952 11970
rect 26016 11906 26032 11970
rect 26096 11906 26112 11970
rect 26176 11906 26192 11970
rect 26256 11906 26264 11970
rect 20944 11362 20952 11426
rect 21016 11362 21032 11426
rect 21096 11362 21112 11426
rect 21176 11362 21192 11426
rect 21256 11362 21264 11426
rect 20944 10338 21264 11362
rect 20944 10274 20952 10338
rect 21016 10274 21032 10338
rect 21096 10274 21112 10338
rect 21176 10274 21192 10338
rect 21256 10274 21264 10338
rect 20944 9250 21264 10274
rect 20944 9186 20952 9250
rect 21016 9186 21032 9250
rect 21096 9186 21112 9250
rect 21176 9186 21192 9250
rect 21256 9186 21264 9250
rect 20944 8162 21264 9186
rect 20944 8098 20952 8162
rect 21016 8098 21032 8162
rect 21096 8098 21112 8162
rect 21176 8098 21192 8162
rect 21256 8098 21264 8162
rect 20944 7074 21264 8098
rect 20944 7010 20952 7074
rect 21016 7010 21032 7074
rect 21096 7010 21112 7074
rect 21176 7010 21192 7074
rect 21256 7010 21264 7074
rect 20944 5986 21264 7010
rect 20944 5922 20952 5986
rect 21016 5922 21032 5986
rect 21096 5922 21112 5986
rect 21176 5922 21192 5986
rect 21256 5922 21264 5986
rect 20944 4898 21264 5922
rect 20944 4834 20952 4898
rect 21016 4834 21032 4898
rect 21096 4834 21112 4898
rect 21176 4834 21192 4898
rect 21256 4834 21264 4898
rect 20944 3810 21264 4834
rect 20944 3746 20952 3810
rect 21016 3746 21032 3810
rect 21096 3746 21112 3810
rect 21176 3746 21192 3810
rect 21256 3746 21264 3810
rect 20944 2722 21264 3746
rect 20944 2658 20952 2722
rect 21016 2658 21032 2722
rect 21096 2658 21112 2722
rect 21176 2658 21192 2722
rect 21256 2658 21264 2722
rect 20944 2098 21264 2658
rect 25944 10882 26264 11906
rect 25944 10818 25952 10882
rect 26016 10818 26032 10882
rect 26096 10818 26112 10882
rect 26176 10818 26192 10882
rect 26256 10818 26264 10882
rect 25944 9794 26264 10818
rect 25944 9730 25952 9794
rect 26016 9730 26032 9794
rect 26096 9730 26112 9794
rect 26176 9730 26192 9794
rect 26256 9730 26264 9794
rect 25944 8706 26264 9730
rect 25944 8642 25952 8706
rect 26016 8642 26032 8706
rect 26096 8642 26112 8706
rect 26176 8642 26192 8706
rect 26256 8642 26264 8706
rect 25944 7618 26264 8642
rect 25944 7554 25952 7618
rect 26016 7554 26032 7618
rect 26096 7554 26112 7618
rect 26176 7554 26192 7618
rect 26256 7554 26264 7618
rect 25944 6530 26264 7554
rect 25944 6466 25952 6530
rect 26016 6466 26032 6530
rect 26096 6466 26112 6530
rect 26176 6466 26192 6530
rect 26256 6466 26264 6530
rect 25944 5442 26264 6466
rect 25944 5378 25952 5442
rect 26016 5378 26032 5442
rect 26096 5378 26112 5442
rect 26176 5378 26192 5442
rect 26256 5378 26264 5442
rect 25944 4354 26264 5378
rect 25944 4290 25952 4354
rect 26016 4290 26032 4354
rect 26096 4290 26112 4354
rect 26176 4290 26192 4354
rect 26256 4290 26264 4354
rect 25944 3266 26264 4290
rect 25944 3202 25952 3266
rect 26016 3202 26032 3266
rect 26096 3202 26112 3266
rect 26176 3202 26192 3266
rect 26256 3202 26264 3266
rect 25944 2178 26264 3202
rect 25944 2114 25952 2178
rect 26016 2114 26032 2178
rect 26096 2114 26112 2178
rect 26176 2114 26192 2178
rect 26256 2114 26264 2178
rect 25944 2098 26264 2114
rect 9627 1702 9693 1703
rect 9627 1638 9628 1702
rect 9692 1638 9693 1702
rect 9627 1637 9693 1638
rect 9630 1431 9690 1637
rect 9627 1430 9693 1431
rect 9627 1366 9628 1430
rect 9692 1366 9693 1430
rect 9627 1365 9693 1366
rect 9627 342 9693 343
rect 9627 278 9628 342
rect 9692 278 9693 342
rect 9627 277 9693 278
rect 9630 71 9690 277
rect 9627 70 9693 71
rect 9627 6 9628 70
rect 9692 6 9693 70
rect 9627 5 9693 6
<< via4 >>
rect 3286 11752 3522 11988
rect 24814 11752 25050 11988
<< metal5 >>
rect 3244 11988 25092 12030
rect 3244 11752 3286 11988
rect 3522 11752 24814 11988
rect 25050 11752 25092 11988
rect 3244 11710 25092 11752
use scs8hd_fill_2  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2690
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2690
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2690
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__15__A
timestamp 1586364061
transform 1 0 1932 0 1 2690
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2690
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2690
box -38 -48 314 592
use scs8hd_buf_2  _35_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2690
box -38 -48 406 592
use scs8hd_buf_2  _15_
timestamp 1586364061
transform 1 0 1380 0 1 2690
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2690
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 3956 0 1 2690
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_23 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 -1 2690
box -38 -48 774 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2690
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_32
timestamp 1586364061
transform 1 0 4048 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2690
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_44
timestamp 1586364061
transform 1 0 5152 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_56
timestamp 1586364061
transform 1 0 6256 0 1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2690
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_68
timestamp 1586364061
transform 1 0 7360 0 1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2690
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 9568 0 1 2690
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2690
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_93
timestamp 1586364061
transform 1 0 9660 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2690
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2690
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_129
timestamp 1586364061
transform 1 0 12972 0 1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2690
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 15180 0 1 2690
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2690
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_141
timestamp 1586364061
transform 1 0 14076 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_154
timestamp 1586364061
transform 1 0 15272 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_166
timestamp 1586364061
transform 1 0 16376 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2690
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2690
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_190
timestamp 1586364061
transform 1 0 18584 0 1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2690
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 20792 0 1 2690
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2690
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2690
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_245 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23644 0 1 2690
box -38 -48 130 592
use scs8hd_decap_6  FILLER_1_239
timestamp 1586364061
transform 1 0 23092 0 1 2690
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2690
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 23736 0 1 2690
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_252
timestamp 1586364061
transform 1 0 24288 0 1 2690
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_257 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24748 0 -1 2690
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_253
timestamp 1586364061
transform 1 0 24380 0 -1 2690
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__12__A
timestamp 1586364061
transform 1 0 24564 0 -1 2690
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__14__A
timestamp 1586364061
transform 1 0 24472 0 1 2690
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 23920 0 -1 2690
box -38 -48 130 592
use scs8hd_buf_2  _14_
timestamp 1586364061
transform 1 0 23920 0 1 2690
box -38 -48 406 592
use scs8hd_buf_2  _12_
timestamp 1586364061
transform 1 0 24012 0 -1 2690
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_256
timestamp 1586364061
transform 1 0 24656 0 1 2690
box -38 -48 1142 592
use scs8hd_buf_2  _16_
timestamp 1586364061
transform 1 0 25116 0 -1 2690
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 26404 0 1 2690
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__16__A
timestamp 1586364061
transform 1 0 25668 0 -1 2690
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_265
timestamp 1586364061
transform 1 0 25484 0 -1 2690
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2690
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_277
timestamp 1586364061
transform 1 0 26588 0 -1 2690
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2690
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2690
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2690
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 26772 0 -1 2690
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2690
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2690
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_288
timestamp 1586364061
transform 1 0 27600 0 1 2690
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_296
timestamp 1586364061
transform 1 0 28336 0 1 2690
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 28888 0 -1 2690
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 28888 0 1 2690
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_298
timestamp 1586364061
transform 1 0 28520 0 -1 2690
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3778
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3778
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_59
timestamp 1586364061
transform 1 0 6532 0 -1 3778
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 -1 3778
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_98
timestamp 1586364061
transform 1 0 10120 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3778
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 -1 3778
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_147
timestamp 1586364061
transform 1 0 14628 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_159
timestamp 1586364061
transform 1 0 15732 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3778
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 -1 3778
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_196
timestamp 1586364061
transform 1 0 19136 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_208
timestamp 1586364061
transform 1 0 20240 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_220
timestamp 1586364061
transform 1 0 21344 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3778
box -38 -48 1142 592
use scs8hd_buf_2  _31_
timestamp 1586364061
transform 1 0 23920 0 -1 3778
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 23552 0 -1 3778
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_245
timestamp 1586364061
transform 1 0 23644 0 -1 3778
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_252
timestamp 1586364061
transform 1 0 24288 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_264
timestamp 1586364061
transform 1 0 25392 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3778
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3778
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_296
timestamp 1586364061
transform 1 0 28336 0 -1 3778
box -38 -48 314 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 28888 0 -1 3778
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3778
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3778
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 3956 0 1 3778
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3778
box -38 -48 406 592
use scs8hd_decap_12  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_44
timestamp 1586364061
transform 1 0 5152 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3778
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 9568 0 1 3778
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_129
timestamp 1586364061
transform 1 0 12972 0 1 3778
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 15180 0 1 3778
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 15548 0 1 3778
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_141
timestamp 1586364061
transform 1 0 14076 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_154
timestamp 1586364061
transform 1 0 15272 0 1 3778
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_183
timestamp 1586364061
transform 1 0 17940 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3778
box -38 -48 1142 592
use scs8hd_buf_2  _30_
timestamp 1586364061
transform 1 0 20884 0 1 3778
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 20792 0 1 3778
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__09__A
timestamp 1586364061
transform 1 0 20424 0 1 3778
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3778
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3778
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 21436 0 1 3778
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3778
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3778
box -38 -48 1142 592
use scs8hd_buf_2  _10_
timestamp 1586364061
transform 1 0 23920 0 1 3778
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__10__A
timestamp 1586364061
transform 1 0 24472 0 1 3778
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_247
timestamp 1586364061
transform 1 0 23828 0 1 3778
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_252
timestamp 1586364061
transform 1 0 24288 0 1 3778
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_256
timestamp 1586364061
transform 1 0 24656 0 1 3778
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 26404 0 1 3778
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_268
timestamp 1586364061
transform 1 0 25760 0 1 3778
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3778
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3778
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_288
timestamp 1586364061
transform 1 0 27600 0 1 3778
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_296
timestamp 1586364061
transform 1 0 28336 0 1 3778
box -38 -48 314 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 28888 0 1 3778
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4866
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_39
timestamp 1586364061
transform 1 0 4692 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4866
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4866
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 6716 0 -1 4866
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_86
timestamp 1586364061
transform 1 0 9016 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_98
timestamp 1586364061
transform 1 0 10120 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4866
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 12328 0 -1 4866
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4866
box -38 -48 1142 592
use scs8hd_buf_2  _29_
timestamp 1586364061
transform 1 0 15548 0 -1 4866
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4866
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_155
timestamp 1586364061
transform 1 0 15364 0 -1 4866
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_161
timestamp 1586364061
transform 1 0 15916 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_173
timestamp 1586364061
transform 1 0 17020 0 -1 4866
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 17940 0 -1 4866
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4866
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_196
timestamp 1586364061
transform 1 0 19136 0 -1 4866
box -38 -48 1142 592
use scs8hd_buf_2  _09_
timestamp 1586364061
transform 1 0 20424 0 -1 4866
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4866
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_214
timestamp 1586364061
transform 1 0 20792 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4866
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 23552 0 -1 4866
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_257
timestamp 1586364061
transform 1 0 24748 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_269
timestamp 1586364061
transform 1 0 25852 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_281
timestamp 1586364061
transform 1 0 26956 0 -1 4866
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_293
timestamp 1586364061
transform 1 0 28060 0 -1 4866
box -38 -48 590 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 28888 0 -1 4866
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4866
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4866
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 3956 0 1 4866
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__07__A
timestamp 1586364061
transform 1 0 4232 0 1 4866
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4866
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4866
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_48
timestamp 1586364061
transform 1 0 5520 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4866
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 9568 0 1 4866
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4866
box -38 -48 774 592
use scs8hd_decap_12  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4866
box -38 -48 774 592
use scs8hd_buf_2  _08_
timestamp 1586364061
transform 1 0 12604 0 1 4866
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__08__A
timestamp 1586364061
transform 1 0 13156 0 1 4866
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__27__A
timestamp 1586364061
transform 1 0 13524 0 1 4866
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_129
timestamp 1586364061
transform 1 0 12972 0 1 4866
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_133
timestamp 1586364061
transform 1 0 13340 0 1 4866
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4866
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 15180 0 1 4866
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4866
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_190
timestamp 1586364061
transform 1 0 18584 0 1 4866
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 20792 0 1 4866
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_202
timestamp 1586364061
transform 1 0 19688 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4866
box -38 -48 1142 592
use scs8hd_buf_2  _28_
timestamp 1586364061
transform 1 0 23920 0 1 4866
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__28__A
timestamp 1586364061
transform 1 0 24472 0 1 4866
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_239
timestamp 1586364061
transform 1 0 23092 0 1 4866
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_247
timestamp 1586364061
transform 1 0 23828 0 1 4866
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_252
timestamp 1586364061
transform 1 0 24288 0 1 4866
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_256
timestamp 1586364061
transform 1 0 24656 0 1 4866
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 26404 0 1 4866
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_268
timestamp 1586364061
transform 1 0 25760 0 1 4866
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_274
timestamp 1586364061
transform 1 0 26312 0 1 4866
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4866
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_288
timestamp 1586364061
transform 1 0 27600 0 1 4866
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_296
timestamp 1586364061
transform 1 0 28336 0 1 4866
box -38 -48 314 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 28888 0 1 4866
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5954
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5954
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5954
box -38 -48 1142 592
use scs8hd_buf_2  _07_
timestamp 1586364061
transform 1 0 4140 0 -1 5954
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 3956 0 1 5954
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5954
box -38 -48 590 592
use scs8hd_decap_12  FILLER_6_37
timestamp 1586364061
transform 1 0 4508 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5954
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_44
timestamp 1586364061
transform 1 0 5152 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5954
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 6716 0 -1 5954
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_74
timestamp 1586364061
transform 1 0 7912 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_68
timestamp 1586364061
transform 1 0 7360 0 1 5954
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 9568 0 1 5954
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_98
timestamp 1586364061
transform 1 0 10120 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_93
timestamp 1586364061
transform 1 0 9660 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5954
box -38 -48 1142 592
use scs8hd_buf_2  _27_
timestamp 1586364061
transform 1 0 12880 0 -1 5954
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 12328 0 -1 5954
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5954
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5954
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_129
timestamp 1586364061
transform 1 0 12972 0 1 5954
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 15180 0 1 5954
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__06__A
timestamp 1586364061
transform 1 0 14720 0 1 5954
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_156
timestamp 1586364061
transform 1 0 15456 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_141
timestamp 1586364061
transform 1 0 14076 0 1 5954
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5954
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5954
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_154
timestamp 1586364061
transform 1 0 15272 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5954
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 17940 0 -1 5954
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5954
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_196
timestamp 1586364061
transform 1 0 19136 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_190
timestamp 1586364061
transform 1 0 18584 0 1 5954
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 20792 0 1 5954
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_208
timestamp 1586364061
transform 1 0 20240 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_202
timestamp 1586364061
transform 1 0 19688 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_215
timestamp 1586364061
transform 1 0 20884 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_220
timestamp 1586364061
transform 1 0 21344 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_227
timestamp 1586364061
transform 1 0 21988 0 1 5954
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 23552 0 -1 5954
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__25__A
timestamp 1586364061
transform 1 0 23920 0 1 5954
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_245
timestamp 1586364061
transform 1 0 23644 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_257
timestamp 1586364061
transform 1 0 24748 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5954
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_247
timestamp 1586364061
transform 1 0 23828 0 1 5954
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_250
timestamp 1586364061
transform 1 0 24104 0 1 5954
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 26404 0 1 5954
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_269
timestamp 1586364061
transform 1 0 25852 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_262
timestamp 1586364061
transform 1 0 25208 0 1 5954
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_274
timestamp 1586364061
transform 1 0 26312 0 1 5954
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5954
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_281
timestamp 1586364061
transform 1 0 26956 0 -1 5954
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_6_293
timestamp 1586364061
transform 1 0 28060 0 -1 5954
box -38 -48 590 592
use scs8hd_decap_8  FILLER_7_288
timestamp 1586364061
transform 1 0 27600 0 1 5954
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_296
timestamp 1586364061
transform 1 0 28336 0 1 5954
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 28888 0 -1 5954
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 28888 0 1 5954
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7042
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7042
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_59
timestamp 1586364061
transform 1 0 6532 0 -1 7042
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 6716 0 -1 7042
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_98
timestamp 1586364061
transform 1 0 10120 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_110
timestamp 1586364061
transform 1 0 11224 0 -1 7042
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 12328 0 -1 7042
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7042
box -38 -48 1142 592
use scs8hd_buf_2  _06_
timestamp 1586364061
transform 1 0 14720 0 -1 7042
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_147
timestamp 1586364061
transform 1 0 14628 0 -1 7042
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_176
timestamp 1586364061
transform 1 0 17296 0 -1 7042
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 17940 0 -1 7042
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7042
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_184
timestamp 1586364061
transform 1 0 18032 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_220
timestamp 1586364061
transform 1 0 21344 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7042
box -38 -48 1142 592
use scs8hd_buf_2  _25_
timestamp 1586364061
transform 1 0 23920 0 -1 7042
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 23552 0 -1 7042
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7042
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_252
timestamp 1586364061
transform 1 0 24288 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_264
timestamp 1586364061
transform 1 0 25392 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7042
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7042
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_296
timestamp 1586364061
transform 1 0 28336 0 -1 7042
box -38 -48 314 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 28888 0 -1 7042
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7042
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7042
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 1 7042
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7042
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_68
timestamp 1586364061
transform 1 0 7360 0 1 7042
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 1 7042
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_80
timestamp 1586364061
transform 1 0 8464 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_93
timestamp 1586364061
transform 1 0 9660 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7042
box -38 -48 1142 592
use scs8hd_buf_2  _05_
timestamp 1586364061
transform 1 0 13064 0 1 7042
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__05__A
timestamp 1586364061
transform 1 0 13616 0 1 7042
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_129
timestamp 1586364061
transform 1 0 12972 0 1 7042
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7042
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7042
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 1 7042
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_150
timestamp 1586364061
transform 1 0 14904 0 1 7042
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7042
box -38 -48 774 592
use scs8hd_buf_2  _04_
timestamp 1586364061
transform 1 0 18400 0 1 7042
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__04__A
timestamp 1586364061
transform 1 0 18952 0 1 7042
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_186
timestamp 1586364061
transform 1 0 18216 0 1 7042
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_192
timestamp 1586364061
transform 1 0 18768 0 1 7042
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7042
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 1 7042
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7042
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7042
box -38 -48 1142 592
use scs8hd_buf_2  _24_
timestamp 1586364061
transform 1 0 22264 0 1 7042
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__24__A
timestamp 1586364061
transform 1 0 22816 0 1 7042
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_227
timestamp 1586364061
transform 1 0 21988 0 1 7042
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7042
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_238
timestamp 1586364061
transform 1 0 23000 0 1 7042
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__03__A
timestamp 1586364061
transform 1 0 23920 0 1 7042
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_246
timestamp 1586364061
transform 1 0 23736 0 1 7042
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_250
timestamp 1586364061
transform 1 0 24104 0 1 7042
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 26404 0 1 7042
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7042
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7042
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7042
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_288
timestamp 1586364061
transform 1 0 27600 0 1 7042
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_296
timestamp 1586364061
transform 1 0 28336 0 1 7042
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 28888 0 1 7042
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8130
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8130
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8130
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 6716 0 -1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_86
timestamp 1586364061
transform 1 0 9016 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8130
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 12328 0 -1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_135
timestamp 1586364061
transform 1 0 13524 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_159
timestamp 1586364061
transform 1 0 15732 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8130
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 17940 0 -1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_184
timestamp 1586364061
transform 1 0 18032 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_220
timestamp 1586364061
transform 1 0 21344 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 8130
box -38 -48 1142 592
use scs8hd_buf_2  _03_
timestamp 1586364061
transform 1 0 23920 0 -1 8130
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 23552 0 -1 8130
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 8130
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_252
timestamp 1586364061
transform 1 0 24288 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_264
timestamp 1586364061
transform 1 0 25392 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8130
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8130
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_296
timestamp 1586364061
transform 1 0 28336 0 -1 8130
box -38 -48 314 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 28888 0 -1 8130
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8130
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 1564 0 1 8130
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8130
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8130
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_44
timestamp 1586364061
transform 1 0 5152 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_68
timestamp 1586364061
transform 1 0 7360 0 1 8130
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_129
timestamp 1586364061
transform 1 0 12972 0 1 8130
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_141
timestamp 1586364061
transform 1 0 14076 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_166
timestamp 1586364061
transform 1 0 16376 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_190
timestamp 1586364061
transform 1 0 18584 0 1 8130
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_202
timestamp 1586364061
transform 1 0 19688 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_215
timestamp 1586364061
transform 1 0 20884 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8130
box -38 -48 1142 592
use scs8hd_buf_2  _23_
timestamp 1586364061
transform 1 0 23920 0 1 8130
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__02__A
timestamp 1586364061
transform 1 0 24472 0 1 8130
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__23__A
timestamp 1586364061
transform 1 0 23736 0 1 8130
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_239
timestamp 1586364061
transform 1 0 23092 0 1 8130
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8130
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_252
timestamp 1586364061
transform 1 0 24288 0 1 8130
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_256
timestamp 1586364061
transform 1 0 24656 0 1 8130
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 1 8130
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8130
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8130
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8130
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_288
timestamp 1586364061
transform 1 0 27600 0 1 8130
box -38 -48 774 592
use scs8hd_decap_3  FILLER_11_296
timestamp 1586364061
transform 1 0 28336 0 1 8130
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 28888 0 1 8130
box -38 -48 314 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 1380 0 -1 9218
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9218
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_31
timestamp 1586364061
transform 1 0 3956 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_43
timestamp 1586364061
transform 1 0 5060 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9218
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6716 0 -1 9218
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_98
timestamp 1586364061
transform 1 0 10120 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9218
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 12328 0 -1 9218
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_123
timestamp 1586364061
transform 1 0 12420 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_159
timestamp 1586364061
transform 1 0 15732 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_171
timestamp 1586364061
transform 1 0 16836 0 -1 9218
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 17940 0 -1 9218
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_196
timestamp 1586364061
transform 1 0 19136 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_208
timestamp 1586364061
transform 1 0 20240 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_220
timestamp 1586364061
transform 1 0 21344 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_232
timestamp 1586364061
transform 1 0 22448 0 -1 9218
box -38 -48 1142 592
use scs8hd_buf_2  _02_
timestamp 1586364061
transform 1 0 23920 0 -1 9218
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 23552 0 -1 9218
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_245
timestamp 1586364061
transform 1 0 23644 0 -1 9218
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_252
timestamp 1586364061
transform 1 0 24288 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_264
timestamp 1586364061
transform 1 0 25392 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9218
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9218
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_296
timestamp 1586364061
transform 1 0 28336 0 -1 9218
box -38 -48 314 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 28888 0 -1 9218
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9218
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__20__A
timestamp 1586364061
transform 1 0 1932 0 1 9218
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10306
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9218
box -38 -48 314 592
use scs8hd_buf_2  _34_
timestamp 1586364061
transform 1 0 1380 0 1 9218
box -38 -48 406 592
use scs8hd_buf_2  _20_
timestamp 1586364061
transform 1 0 1380 0 -1 10306
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9218
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 2300 0 1 9218
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9218
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 3956 0 1 9218
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9218
box -38 -48 406 592
use scs8hd_decap_12  FILLER_13_32
timestamp 1586364061
transform 1 0 4048 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_31
timestamp 1586364061
transform 1 0 3956 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_55
timestamp 1586364061
transform 1 0 6164 0 -1 10306
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 6716 0 -1 10306
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7912 0 -1 10306
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8280 0 -1 10306
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_68
timestamp 1586364061
transform 1 0 7360 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10306
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10306
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 9568 0 1 9218
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_92
timestamp 1586364061
transform 1 0 9568 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10306
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 12328 0 -1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_123
timestamp 1586364061
transform 1 0 12420 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 15180 0 1 9218
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_159
timestamp 1586364061
transform 1 0 15732 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 17940 0 -1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_190
timestamp 1586364061
transform 1 0 18584 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_184
timestamp 1586364061
transform 1 0 18032 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 20792 0 1 9218
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_215
timestamp 1586364061
transform 1 0 20884 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_208
timestamp 1586364061
transform 1 0 20240 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_220
timestamp 1586364061
transform 1 0 21344 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10306
box -38 -48 1142 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 23920 0 1 9218
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 23552 0 -1 10306
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 24472 0 1 9218
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9218
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_247
timestamp 1586364061
transform 1 0 23828 0 1 9218
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_252
timestamp 1586364061
transform 1 0 24288 0 1 9218
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_256
timestamp 1586364061
transform 1 0 24656 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_245
timestamp 1586364061
transform 1 0 23644 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_257
timestamp 1586364061
transform 1 0 24748 0 -1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 26404 0 1 9218
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_268
timestamp 1586364061
transform 1 0 25760 0 1 9218
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_274
timestamp 1586364061
transform 1 0 26312 0 1 9218
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9218
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_269
timestamp 1586364061
transform 1 0 25852 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_288
timestamp 1586364061
transform 1 0 27600 0 1 9218
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_296
timestamp 1586364061
transform 1 0 28336 0 1 9218
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_281
timestamp 1586364061
transform 1 0 26956 0 -1 10306
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_293
timestamp 1586364061
transform 1 0 28060 0 -1 10306
box -38 -48 590 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 28888 0 1 9218
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 28888 0 -1 10306
box -38 -48 314 592
use scs8hd_buf_2  _32_
timestamp 1586364061
transform 1 0 1380 0 1 10306
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10306
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 1932 0 1 10306
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 2300 0 1 10306
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10306
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10306
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 1 10306
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10306
box -38 -48 406 592
use scs8hd_decap_12  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10306
box -38 -48 774 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7912 0 1 10306
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7728 0 1 10306
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7360 0 1 10306
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 1 10306
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10306
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_70
timestamp 1586364061
transform 1 0 7544 0 1 10306
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 1 10306
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8924 0 1 10306
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10306
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10306
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_129
timestamp 1586364061
transform 1 0 12972 0 1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 15180 0 1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_141
timestamp 1586364061
transform 1 0 14076 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_190
timestamp 1586364061
transform 1 0 18584 0 1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 20792 0 1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_215
timestamp 1586364061
transform 1 0 20884 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10306
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 23920 0 1 10306
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_239
timestamp 1586364061
transform 1 0 23092 0 1 10306
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_247
timestamp 1586364061
transform 1 0 23828 0 1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_250
timestamp 1586364061
transform 1 0 24104 0 1 10306
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 26404 0 1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_262
timestamp 1586364061
transform 1 0 25208 0 1 10306
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_15_274
timestamp 1586364061
transform 1 0 26312 0 1 10306
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10306
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_288
timestamp 1586364061
transform 1 0 27600 0 1 10306
box -38 -48 774 592
use scs8hd_decap_3  FILLER_15_296
timestamp 1586364061
transform 1 0 28336 0 1 10306
box -38 -48 314 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 28888 0 1 10306
box -38 -48 314 592
use scs8hd_buf_2  _33_
timestamp 1586364061
transform 1 0 1380 0 -1 11394
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11394
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_31
timestamp 1586364061
transform 1 0 3956 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_55
timestamp 1586364061
transform 1 0 6164 0 -1 11394
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7728 0 -1 11394
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 -1 11394
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11394
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11394
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11394
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 -1 11394
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 12144 0 -1 11394
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_123
timestamp 1586364061
transform 1 0 12420 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_147
timestamp 1586364061
transform 1 0 14628 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_159
timestamp 1586364061
transform 1 0 15732 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11394
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 -1 11394
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_184
timestamp 1586364061
transform 1 0 18032 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_196
timestamp 1586364061
transform 1 0 19136 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_208
timestamp 1586364061
transform 1 0 20240 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_220
timestamp 1586364061
transform 1 0 21344 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_232
timestamp 1586364061
transform 1 0 22448 0 -1 11394
box -38 -48 1142 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 23920 0 -1 11394
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 23552 0 -1 11394
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_245
timestamp 1586364061
transform 1 0 23644 0 -1 11394
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_252
timestamp 1586364061
transform 1 0 24288 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_264
timestamp 1586364061
transform 1 0 25392 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11394
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_288
timestamp 1586364061
transform 1 0 27600 0 -1 11394
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_296
timestamp 1586364061
transform 1 0 28336 0 -1 11394
box -38 -48 314 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 28888 0 -1 11394
box -38 -48 314 592
use scs8hd_buf_2  _13_
timestamp 1586364061
transform 1 0 1380 0 1 11394
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11394
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__13__A
timestamp 1586364061
transform 1 0 1932 0 1 11394
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11394
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11394
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 3956 0 1 11394
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11394
box -38 -48 774 592
use scs8hd_decap_12  FILLER_17_32
timestamp 1586364061
transform 1 0 4048 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11394
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7912 0 1 11394
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8280 0 1 11394
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11394
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_76
timestamp 1586364061
transform 1 0 8096 0 1 11394
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 9568 0 1 11394
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8648 0 1 11394
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11394
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_84
timestamp 1586364061
transform 1 0 8832 0 1 11394
box -38 -48 774 592
use scs8hd_decap_12  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11394
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 11960 0 1 11394
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11394
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11394
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 12144 0 1 11394
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13156 0 1 11394
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13524 0 1 11394
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_129
timestamp 1586364061
transform 1 0 12972 0 1 11394
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_133
timestamp 1586364061
transform 1 0 13340 0 1 11394
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11394
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 15180 0 1 11394
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 13892 0 1 11394
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_154
timestamp 1586364061
transform 1 0 15272 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_190
timestamp 1586364061
transform 1 0 18584 0 1 11394
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 20792 0 1 11394
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_202
timestamp 1586364061
transform 1 0 19688 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_227
timestamp 1586364061
transform 1 0 21988 0 1 11394
box -38 -48 1142 592
use scs8hd_buf_2  _19_
timestamp 1586364061
transform 1 0 23920 0 1 11394
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__19__A
timestamp 1586364061
transform 1 0 24472 0 1 11394
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11394
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_247
timestamp 1586364061
transform 1 0 23828 0 1 11394
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_252
timestamp 1586364061
transform 1 0 24288 0 1 11394
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_256
timestamp 1586364061
transform 1 0 24656 0 1 11394
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 26404 0 1 11394
box -38 -48 130 592
use scs8hd_decap_6  FILLER_17_268
timestamp 1586364061
transform 1 0 25760 0 1 11394
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11394
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11394
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_288
timestamp 1586364061
transform 1 0 27600 0 1 11394
box -38 -48 774 592
use scs8hd_decap_3  FILLER_17_296
timestamp 1586364061
transform 1 0 28336 0 1 11394
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 28888 0 1 11394
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12482
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__26__A
timestamp 1586364061
transform 1 0 1564 0 -1 12482
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12482
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_31
timestamp 1586364061
transform 1 0 3956 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_55
timestamp 1586364061
transform 1 0 6164 0 -1 12482
box -38 -48 590 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 12482
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 -1 12482
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_95
timestamp 1586364061
transform 1 0 9844 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12482
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12482
box -38 -48 130 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13064 0 -1 12482
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 -1 12482
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 12144 0 -1 12482
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12482
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12482
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_139
timestamp 1586364061
transform 1 0 13892 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12482
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 17940 0 -1 12482
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_196
timestamp 1586364061
transform 1 0 19136 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_208
timestamp 1586364061
transform 1 0 20240 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_220
timestamp 1586364061
transform 1 0 21344 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_232
timestamp 1586364061
transform 1 0 22448 0 -1 12482
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 23552 0 -1 12482
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_245
timestamp 1586364061
transform 1 0 23644 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_257
timestamp 1586364061
transform 1 0 24748 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_269
timestamp 1586364061
transform 1 0 25852 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_281
timestamp 1586364061
transform 1 0 26956 0 -1 12482
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_293
timestamp 1586364061
transform 1 0 28060 0 -1 12482
box -38 -48 590 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 28888 0 -1 12482
box -38 -48 314 592
use scs8hd_buf_2  _11_
timestamp 1586364061
transform 1 0 1380 0 1 12482
box -38 -48 406 592
use scs8hd_buf_2  _26_
timestamp 1586364061
transform 1 0 1380 0 -1 13570
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12482
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13570
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__11__A
timestamp 1586364061
transform 1 0 1932 0 1 12482
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12482
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 3956 0 1 12482
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12482
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_31
timestamp 1586364061
transform 1 0 3956 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_44
timestamp 1586364061
transform 1 0 5152 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13570
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 6716 0 -1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_68
timestamp 1586364061
transform 1 0 7360 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 9568 0 1 12482
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_80
timestamp 1586364061
transform 1 0 8464 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_98
timestamp 1586364061
transform 1 0 10120 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_110
timestamp 1586364061
transform 1 0 11224 0 -1 13570
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13524 0 -1 13570
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 12328 0 -1 13570
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13524 0 1 12482
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_129
timestamp 1586364061
transform 1 0 12972 0 1 12482
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12482
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 15180 0 1 12482
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 1 12482
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14260 0 1 12482
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_141
timestamp 1586364061
transform 1 0 14076 0 1 12482
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_145
timestamp 1586364061
transform 1 0 14444 0 1 12482
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_166
timestamp 1586364061
transform 1 0 16376 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_178
timestamp 1586364061
transform 1 0 17480 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13570
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1586364061
transform 1 0 19136 0 -1 13570
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 17940 0 -1 13570
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1586364061
transform 1 0 19136 0 1 12482
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_190
timestamp 1586364061
transform 1 0 18584 0 1 12482
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_198
timestamp 1586364061
transform 1 0 19320 0 1 12482
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13570
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_184
timestamp 1586364061
transform 1 0 18032 0 -1 13570
box -38 -48 1142 592
use scs8hd_conb_1  _01_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 1 12482
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 20792 0 1 12482
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1586364061
transform 1 0 19504 0 1 12482
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1586364061
transform 1 0 19872 0 1 12482
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_202
timestamp 1586364061
transform 1 0 19688 0 1 12482
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_206
timestamp 1586364061
transform 1 0 20056 0 1 12482
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_218
timestamp 1586364061
transform 1 0 21160 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_205
timestamp 1586364061
transform 1 0 19964 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_217
timestamp 1586364061
transform 1 0 21068 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_229
timestamp 1586364061
transform 1 0 22172 0 -1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 23552 0 -1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_242
timestamp 1586364061
transform 1 0 23368 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_241
timestamp 1586364061
transform 1 0 23276 0 -1 13570
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_245
timestamp 1586364061
transform 1 0 23644 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_257
timestamp 1586364061
transform 1 0 24748 0 -1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 26404 0 1 12482
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_266
timestamp 1586364061
transform 1 0 25576 0 1 12482
box -38 -48 774 592
use scs8hd_fill_1  FILLER_19_274
timestamp 1586364061
transform 1 0 26312 0 1 12482
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_276
timestamp 1586364061
transform 1 0 26496 0 1 12482
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_269
timestamp 1586364061
transform 1 0 25852 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_288
timestamp 1586364061
transform 1 0 27600 0 1 12482
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_296
timestamp 1586364061
transform 1 0 28336 0 1 12482
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_281
timestamp 1586364061
transform 1 0 26956 0 -1 13570
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_293
timestamp 1586364061
transform 1 0 28060 0 -1 13570
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 28888 0 1 12482
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 28888 0 -1 13570
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13570
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 3956 0 1 13570
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13570
box -38 -48 406 592
use scs8hd_decap_12  FILLER_21_32
timestamp 1586364061
transform 1 0 4048 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_56
timestamp 1586364061
transform 1 0 6256 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_68
timestamp 1586364061
transform 1 0 7360 0 1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 9568 0 1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_105
timestamp 1586364061
transform 1 0 10764 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_117
timestamp 1586364061
transform 1 0 11868 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_129
timestamp 1586364061
transform 1 0 12972 0 1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 15180 0 1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_166
timestamp 1586364061
transform 1 0 16376 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_190
timestamp 1586364061
transform 1 0 18584 0 1 13570
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_198
timestamp 1586364061
transform 1 0 19320 0 1 13570
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 20792 0 1 13570
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1586364061
transform 1 0 19412 0 1 13570
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1586364061
transform 1 0 19780 0 1 13570
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1586364061
transform 1 0 20148 0 1 13570
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_201
timestamp 1586364061
transform 1 0 19596 0 1 13570
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_205
timestamp 1586364061
transform 1 0 19964 0 1 13570
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_209
timestamp 1586364061
transform 1 0 20332 0 1 13570
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_215
timestamp 1586364061
transform 1 0 20884 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_227
timestamp 1586364061
transform 1 0 21988 0 1 13570
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__22__A
timestamp 1586364061
transform 1 0 23920 0 1 13570
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_239
timestamp 1586364061
transform 1 0 23092 0 1 13570
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_247
timestamp 1586364061
transform 1 0 23828 0 1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_250
timestamp 1586364061
transform 1 0 24104 0 1 13570
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 26404 0 1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_262
timestamp 1586364061
transform 1 0 25208 0 1 13570
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_21_274
timestamp 1586364061
transform 1 0 26312 0 1 13570
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13570
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_288
timestamp 1586364061
transform 1 0 27600 0 1 13570
box -38 -48 774 592
use scs8hd_decap_3  FILLER_21_296
timestamp 1586364061
transform 1 0 28336 0 1 13570
box -38 -48 314 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 28888 0 1 13570
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14658
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_39
timestamp 1586364061
transform 1 0 4692 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14658
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_59
timestamp 1586364061
transform 1 0 6532 0 -1 14658
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 6716 0 -1 14658
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_62
timestamp 1586364061
transform 1 0 6808 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_74
timestamp 1586364061
transform 1 0 7912 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_86
timestamp 1586364061
transform 1 0 9016 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_98
timestamp 1586364061
transform 1 0 10120 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14658
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 12328 0 -1 14658
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_135
timestamp 1586364061
transform 1 0 13524 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_147
timestamp 1586364061
transform 1 0 14628 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_159
timestamp 1586364061
transform 1 0 15732 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_171
timestamp 1586364061
transform 1 0 16836 0 -1 14658
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 17940 0 -1 14658
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1586364061
transform 1 0 18952 0 -1 14658
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_184
timestamp 1586364061
transform 1 0 18032 0 -1 14658
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_192
timestamp 1586364061
transform 1 0 18768 0 -1 14658
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14658
box -38 -48 314 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1586364061
transform 1 0 19412 0 -1 14658
box -38 -48 866 592
use scs8hd_decap_12  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_220
timestamp 1586364061
transform 1 0 21344 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_232
timestamp 1586364061
transform 1 0 22448 0 -1 14658
box -38 -48 1142 592
use scs8hd_buf_2  _22_
timestamp 1586364061
transform 1 0 23920 0 -1 14658
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 23552 0 -1 14658
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_245
timestamp 1586364061
transform 1 0 23644 0 -1 14658
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_264
timestamp 1586364061
transform 1 0 25392 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14658
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_288
timestamp 1586364061
transform 1 0 27600 0 -1 14658
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_296
timestamp 1586364061
transform 1 0 28336 0 -1 14658
box -38 -48 314 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 28888 0 -1 14658
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14658
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14658
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 1 14658
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14658
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_44
timestamp 1586364061
transform 1 0 5152 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_68
timestamp 1586364061
transform 1 0 7360 0 1 14658
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 1 14658
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_129
timestamp 1586364061
transform 1 0 12972 0 1 14658
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 1 14658
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_178
timestamp 1586364061
transform 1 0 17480 0 1 14658
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1586364061
transform 1 0 18952 0 1 14658
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1586364061
transform 1 0 18768 0 1 14658
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_190
timestamp 1586364061
transform 1 0 18584 0 1 14658
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 1 14658
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_203
timestamp 1586364061
transform 1 0 19780 0 1 14658
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_211
timestamp 1586364061
transform 1 0 20516 0 1 14658
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_215
timestamp 1586364061
transform 1 0 20884 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_227
timestamp 1586364061
transform 1 0 21988 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_239
timestamp 1586364061
transform 1 0 23092 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_251
timestamp 1586364061
transform 1 0 24196 0 1 14658
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 26404 0 1 14658
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14658
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_288
timestamp 1586364061
transform 1 0 27600 0 1 14658
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_296
timestamp 1586364061
transform 1 0 28336 0 1 14658
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 28888 0 1 14658
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15746
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_39
timestamp 1586364061
transform 1 0 4692 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15746
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15746
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 6716 0 -1 15746
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7084 0 -1 15746
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15746
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_103
timestamp 1586364061
transform 1 0 10580 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15746
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 12328 0 -1 15746
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15746
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_147
timestamp 1586364061
transform 1 0 14628 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_159
timestamp 1586364061
transform 1 0 15732 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_171
timestamp 1586364061
transform 1 0 16836 0 -1 15746
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 17940 0 -1 15746
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1586364061
transform 1 0 18952 0 -1 15746
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_184
timestamp 1586364061
transform 1 0 18032 0 -1 15746
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15746
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_196
timestamp 1586364061
transform 1 0 19136 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_208
timestamp 1586364061
transform 1 0 20240 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_220
timestamp 1586364061
transform 1 0 21344 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_232
timestamp 1586364061
transform 1 0 22448 0 -1 15746
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 23552 0 -1 15746
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_245
timestamp 1586364061
transform 1 0 23644 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_257
timestamp 1586364061
transform 1 0 24748 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_269
timestamp 1586364061
transform 1 0 25852 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_281
timestamp 1586364061
transform 1 0 26956 0 -1 15746
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_293
timestamp 1586364061
transform 1 0 28060 0 -1 15746
box -38 -48 590 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 28888 0 -1 15746
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15746
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15746
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 3956 0 1 15746
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15746
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_32
timestamp 1586364061
transform 1 0 4048 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_44
timestamp 1586364061
transform 1 0 5152 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15746
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_1_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 1 15746
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6900 0 1 15746
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15746
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 9568 0 1 15746
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_84
timestamp 1586364061
transform 1 0 8832 0 1 15746
box -38 -48 774 592
use scs8hd_decap_12  FILLER_25_93
timestamp 1586364061
transform 1 0 9660 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_105
timestamp 1586364061
transform 1 0 10764 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15746
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 13064 0 1 15746
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 13432 0 1 15746
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_129
timestamp 1586364061
transform 1 0 12972 0 1 15746
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15746
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15746
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 15180 0 1 15746
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_148
timestamp 1586364061
transform 1 0 14720 0 1 15746
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15746
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_190
timestamp 1586364061
transform 1 0 18584 0 1 15746
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 20792 0 1 15746
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_202
timestamp 1586364061
transform 1 0 19688 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_227
timestamp 1586364061
transform 1 0 21988 0 1 15746
box -38 -48 1142 592
use scs8hd_buf_2  _21_
timestamp 1586364061
transform 1 0 23920 0 1 15746
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__21__A
timestamp 1586364061
transform 1 0 24472 0 1 15746
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_239
timestamp 1586364061
transform 1 0 23092 0 1 15746
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_247
timestamp 1586364061
transform 1 0 23828 0 1 15746
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_252
timestamp 1586364061
transform 1 0 24288 0 1 15746
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_256
timestamp 1586364061
transform 1 0 24656 0 1 15746
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 26404 0 1 15746
box -38 -48 130 592
use scs8hd_decap_6  FILLER_25_268
timestamp 1586364061
transform 1 0 25760 0 1 15746
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15746
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15746
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_288
timestamp 1586364061
transform 1 0 27600 0 1 15746
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_296
timestamp 1586364061
transform 1 0 28336 0 1 15746
box -38 -48 314 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 28888 0 1 15746
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16834
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16834
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16834
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_39
timestamp 1586364061
transform 1 0 4692 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16834
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16834
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_59
timestamp 1586364061
transform 1 0 6532 0 -1 16834
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16834
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 -1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_62
timestamp 1586364061
transform 1 0 6808 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_68
timestamp 1586364061
transform 1 0 7360 0 1 16834
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 9568 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_98
timestamp 1586364061
transform 1 0 10120 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16834
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 13064 0 -1 16834
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 -1 16834
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16834
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_129
timestamp 1586364061
transform 1 0 12972 0 1 16834
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 15180 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_141
timestamp 1586364061
transform 1 0 14076 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16834
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1586364061
transform 1 0 17480 0 1 16834
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_173
timestamp 1586364061
transform 1 0 17020 0 -1 16834
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_166
timestamp 1586364061
transform 1 0 16376 0 1 16834
box -38 -48 1142 592
use scs8hd_mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 16834
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 17940 0 -1 16834
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1586364061
transform 1 0 17848 0 1 16834
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 -1 16834
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_181
timestamp 1586364061
transform 1 0 17756 0 -1 16834
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16834
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16834
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16834
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16834
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 20792 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_200
timestamp 1586364061
transform 1 0 19504 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16834
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_213
timestamp 1586364061
transform 1 0 20700 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_215
timestamp 1586364061
transform 1 0 20884 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_236
timestamp 1586364061
transform 1 0 22816 0 -1 16834
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16834
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 23552 0 -1 16834
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 23920 0 1 16834
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_245
timestamp 1586364061
transform 1 0 23644 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_257
timestamp 1586364061
transform 1 0 24748 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_239
timestamp 1586364061
transform 1 0 23092 0 1 16834
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_247
timestamp 1586364061
transform 1 0 23828 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_250
timestamp 1586364061
transform 1 0 24104 0 1 16834
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 26404 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_269
timestamp 1586364061
transform 1 0 25852 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_262
timestamp 1586364061
transform 1 0 25208 0 1 16834
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_274
timestamp 1586364061
transform 1 0 26312 0 1 16834
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16834
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_281
timestamp 1586364061
transform 1 0 26956 0 -1 16834
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_293
timestamp 1586364061
transform 1 0 28060 0 -1 16834
box -38 -48 590 592
use scs8hd_decap_8  FILLER_27_288
timestamp 1586364061
transform 1 0 27600 0 1 16834
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_296
timestamp 1586364061
transform 1 0 28336 0 1 16834
box -38 -48 314 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 28888 0 -1 16834
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 28888 0 1 16834
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17922
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17922
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17922
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 6716 0 -1 17922
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_62
timestamp 1586364061
transform 1 0 6808 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_98
timestamp 1586364061
transform 1 0 10120 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17922
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 12328 0 -1 17922
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_123
timestamp 1586364061
transform 1 0 12420 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_147
timestamp 1586364061
transform 1 0 14628 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_159
timestamp 1586364061
transform 1 0 15732 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_171
timestamp 1586364061
transform 1 0 16836 0 -1 17922
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 17940 0 -1 17922
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_208
timestamp 1586364061
transform 1 0 20240 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_220
timestamp 1586364061
transform 1 0 21344 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_232
timestamp 1586364061
transform 1 0 22448 0 -1 17922
box -38 -48 1142 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 23920 0 -1 17922
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 23552 0 -1 17922
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_245
timestamp 1586364061
transform 1 0 23644 0 -1 17922
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_252
timestamp 1586364061
transform 1 0 24288 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_264
timestamp 1586364061
transform 1 0 25392 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17922
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_288
timestamp 1586364061
transform 1 0 27600 0 -1 17922
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_296
timestamp 1586364061
transform 1 0 28336 0 -1 17922
box -38 -48 314 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 28888 0 -1 17922
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17922
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17922
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 3956 0 1 17922
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17922
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_56
timestamp 1586364061
transform 1 0 6256 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_68
timestamp 1586364061
transform 1 0 7360 0 1 17922
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 9568 0 1 17922
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8556 0 1 17922
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8924 0 1 17922
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17922
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17922
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_87
timestamp 1586364061
transform 1 0 9108 0 1 17922
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17922
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_129
timestamp 1586364061
transform 1 0 12972 0 1 17922
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 15180 0 1 17922
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__CLK
timestamp 1586364061
transform 1 0 15456 0 1 17922
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17922
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_154
timestamp 1586364061
transform 1 0 15272 0 1 17922
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_158
timestamp 1586364061
transform 1 0 15640 0 1 17922
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.scs8hd_dfxbp_1_3__D
timestamp 1586364061
transform 1 0 15824 0 1 17922
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_162
timestamp 1586364061
transform 1 0 16008 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_186
timestamp 1586364061
transform 1 0 18216 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_198
timestamp 1586364061
transform 1 0 19320 0 1 17922
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 20792 0 1 17922
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20608 0 1 17922
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_210
timestamp 1586364061
transform 1 0 20424 0 1 17922
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_215
timestamp 1586364061
transform 1 0 20884 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_227
timestamp 1586364061
transform 1 0 21988 0 1 17922
box -38 -48 1142 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 23920 0 1 17922
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 24472 0 1 17922
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 23736 0 1 17922
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_239
timestamp 1586364061
transform 1 0 23092 0 1 17922
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17922
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_252
timestamp 1586364061
transform 1 0 24288 0 1 17922
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_256
timestamp 1586364061
transform 1 0 24656 0 1 17922
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 26404 0 1 17922
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__18__A
timestamp 1586364061
transform 1 0 25024 0 1 17922
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_262
timestamp 1586364061
transform 1 0 25208 0 1 17922
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17922
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_276
timestamp 1586364061
transform 1 0 26496 0 1 17922
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_288
timestamp 1586364061
transform 1 0 27600 0 1 17922
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_296
timestamp 1586364061
transform 1 0 28336 0 1 17922
box -38 -48 314 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 28888 0 1 17922
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19010
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_51
timestamp 1586364061
transform 1 0 5796 0 -1 19010
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19010
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 6716 0 -1 19010
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_62
timestamp 1586364061
transform 1 0 6808 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_74
timestamp 1586364061
transform 1 0 7912 0 -1 19010
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8556 0 -1 19010
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19010
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_100
timestamp 1586364061
transform 1 0 10304 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_112
timestamp 1586364061
transform 1 0 11408 0 -1 19010
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 12328 0 -1 19010
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_120
timestamp 1586364061
transform 1 0 12144 0 -1 19010
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_123
timestamp 1586364061
transform 1 0 12420 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19010
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_ipin_0.scs8hd_dfxbp_1_3_
timestamp 1586364061
transform 1 0 15364 0 -1 19010
box -38 -48 1786 592
use scs8hd_decap_8  FILLER_30_147
timestamp 1586364061
transform 1 0 14628 0 -1 19010
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_174
timestamp 1586364061
transform 1 0 17112 0 -1 19010
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 17940 0 -1 19010
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_182
timestamp 1586364061
transform 1 0 17848 0 -1 19010
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_184
timestamp 1586364061
transform 1 0 18032 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_196
timestamp 1586364061
transform 1 0 19136 0 -1 19010
box -38 -48 1142 592
use scs8hd_buf_1  mux_bottom_ipin_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20608 0 -1 19010
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_208
timestamp 1586364061
transform 1 0 20240 0 -1 19010
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19010
box -38 -48 1142 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 23920 0 -1 19010
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 23552 0 -1 19010
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19010
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_243
timestamp 1586364061
transform 1 0 23460 0 -1 19010
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_245
timestamp 1586364061
transform 1 0 23644 0 -1 19010
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_252
timestamp 1586364061
transform 1 0 24288 0 -1 19010
box -38 -48 774 592
use scs8hd_buf_2  _18_
timestamp 1586364061
transform 1 0 25024 0 -1 19010
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_264
timestamp 1586364061
transform 1 0 25392 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19010
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_288
timestamp 1586364061
transform 1 0 27600 0 -1 19010
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_296
timestamp 1586364061
transform 1 0 28336 0 -1 19010
box -38 -48 314 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 28888 0 -1 19010
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19010
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19010
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 1 19010
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19010
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_68
timestamp 1586364061
transform 1 0 7360 0 1 19010
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 1 19010
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_129
timestamp 1586364061
transform 1 0 12972 0 1 19010
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 15180 0 1 19010
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_141
timestamp 1586364061
transform 1 0 14076 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_154
timestamp 1586364061
transform 1 0 15272 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_178
timestamp 1586364061
transform 1 0 17480 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_190
timestamp 1586364061
transform 1 0 18584 0 1 19010
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 20792 0 1 19010
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_202
timestamp 1586364061
transform 1 0 19688 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_215
timestamp 1586364061
transform 1 0 20884 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_227
timestamp 1586364061
transform 1 0 21988 0 1 19010
box -38 -48 1142 592
use scs8hd_buf_2  _17_
timestamp 1586364061
transform 1 0 23920 0 1 19010
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__17__A
timestamp 1586364061
transform 1 0 24472 0 1 19010
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_239
timestamp 1586364061
transform 1 0 23092 0 1 19010
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_247
timestamp 1586364061
transform 1 0 23828 0 1 19010
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_252
timestamp 1586364061
transform 1 0 24288 0 1 19010
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_256
timestamp 1586364061
transform 1 0 24656 0 1 19010
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 26404 0 1 19010
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_268
timestamp 1586364061
transform 1 0 25760 0 1 19010
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_274
timestamp 1586364061
transform 1 0 26312 0 1 19010
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19010
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_288
timestamp 1586364061
transform 1 0 27600 0 1 19010
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_296
timestamp 1586364061
transform 1 0 28336 0 1 19010
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 28888 0 1 19010
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20098
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_39
timestamp 1586364061
transform 1 0 4692 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_51
timestamp 1586364061
transform 1 0 5796 0 -1 20098
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20098
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 6716 0 -1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_62
timestamp 1586364061
transform 1 0 6808 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_86
timestamp 1586364061
transform 1 0 9016 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_98
timestamp 1586364061
transform 1 0 10120 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_110
timestamp 1586364061
transform 1 0 11224 0 -1 20098
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 12328 0 -1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_135
timestamp 1586364061
transform 1 0 13524 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_147
timestamp 1586364061
transform 1 0 14628 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_159
timestamp 1586364061
transform 1 0 15732 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20098
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 17940 0 -1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_184
timestamp 1586364061
transform 1 0 18032 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_196
timestamp 1586364061
transform 1 0 19136 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_208
timestamp 1586364061
transform 1 0 20240 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_220
timestamp 1586364061
transform 1 0 21344 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_232
timestamp 1586364061
transform 1 0 22448 0 -1 20098
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 23552 0 -1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_245
timestamp 1586364061
transform 1 0 23644 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_257
timestamp 1586364061
transform 1 0 24748 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_269
timestamp 1586364061
transform 1 0 25852 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_281
timestamp 1586364061
transform 1 0 26956 0 -1 20098
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_293
timestamp 1586364061
transform 1 0 28060 0 -1 20098
box -38 -48 590 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 28888 0 -1 20098
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20098
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21186
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 3956 0 1 20098
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20098
box -38 -48 406 592
use scs8hd_decap_12  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_39
timestamp 1586364061
transform 1 0 4692 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_44
timestamp 1586364061
transform 1 0 5152 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_51
timestamp 1586364061
transform 1 0 5796 0 -1 21186
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_59
timestamp 1586364061
transform 1 0 6532 0 -1 21186
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 -1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_62
timestamp 1586364061
transform 1 0 6808 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_74
timestamp 1586364061
transform 1 0 7912 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 9568 0 1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_80
timestamp 1586364061
transform 1 0 8464 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_93
timestamp 1586364061
transform 1 0 9660 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_86
timestamp 1586364061
transform 1 0 9016 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_98
timestamp 1586364061
transform 1 0 10120 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_110
timestamp 1586364061
transform 1 0 11224 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 -1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_129
timestamp 1586364061
transform 1 0 12972 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_135
timestamp 1586364061
transform 1 0 13524 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 15180 0 1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_141
timestamp 1586364061
transform 1 0 14076 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_147
timestamp 1586364061
transform 1 0 14628 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_166
timestamp 1586364061
transform 1 0 16376 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_178
timestamp 1586364061
transform 1 0 17480 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_159
timestamp 1586364061
transform 1 0 15732 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_171
timestamp 1586364061
transform 1 0 16836 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 17940 0 -1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_190
timestamp 1586364061
transform 1 0 18584 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_184
timestamp 1586364061
transform 1 0 18032 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_196
timestamp 1586364061
transform 1 0 19136 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 20792 0 1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_215
timestamp 1586364061
transform 1 0 20884 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_208
timestamp 1586364061
transform 1 0 20240 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_227
timestamp 1586364061
transform 1 0 21988 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_220
timestamp 1586364061
transform 1 0 21344 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_232
timestamp 1586364061
transform 1 0 22448 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 23552 0 -1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_239
timestamp 1586364061
transform 1 0 23092 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_251
timestamp 1586364061
transform 1 0 24196 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_245
timestamp 1586364061
transform 1 0 23644 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_257
timestamp 1586364061
transform 1 0 24748 0 -1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 26404 0 1 20098
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_263
timestamp 1586364061
transform 1 0 25300 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_276
timestamp 1586364061
transform 1 0 26496 0 1 20098
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_269
timestamp 1586364061
transform 1 0 25852 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_288
timestamp 1586364061
transform 1 0 27600 0 1 20098
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_296
timestamp 1586364061
transform 1 0 28336 0 1 20098
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_281
timestamp 1586364061
transform 1 0 26956 0 -1 21186
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_293
timestamp 1586364061
transform 1 0 28060 0 -1 21186
box -38 -48 590 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 28888 0 1 20098
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 28888 0 -1 21186
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21186
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 3956 0 1 21186
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21186
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21186
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 6808 0 1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 9660 0 1 21186
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21186
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21186
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 12512 0 1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 15364 0 1 21186
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21186
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 18216 0 1 21186
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21186
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 21068 0 1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21186
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21186
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23920 0 1 21186
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_242
timestamp 1586364061
transform 1 0 23368 0 1 21186
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_249
timestamp 1586364061
transform 1 0 24012 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_261
timestamp 1586364061
transform 1 0 25116 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_273
timestamp 1586364061
transform 1 0 26220 0 1 21186
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26772 0 1 21186
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_280
timestamp 1586364061
transform 1 0 26864 0 1 21186
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_292
timestamp 1586364061
transform 1 0 27968 0 1 21186
box -38 -48 590 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 28888 0 1 21186
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_298
timestamp 1586364061
transform 1 0 28520 0 1 21186
box -38 -48 130 592
<< labels >>
rlabel metal2 s 11150 23490 11206 23970 6 ccff_head
port 0 nsew default input
rlabel metal2 s 18694 23490 18750 23970 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 12218 480 12338 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 18202 480 18322 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 18746 480 18866 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 19290 480 19410 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 19970 480 20090 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 20514 480 20634 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 21194 480 21314 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 21738 480 21858 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 22282 480 22402 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 22962 480 23082 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 23506 480 23626 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 12762 480 12882 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 13306 480 13426 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 13986 480 14106 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 14530 480 14650 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 15210 480 15330 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 15754 480 15874 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 16298 480 16418 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 16978 480 17098 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 17522 480 17642 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 250 480 370 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 6234 480 6354 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 6778 480 6898 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 7322 480 7442 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 8002 480 8122 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 8546 480 8666 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 9226 480 9346 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 9770 480 9890 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 10314 480 10434 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 10994 480 11114 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 11538 480 11658 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 794 480 914 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 1338 480 1458 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 2018 480 2138 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 2562 480 2682 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 3242 480 3362 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 3786 480 3906 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 4330 480 4450 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 5010 480 5130 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 5554 480 5674 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 29520 12218 30000 12338 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 29520 18202 30000 18322 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 29520 18746 30000 18866 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 29520 19290 30000 19410 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 29520 19970 30000 20090 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 29520 20514 30000 20634 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 29520 21194 30000 21314 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 29520 21738 30000 21858 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 29520 22282 30000 22402 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 29520 22962 30000 23082 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 29520 23506 30000 23626 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 29520 12762 30000 12882 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 29520 13306 30000 13426 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 29520 13986 30000 14106 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 29520 14530 30000 14650 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 29520 15210 30000 15330 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 29520 15754 30000 15874 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 29520 16298 30000 16418 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 29520 16978 30000 17098 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 29520 17522 30000 17642 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 29520 250 30000 370 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 29520 6234 30000 6354 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 29520 6778 30000 6898 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 29520 7322 30000 7442 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 29520 8002 30000 8122 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 29520 8546 30000 8666 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 29520 9226 30000 9346 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 29520 9770 30000 9890 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 29520 10314 30000 10434 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 29520 10994 30000 11114 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 29520 11538 30000 11658 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 29520 794 30000 914 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 29520 1338 30000 1458 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 29520 2018 30000 2138 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 29520 2562 30000 2682 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 29520 3242 30000 3362 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 29520 3786 30000 3906 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 29520 4330 30000 4450 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 29520 5010 30000 5130 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 29520 5554 30000 5674 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 3698 23490 3754 23970 6 prog_clk
port 82 nsew default input
rlabel metal2 s 26146 23490 26202 23970 6 top_grid_pin_0_
port 83 nsew default tristate
rlabel metal4 s 5944 2098 6264 21778 6 vpwr
port 84 nsew default input
rlabel metal4 s 10944 2098 11264 21778 6 vgnd
port 85 nsew default input
<< properties >>
string FIXED_BBOX 0 1 30000 23970
<< end >>
