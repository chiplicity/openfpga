magic
tech sky130A
magscale 1 2
timestamp 1606928802
<< locali >>
rect 9413 13243 9447 13345
rect 8493 12087 8527 12393
rect 9413 12155 9447 12257
rect 3525 11679 3559 11849
rect 3617 11543 3651 11713
rect 6561 10455 6595 10693
rect 6653 9435 6687 9673
rect 7757 9367 7791 9605
rect 11897 8959 11931 9061
rect 15117 9027 15151 9129
rect 15117 8823 15151 8993
rect 4353 8483 4387 8585
rect 3801 7735 3835 8041
rect 4905 7735 4939 7973
rect 16221 7735 16255 7837
rect 3893 6783 3927 6885
rect 3341 6171 3375 6341
rect 3709 6103 3743 6273
rect 8677 5083 8711 5321
rect 12265 4607 12299 4709
rect 5181 3519 5215 3689
rect 6837 3519 6871 3689
rect 10517 3383 10551 3553
rect 12081 3451 12115 3689
rect 12265 2839 12299 3145
rect 6929 2499 6963 2601
<< viali >>
rect 15945 14501 15979 14535
rect 16865 14501 16899 14535
rect 2145 14433 2179 14467
rect 3341 14433 3375 14467
rect 5089 14433 5123 14467
rect 17509 14433 17543 14467
rect 17601 14433 17635 14467
rect 2237 14365 2271 14399
rect 2421 14365 2455 14399
rect 3433 14365 3467 14399
rect 3525 14365 3559 14399
rect 5181 14365 5215 14399
rect 5273 14365 5307 14399
rect 15853 14365 15887 14399
rect 17693 14365 17727 14399
rect 1777 14229 1811 14263
rect 2973 14229 3007 14263
rect 4721 14229 4755 14263
rect 17141 14229 17175 14263
rect 2053 14025 2087 14059
rect 4721 14025 4755 14059
rect 6837 14025 6871 14059
rect 8125 14025 8159 14059
rect 17509 14025 17543 14059
rect 3709 13957 3743 13991
rect 5733 13957 5767 13991
rect 10149 13957 10183 13991
rect 14197 13957 14231 13991
rect 18245 13957 18279 13991
rect 2605 13889 2639 13923
rect 4261 13889 4295 13923
rect 5365 13889 5399 13923
rect 6377 13889 6411 13923
rect 7481 13889 7515 13923
rect 8585 13889 8619 13923
rect 8769 13889 8803 13923
rect 9689 13889 9723 13923
rect 10793 13889 10827 13923
rect 13737 13889 13771 13923
rect 14749 13889 14783 13923
rect 16037 13889 16071 13923
rect 17049 13889 17083 13923
rect 4169 13821 4203 13855
rect 5181 13821 5215 13855
rect 7297 13821 7331 13855
rect 10609 13821 10643 13855
rect 12817 13821 12851 13855
rect 13001 13821 13035 13855
rect 13369 13821 13403 13855
rect 14657 13821 14691 13855
rect 15520 13821 15554 13855
rect 17325 13821 17359 13855
rect 18061 13821 18095 13855
rect 2513 13753 2547 13787
rect 4077 13753 4111 13787
rect 9505 13753 9539 13787
rect 16129 13753 16163 13787
rect 2421 13685 2455 13719
rect 5089 13685 5123 13719
rect 6101 13685 6135 13719
rect 6193 13685 6227 13719
rect 7205 13685 7239 13719
rect 8493 13685 8527 13719
rect 9137 13685 9171 13719
rect 9597 13685 9631 13719
rect 10517 13685 10551 13719
rect 14565 13685 14599 13719
rect 15623 13685 15657 13719
rect 1961 13481 1995 13515
rect 2329 13481 2363 13515
rect 2973 13481 3007 13515
rect 4813 13481 4847 13515
rect 5825 13481 5859 13515
rect 8217 13481 8251 13515
rect 8953 13481 8987 13515
rect 14197 13481 14231 13515
rect 14565 13481 14599 13515
rect 15301 13481 15335 13515
rect 16313 13481 16347 13515
rect 17325 13481 17359 13515
rect 7104 13413 7138 13447
rect 10333 13413 10367 13447
rect 12265 13413 12299 13447
rect 17785 13413 17819 13447
rect 2421 13345 2455 13379
rect 3341 13345 3375 13379
rect 5181 13345 5215 13379
rect 6193 13345 6227 13379
rect 9413 13345 9447 13379
rect 11345 13345 11379 13379
rect 11437 13345 11471 13379
rect 11989 13345 12023 13379
rect 13553 13345 13587 13379
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 16681 13345 16715 13379
rect 17693 13345 17727 13379
rect 2513 13277 2547 13311
rect 3433 13277 3467 13311
rect 3525 13277 3559 13311
rect 5273 13277 5307 13311
rect 5457 13277 5491 13311
rect 6285 13277 6319 13311
rect 6469 13277 6503 13311
rect 6837 13277 6871 13311
rect 9045 13277 9079 13311
rect 9137 13277 9171 13311
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 11529 13277 11563 13311
rect 13645 13277 13679 13311
rect 13737 13277 13771 13311
rect 14657 13277 14691 13311
rect 14841 13277 14875 13311
rect 15945 13277 15979 13311
rect 16773 13277 16807 13311
rect 16865 13277 16899 13311
rect 17877 13277 17911 13311
rect 9413 13209 9447 13243
rect 8585 13141 8619 13175
rect 9965 13141 9999 13175
rect 10977 13141 11011 13175
rect 13185 13141 13219 13175
rect 1869 12937 1903 12971
rect 4261 12937 4295 12971
rect 11161 12937 11195 12971
rect 16313 12937 16347 12971
rect 16589 12937 16623 12971
rect 8217 12869 8251 12903
rect 13829 12869 13863 12903
rect 2421 12801 2455 12835
rect 5273 12801 5307 12835
rect 6377 12801 6411 12835
rect 10793 12801 10827 12835
rect 11713 12801 11747 12835
rect 14473 12801 14507 12835
rect 17233 12801 17267 12835
rect 2237 12733 2271 12767
rect 2881 12733 2915 12767
rect 5181 12733 5215 12767
rect 6837 12733 6871 12767
rect 8493 12733 8527 12767
rect 8760 12733 8794 12767
rect 10517 12733 10551 12767
rect 12449 12733 12483 12767
rect 12716 12733 12750 12767
rect 14933 12733 14967 12767
rect 15200 12733 15234 12767
rect 3148 12665 3182 12699
rect 5089 12665 5123 12699
rect 6101 12665 6135 12699
rect 7104 12665 7138 12699
rect 10609 12665 10643 12699
rect 11621 12665 11655 12699
rect 16957 12665 16991 12699
rect 2329 12597 2363 12631
rect 4721 12597 4755 12631
rect 5733 12597 5767 12631
rect 6193 12597 6227 12631
rect 9873 12597 9907 12631
rect 10149 12597 10183 12631
rect 11529 12597 11563 12631
rect 17049 12597 17083 12631
rect 1961 12393 1995 12427
rect 2973 12393 3007 12427
rect 3433 12393 3467 12427
rect 5457 12393 5491 12427
rect 5733 12393 5767 12427
rect 8033 12393 8067 12427
rect 8493 12393 8527 12427
rect 8585 12393 8619 12427
rect 9689 12393 9723 12427
rect 11621 12393 11655 12427
rect 14657 12393 14691 12427
rect 15301 12393 15335 12427
rect 4344 12325 4378 12359
rect 7941 12325 7975 12359
rect 2329 12257 2363 12291
rect 2421 12257 2455 12291
rect 3341 12257 3375 12291
rect 6929 12257 6963 12291
rect 2605 12189 2639 12223
rect 3617 12189 3651 12223
rect 4077 12189 4111 12223
rect 7021 12189 7055 12223
rect 7205 12189 7239 12223
rect 8125 12189 8159 12223
rect 10508 12325 10542 12359
rect 13544 12325 13578 12359
rect 8953 12257 8987 12291
rect 9413 12257 9447 12291
rect 12633 12257 12667 12291
rect 15669 12257 15703 12291
rect 16672 12257 16706 12291
rect 9045 12189 9079 12223
rect 9229 12189 9263 12223
rect 10241 12189 10275 12223
rect 12725 12189 12759 12223
rect 12909 12189 12943 12223
rect 13277 12189 13311 12223
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 16405 12189 16439 12223
rect 9413 12121 9447 12155
rect 6561 12053 6595 12087
rect 7573 12053 7607 12087
rect 8493 12053 8527 12087
rect 12265 12053 12299 12087
rect 17785 12053 17819 12087
rect 2697 11849 2731 11883
rect 3525 11849 3559 11883
rect 9321 11849 9355 11883
rect 13093 11849 13127 11883
rect 14105 11849 14139 11883
rect 1685 11781 1719 11815
rect 2329 11713 2363 11747
rect 3341 11713 3375 11747
rect 2053 11645 2087 11679
rect 3525 11645 3559 11679
rect 3617 11713 3651 11747
rect 6377 11713 6411 11747
rect 9873 11713 9907 11747
rect 10977 11713 11011 11747
rect 11989 11713 12023 11747
rect 13553 11713 13587 11747
rect 13737 11713 13771 11747
rect 14657 11713 14691 11747
rect 3065 11577 3099 11611
rect 3709 11645 3743 11679
rect 3965 11645 3999 11679
rect 6101 11645 6135 11679
rect 7481 11645 7515 11679
rect 7573 11645 7607 11679
rect 7840 11645 7874 11679
rect 9689 11645 9723 11679
rect 11713 11645 11747 11679
rect 14473 11645 14507 11679
rect 14565 11645 14599 11679
rect 15393 11645 15427 11679
rect 6193 11577 6227 11611
rect 10793 11577 10827 11611
rect 15638 11577 15672 11611
rect 2145 11509 2179 11543
rect 3157 11509 3191 11543
rect 3617 11509 3651 11543
rect 5089 11509 5123 11543
rect 5733 11509 5767 11543
rect 7297 11509 7331 11543
rect 8953 11509 8987 11543
rect 9781 11509 9815 11543
rect 10333 11509 10367 11543
rect 10701 11509 10735 11543
rect 11345 11509 11379 11543
rect 11805 11509 11839 11543
rect 13461 11509 13495 11543
rect 16773 11509 16807 11543
rect 1685 11305 1719 11339
rect 8585 11305 8619 11339
rect 10517 11305 10551 11339
rect 14197 11305 14231 11339
rect 14473 11305 14507 11339
rect 16681 11305 16715 11339
rect 16957 11305 16991 11339
rect 7941 11237 7975 11271
rect 8953 11237 8987 11271
rect 11428 11237 11462 11271
rect 17325 11237 17359 11271
rect 1501 11169 1535 11203
rect 2053 11169 2087 11203
rect 2320 11169 2354 11203
rect 4344 11169 4378 11203
rect 6745 11169 6779 11203
rect 8033 11169 8067 11203
rect 9045 11169 9079 11203
rect 10609 11169 10643 11203
rect 13084 11169 13118 11203
rect 15568 11169 15602 11203
rect 17417 11169 17451 11203
rect 4077 11101 4111 11135
rect 6837 11101 6871 11135
rect 7021 11101 7055 11135
rect 8217 11101 8251 11135
rect 9229 11101 9263 11135
rect 10793 11101 10827 11135
rect 11161 11101 11195 11135
rect 12817 11101 12851 11135
rect 15301 11101 15335 11135
rect 17601 11101 17635 11135
rect 3433 11033 3467 11067
rect 5457 11033 5491 11067
rect 6377 11033 6411 11067
rect 7573 11033 7607 11067
rect 10149 11033 10183 11067
rect 12541 11033 12575 11067
rect 3709 10761 3743 10795
rect 4721 10761 4755 10795
rect 8217 10761 8251 10795
rect 9873 10761 9907 10795
rect 17509 10761 17543 10795
rect 6561 10693 6595 10727
rect 11805 10693 11839 10727
rect 1409 10625 1443 10659
rect 2329 10625 2363 10659
rect 2513 10625 2547 10659
rect 4353 10625 4387 10659
rect 5273 10625 5307 10659
rect 6285 10625 6319 10659
rect 2237 10557 2271 10591
rect 2881 10557 2915 10591
rect 3617 10557 3651 10591
rect 4077 10557 4111 10591
rect 5181 10557 5215 10591
rect 4169 10489 4203 10523
rect 6837 10625 6871 10659
rect 15761 10625 15795 10659
rect 8493 10557 8527 10591
rect 8749 10557 8783 10591
rect 10149 10557 10183 10591
rect 11989 10557 12023 10591
rect 12909 10557 12943 10591
rect 13277 10557 13311 10591
rect 16129 10557 16163 10591
rect 7082 10489 7116 10523
rect 10394 10489 10428 10523
rect 13522 10489 13556 10523
rect 16396 10489 16430 10523
rect 1869 10421 1903 10455
rect 3065 10421 3099 10455
rect 3433 10421 3467 10455
rect 5089 10421 5123 10455
rect 5733 10421 5767 10455
rect 6101 10421 6135 10455
rect 6193 10421 6227 10455
rect 6561 10421 6595 10455
rect 11529 10421 11563 10455
rect 12725 10421 12759 10455
rect 14657 10421 14691 10455
rect 15117 10421 15151 10455
rect 15485 10421 15519 10455
rect 15577 10421 15611 10455
rect 2789 10217 2823 10251
rect 7113 10217 7147 10251
rect 7573 10217 7607 10251
rect 9045 10217 9079 10251
rect 11069 10217 11103 10251
rect 11989 10217 12023 10251
rect 13001 10217 13035 10251
rect 14381 10217 14415 10251
rect 17141 10217 17175 10251
rect 1676 10149 1710 10183
rect 4813 10149 4847 10183
rect 7941 10149 7975 10183
rect 12357 10149 12391 10183
rect 13461 10149 13495 10183
rect 17509 10149 17543 10183
rect 3065 10081 3099 10115
rect 5457 10081 5491 10115
rect 5724 10081 5758 10115
rect 7297 10081 7331 10115
rect 8033 10081 8067 10115
rect 8953 10081 8987 10115
rect 9689 10081 9723 10115
rect 9956 10081 9990 10115
rect 13369 10081 13403 10115
rect 15669 10081 15703 10115
rect 16497 10081 16531 10115
rect 16589 10081 16623 10115
rect 1409 10013 1443 10047
rect 4905 10013 4939 10047
rect 5089 10013 5123 10047
rect 8125 10013 8159 10047
rect 9137 10013 9171 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 13553 10013 13587 10047
rect 14473 10013 14507 10047
rect 14565 10013 14599 10047
rect 16773 10013 16807 10047
rect 17601 10013 17635 10047
rect 17785 10013 17819 10047
rect 18153 10013 18187 10047
rect 6837 9945 6871 9979
rect 14013 9945 14047 9979
rect 3249 9877 3283 9911
rect 4445 9877 4479 9911
rect 8585 9877 8619 9911
rect 15485 9877 15519 9911
rect 16129 9877 16163 9911
rect 4721 9673 4755 9707
rect 6653 9673 6687 9707
rect 6837 9673 6871 9707
rect 11345 9673 11379 9707
rect 5733 9605 5767 9639
rect 2329 9537 2363 9571
rect 5365 9537 5399 9571
rect 6377 9537 6411 9571
rect 1685 9469 1719 9503
rect 3985 9469 4019 9503
rect 5089 9469 5123 9503
rect 7757 9605 7791 9639
rect 7849 9605 7883 9639
rect 9505 9605 9539 9639
rect 10333 9605 10367 9639
rect 13829 9605 13863 9639
rect 7389 9537 7423 9571
rect 2574 9401 2608 9435
rect 6101 9401 6135 9435
rect 6653 9401 6687 9435
rect 7205 9401 7239 9435
rect 8401 9537 8435 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 10977 9537 11011 9571
rect 11989 9537 12023 9571
rect 12449 9537 12483 9571
rect 16313 9537 16347 9571
rect 8309 9469 8343 9503
rect 10793 9469 10827 9503
rect 14105 9469 14139 9503
rect 14372 9469 14406 9503
rect 8217 9401 8251 9435
rect 8861 9401 8895 9435
rect 12716 9401 12750 9435
rect 16580 9401 16614 9435
rect 1869 9333 1903 9367
rect 3709 9333 3743 9367
rect 4169 9333 4203 9367
rect 5181 9333 5215 9367
rect 6193 9333 6227 9367
rect 7297 9333 7331 9367
rect 7757 9333 7791 9367
rect 9873 9333 9907 9367
rect 10701 9333 10735 9367
rect 11713 9333 11747 9367
rect 11805 9333 11839 9367
rect 15485 9333 15519 9367
rect 17693 9333 17727 9367
rect 1961 9129 1995 9163
rect 2329 9129 2363 9163
rect 7113 9129 7147 9163
rect 8769 9129 8803 9163
rect 10149 9129 10183 9163
rect 12081 9129 12115 9163
rect 12449 9129 12483 9163
rect 13093 9129 13127 9163
rect 13461 9129 13495 9163
rect 13553 9129 13587 9163
rect 15117 9129 15151 9163
rect 2421 9061 2455 9095
rect 4322 9061 4356 9095
rect 6000 9061 6034 9095
rect 7634 9061 7668 9095
rect 10609 9061 10643 9095
rect 11897 9061 11931 9095
rect 1409 8993 1443 9027
rect 3341 8993 3375 9027
rect 5733 8993 5767 9027
rect 10517 8993 10551 9027
rect 11437 8993 11471 9027
rect 15393 9061 15427 9095
rect 12541 8993 12575 9027
rect 14565 8993 14599 9027
rect 15117 8993 15151 9027
rect 16293 8993 16327 9027
rect 17877 8993 17911 9027
rect 2605 8925 2639 8959
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 4077 8925 4111 8959
rect 7389 8925 7423 8959
rect 10793 8925 10827 8959
rect 11529 8925 11563 8959
rect 11713 8925 11747 8959
rect 11897 8925 11931 8959
rect 12725 8925 12759 8959
rect 13645 8925 13679 8959
rect 14657 8925 14691 8959
rect 14749 8925 14783 8959
rect 1593 8857 1627 8891
rect 16037 8925 16071 8959
rect 2973 8789 3007 8823
rect 5457 8789 5491 8823
rect 11069 8789 11103 8823
rect 14197 8789 14231 8823
rect 15117 8789 15151 8823
rect 17417 8789 17451 8823
rect 18061 8789 18095 8823
rect 3525 8585 3559 8619
rect 4353 8585 4387 8619
rect 6837 8585 6871 8619
rect 8493 8585 8527 8619
rect 11069 8585 11103 8619
rect 11345 8585 11379 8619
rect 14105 8585 14139 8619
rect 6377 8517 6411 8551
rect 7849 8517 7883 8551
rect 12449 8517 12483 8551
rect 16773 8517 16807 8551
rect 18245 8517 18279 8551
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 4997 8449 5031 8483
rect 7481 8449 7515 8483
rect 11897 8449 11931 8483
rect 13001 8449 13035 8483
rect 14565 8449 14599 8483
rect 14657 8449 14691 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 1409 8381 1443 8415
rect 1676 8381 1710 8415
rect 7665 8381 7699 8415
rect 8677 8381 8711 8415
rect 10517 8381 10551 8415
rect 11253 8381 11287 8415
rect 15117 8381 15151 8415
rect 15384 8381 15418 8415
rect 18061 8381 18095 8415
rect 3893 8313 3927 8347
rect 5264 8313 5298 8347
rect 7205 8313 7239 8347
rect 7297 8313 7331 8347
rect 8033 8313 8067 8347
rect 8953 8313 8987 8347
rect 11713 8313 11747 8347
rect 11805 8313 11839 8347
rect 12909 8313 12943 8347
rect 2789 8245 2823 8279
rect 4537 8245 4571 8279
rect 12817 8245 12851 8279
rect 14473 8245 14507 8279
rect 16497 8245 16531 8279
rect 17141 8245 17175 8279
rect 2329 8041 2363 8075
rect 2973 8041 3007 8075
rect 3341 8041 3375 8075
rect 3801 8041 3835 8075
rect 4077 8041 4111 8075
rect 5549 8041 5583 8075
rect 6561 8041 6595 8075
rect 7297 8041 7331 8075
rect 7757 8041 7791 8075
rect 10885 8041 10919 8075
rect 12725 8041 12759 8075
rect 13001 8041 13035 8075
rect 14841 8041 14875 8075
rect 17325 8041 17359 8075
rect 17693 8041 17727 8075
rect 2421 7973 2455 8007
rect 3433 7973 3467 8007
rect 1409 7905 1443 7939
rect 2605 7837 2639 7871
rect 3617 7837 3651 7871
rect 1593 7769 1627 7803
rect 4905 7973 4939 8007
rect 7665 7973 7699 8007
rect 11612 7973 11646 8007
rect 13728 7973 13762 8007
rect 15669 7973 15703 8007
rect 16681 7973 16715 8007
rect 16773 7973 16807 8007
rect 4445 7905 4479 7939
rect 4537 7905 4571 7939
rect 4629 7837 4663 7871
rect 1961 7701 1995 7735
rect 3801 7701 3835 7735
rect 5457 7905 5491 7939
rect 8125 7905 8159 7939
rect 8392 7905 8426 7939
rect 10057 7905 10091 7939
rect 13461 7905 13495 7939
rect 5641 7837 5675 7871
rect 6653 7837 6687 7871
rect 6837 7837 6871 7871
rect 7849 7837 7883 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 11345 7837 11379 7871
rect 15761 7837 15795 7871
rect 15853 7837 15887 7871
rect 16221 7837 16255 7871
rect 16865 7837 16899 7871
rect 17785 7837 17819 7871
rect 17877 7837 17911 7871
rect 9689 7769 9723 7803
rect 15301 7769 15335 7803
rect 4905 7701 4939 7735
rect 5089 7701 5123 7735
rect 6193 7701 6227 7735
rect 9505 7701 9539 7735
rect 16221 7701 16255 7735
rect 16313 7701 16347 7735
rect 3801 7497 3835 7531
rect 6285 7497 6319 7531
rect 7205 7497 7239 7531
rect 11897 7497 11931 7531
rect 12449 7497 12483 7531
rect 13461 7497 13495 7531
rect 16497 7497 16531 7531
rect 18245 7497 18279 7531
rect 1685 7361 1719 7395
rect 3341 7361 3375 7395
rect 4445 7361 4479 7395
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 10517 7361 10551 7395
rect 12909 7361 12943 7395
rect 13093 7361 13127 7395
rect 14013 7361 14047 7395
rect 15117 7361 15151 7395
rect 16129 7361 16163 7395
rect 17049 7361 17083 7395
rect 1952 7293 1986 7327
rect 4169 7293 4203 7327
rect 4905 7293 4939 7327
rect 8677 7293 8711 7327
rect 8933 7293 8967 7327
rect 10784 7293 10818 7327
rect 13829 7293 13863 7327
rect 13921 7293 13955 7327
rect 14841 7293 14875 7327
rect 15853 7293 15887 7327
rect 15945 7293 15979 7327
rect 16865 7293 16899 7327
rect 18061 7293 18095 7327
rect 5172 7225 5206 7259
rect 16957 7225 16991 7259
rect 3065 7157 3099 7191
rect 4261 7157 4295 7191
rect 7573 7157 7607 7191
rect 10057 7157 10091 7191
rect 12817 7157 12851 7191
rect 14473 7157 14507 7191
rect 14933 7157 14967 7191
rect 15485 7157 15519 7191
rect 6377 6953 6411 6987
rect 8769 6953 8803 6987
rect 9873 6953 9907 6987
rect 11713 6953 11747 6987
rect 12725 6953 12759 6987
rect 13737 6953 13771 6987
rect 15669 6953 15703 6987
rect 16773 6953 16807 6987
rect 17877 6953 17911 6987
rect 3893 6885 3927 6919
rect 16681 6885 16715 6919
rect 1685 6817 1719 6851
rect 2596 6817 2630 6851
rect 4344 6817 4378 6851
rect 5733 6817 5767 6851
rect 6745 6817 6779 6851
rect 7656 6817 7690 6851
rect 10057 6817 10091 6851
rect 10333 6817 10367 6851
rect 10600 6817 10634 6851
rect 12173 6817 12207 6851
rect 17969 6817 18003 6851
rect 2329 6749 2363 6783
rect 3893 6749 3927 6783
rect 4077 6749 4111 6783
rect 6837 6749 6871 6783
rect 7021 6749 7055 6783
rect 7389 6749 7423 6783
rect 12817 6749 12851 6783
rect 13001 6749 13035 6783
rect 13829 6749 13863 6783
rect 14013 6749 14047 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 16865 6749 16899 6783
rect 18061 6749 18095 6783
rect 3709 6681 3743 6715
rect 15301 6681 15335 6715
rect 16313 6681 16347 6715
rect 17509 6681 17543 6715
rect 1869 6613 1903 6647
rect 5457 6613 5491 6647
rect 5917 6613 5951 6647
rect 11989 6613 12023 6647
rect 12357 6613 12391 6647
rect 13369 6613 13403 6647
rect 3433 6409 3467 6443
rect 8217 6409 8251 6443
rect 11345 6409 11379 6443
rect 13093 6409 13127 6443
rect 15485 6409 15519 6443
rect 17601 6409 17635 6443
rect 18245 6409 18279 6443
rect 3341 6341 3375 6375
rect 3801 6341 3835 6375
rect 6009 6341 6043 6375
rect 2053 6273 2087 6307
rect 2881 6273 2915 6307
rect 3065 6273 3099 6307
rect 2789 6205 2823 6239
rect 3709 6273 3743 6307
rect 4445 6273 4479 6307
rect 5365 6273 5399 6307
rect 11805 6273 11839 6307
rect 11989 6273 12023 6307
rect 13737 6273 13771 6307
rect 16313 6273 16347 6307
rect 3617 6205 3651 6239
rect 1869 6137 1903 6171
rect 3341 6137 3375 6171
rect 5273 6205 5307 6239
rect 5825 6205 5859 6239
rect 6653 6205 6687 6239
rect 6837 6205 6871 6239
rect 9229 6205 9263 6239
rect 11713 6205 11747 6239
rect 14105 6205 14139 6239
rect 17417 6205 17451 6239
rect 18061 6205 18095 6239
rect 7104 6137 7138 6171
rect 9496 6137 9530 6171
rect 13461 6137 13495 6171
rect 14372 6137 14406 6171
rect 16129 6137 16163 6171
rect 1409 6069 1443 6103
rect 1777 6069 1811 6103
rect 2421 6069 2455 6103
rect 3709 6069 3743 6103
rect 4169 6069 4203 6103
rect 4261 6069 4295 6103
rect 4813 6069 4847 6103
rect 5181 6069 5215 6103
rect 6469 6069 6503 6103
rect 8769 6069 8803 6103
rect 10609 6069 10643 6103
rect 13553 6069 13587 6103
rect 15761 6069 15795 6103
rect 16221 6069 16255 6103
rect 4169 5865 4203 5899
rect 4629 5865 4663 5899
rect 5273 5865 5307 5899
rect 6929 5865 6963 5899
rect 9229 5865 9263 5899
rect 14013 5865 14047 5899
rect 18061 5865 18095 5899
rect 5816 5797 5850 5831
rect 1593 5729 1627 5763
rect 1860 5729 1894 5763
rect 3249 5729 3283 5763
rect 4537 5729 4571 5763
rect 5457 5729 5491 5763
rect 5549 5729 5583 5763
rect 7205 5729 7239 5763
rect 8116 5729 8150 5763
rect 10149 5729 10183 5763
rect 10416 5729 10450 5763
rect 12900 5729 12934 5763
rect 14749 5729 14783 5763
rect 15669 5729 15703 5763
rect 16773 5729 16807 5763
rect 17325 5729 17359 5763
rect 17877 5729 17911 5763
rect 4721 5661 4755 5695
rect 7849 5661 7883 5695
rect 12633 5661 12667 5695
rect 15761 5661 15795 5695
rect 15945 5661 15979 5695
rect 17509 5593 17543 5627
rect 2973 5525 3007 5559
rect 3433 5525 3467 5559
rect 7389 5525 7423 5559
rect 11529 5525 11563 5559
rect 15301 5525 15335 5559
rect 16957 5525 16991 5559
rect 6101 5321 6135 5355
rect 7849 5321 7883 5355
rect 8677 5321 8711 5355
rect 8861 5321 8895 5355
rect 9873 5321 9907 5355
rect 13829 5321 13863 5355
rect 16037 5321 16071 5355
rect 1409 5185 1443 5219
rect 4537 5185 4571 5219
rect 5457 5185 5491 5219
rect 7389 5185 7423 5219
rect 8309 5185 8343 5219
rect 8401 5185 8435 5219
rect 1676 5117 1710 5151
rect 3065 5117 3099 5151
rect 5917 5117 5951 5151
rect 7205 5117 7239 5151
rect 8217 5117 8251 5151
rect 9505 5185 9539 5219
rect 10425 5185 10459 5219
rect 11805 5185 11839 5219
rect 11989 5185 12023 5219
rect 16589 5185 16623 5219
rect 9229 5117 9263 5151
rect 10241 5117 10275 5151
rect 12449 5117 12483 5151
rect 14381 5117 14415 5151
rect 14648 5117 14682 5151
rect 17417 5117 17451 5151
rect 18061 5117 18095 5151
rect 3341 5049 3375 5083
rect 4261 5049 4295 5083
rect 7297 5049 7331 5083
rect 8677 5049 8711 5083
rect 9321 5049 9355 5083
rect 11713 5049 11747 5083
rect 12716 5049 12750 5083
rect 16405 5049 16439 5083
rect 2789 4981 2823 5015
rect 3893 4981 3927 5015
rect 4353 4981 4387 5015
rect 4905 4981 4939 5015
rect 5273 4981 5307 5015
rect 5365 4981 5399 5015
rect 6837 4981 6871 5015
rect 10333 4981 10367 5015
rect 10885 4981 10919 5015
rect 11345 4981 11379 5015
rect 15761 4981 15795 5015
rect 16497 4981 16531 5015
rect 17601 4981 17635 5015
rect 18245 4981 18279 5015
rect 6193 4777 6227 4811
rect 11713 4777 11747 4811
rect 13093 4777 13127 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15301 4777 15335 4811
rect 15669 4777 15703 4811
rect 15761 4777 15795 4811
rect 6101 4709 6135 4743
rect 7205 4709 7239 4743
rect 8116 4709 8150 4743
rect 11805 4709 11839 4743
rect 12265 4709 12299 4743
rect 13001 4709 13035 4743
rect 14105 4709 14139 4743
rect 1501 4641 1535 4675
rect 2320 4641 2354 4675
rect 4344 4641 4378 4675
rect 7113 4641 7147 4675
rect 9689 4641 9723 4675
rect 9956 4641 9990 4675
rect 12541 4641 12575 4675
rect 17877 4641 17911 4675
rect 2053 4573 2087 4607
rect 4077 4573 4111 4607
rect 6377 4573 6411 4607
rect 7297 4573 7331 4607
rect 7849 4573 7883 4607
rect 11897 4573 11931 4607
rect 12265 4573 12299 4607
rect 13277 4573 13311 4607
rect 14289 4573 14323 4607
rect 15945 4573 15979 4607
rect 9229 4505 9263 4539
rect 1685 4437 1719 4471
rect 3433 4437 3467 4471
rect 5457 4437 5491 4471
rect 5733 4437 5767 4471
rect 6745 4437 6779 4471
rect 11069 4437 11103 4471
rect 11345 4437 11379 4471
rect 12357 4437 12391 4471
rect 12633 4437 12667 4471
rect 18061 4437 18095 4471
rect 3985 4233 4019 4267
rect 15025 4233 15059 4267
rect 2605 4097 2639 4131
rect 5457 4097 5491 4131
rect 8309 4097 8343 4131
rect 9321 4097 9355 4131
rect 9965 4097 9999 4131
rect 13093 4097 13127 4131
rect 13277 4097 13311 4131
rect 1593 4029 1627 4063
rect 4261 4029 4295 4063
rect 5273 4029 5307 4063
rect 5917 4029 5951 4063
rect 6837 4029 6871 4063
rect 8217 4029 8251 4063
rect 9781 4029 9815 4063
rect 10701 4029 10735 4063
rect 13001 4029 13035 4063
rect 13645 4029 13679 4063
rect 17417 4029 17451 4063
rect 18061 4029 18095 4063
rect 1869 3961 1903 3995
rect 2872 3961 2906 3995
rect 6193 3961 6227 3995
rect 7113 3961 7147 3995
rect 9137 3961 9171 3995
rect 10946 3961 10980 3995
rect 13912 3961 13946 3995
rect 4445 3893 4479 3927
rect 4905 3893 4939 3927
rect 5365 3893 5399 3927
rect 7757 3893 7791 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 9229 3893 9263 3927
rect 12081 3893 12115 3927
rect 12633 3893 12667 3927
rect 17601 3893 17635 3927
rect 18245 3893 18279 3927
rect 1593 3689 1627 3723
rect 1961 3689 1995 3723
rect 3433 3689 3467 3723
rect 4629 3689 4663 3723
rect 5181 3689 5215 3723
rect 1409 3553 1443 3587
rect 2329 3553 2363 3587
rect 3341 3553 3375 3587
rect 6837 3689 6871 3723
rect 8585 3689 8619 3723
rect 9045 3689 9079 3723
rect 9689 3689 9723 3723
rect 10057 3689 10091 3723
rect 10701 3689 10735 3723
rect 12081 3689 12115 3723
rect 14289 3689 14323 3723
rect 5518 3621 5552 3655
rect 8953 3621 8987 3655
rect 10149 3621 10183 3655
rect 7185 3553 7219 3587
rect 10517 3553 10551 3587
rect 11069 3553 11103 3587
rect 2421 3485 2455 3519
rect 2605 3485 2639 3519
rect 3525 3485 3559 3519
rect 4721 3485 4755 3519
rect 4905 3485 4939 3519
rect 5181 3485 5215 3519
rect 5273 3485 5307 3519
rect 6837 3485 6871 3519
rect 6929 3485 6963 3519
rect 9229 3485 9263 3519
rect 10241 3485 10275 3519
rect 11161 3485 11195 3519
rect 11253 3485 11287 3519
rect 12440 3553 12474 3587
rect 14197 3553 14231 3587
rect 17233 3553 17267 3587
rect 17785 3553 17819 3587
rect 12173 3485 12207 3519
rect 14381 3485 14415 3519
rect 12081 3417 12115 3451
rect 13553 3417 13587 3451
rect 2973 3349 3007 3383
rect 4261 3349 4295 3383
rect 6653 3349 6687 3383
rect 8309 3349 8343 3383
rect 10517 3349 10551 3383
rect 13829 3349 13863 3383
rect 17417 3349 17451 3383
rect 17969 3349 18003 3383
rect 2697 3145 2731 3179
rect 4629 3145 4663 3179
rect 8493 3145 8527 3179
rect 12265 3145 12299 3179
rect 13461 3145 13495 3179
rect 16313 3145 16347 3179
rect 10517 3077 10551 3111
rect 3249 3009 3283 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 6101 3009 6135 3043
rect 6193 3009 6227 3043
rect 8033 3009 8067 3043
rect 9045 3009 9079 3043
rect 10057 3009 10091 3043
rect 11069 3009 11103 3043
rect 1593 2941 1627 2975
rect 3893 2941 3927 2975
rect 7205 2941 7239 2975
rect 8953 2941 8987 2975
rect 9873 2941 9907 2975
rect 10885 2941 10919 2975
rect 11621 2941 11655 2975
rect 1869 2873 1903 2907
rect 3157 2873 3191 2907
rect 4169 2873 4203 2907
rect 4997 2873 5031 2907
rect 11897 2873 11931 2907
rect 12449 3077 12483 3111
rect 13093 3009 13127 3043
rect 13921 3009 13955 3043
rect 14013 3009 14047 3043
rect 14473 2941 14507 2975
rect 15209 2941 15243 2975
rect 15485 2941 15519 2975
rect 16129 2941 16163 2975
rect 16865 2941 16899 2975
rect 17417 2941 17451 2975
rect 18061 2941 18095 2975
rect 12817 2873 12851 2907
rect 14749 2873 14783 2907
rect 3065 2805 3099 2839
rect 5641 2805 5675 2839
rect 6009 2805 6043 2839
rect 8861 2805 8895 2839
rect 9505 2805 9539 2839
rect 9965 2805 9999 2839
rect 10977 2805 11011 2839
rect 12265 2805 12299 2839
rect 12909 2805 12943 2839
rect 13829 2805 13863 2839
rect 17049 2805 17083 2839
rect 17601 2805 17635 2839
rect 18245 2805 18279 2839
rect 1685 2601 1719 2635
rect 2973 2601 3007 2635
rect 3433 2601 3467 2635
rect 4077 2601 4111 2635
rect 4997 2601 5031 2635
rect 6469 2601 6503 2635
rect 6929 2601 6963 2635
rect 9137 2601 9171 2635
rect 11345 2601 11379 2635
rect 11805 2601 11839 2635
rect 4905 2533 4939 2567
rect 11713 2533 11747 2567
rect 14933 2533 14967 2567
rect 1501 2465 1535 2499
rect 2053 2465 2087 2499
rect 3341 2465 3375 2499
rect 5549 2465 5583 2499
rect 6285 2465 6319 2499
rect 6929 2465 6963 2499
rect 7021 2465 7055 2499
rect 7757 2465 7791 2499
rect 9045 2465 9079 2499
rect 9781 2465 9815 2499
rect 10701 2465 10735 2499
rect 13185 2465 13219 2499
rect 13921 2465 13955 2499
rect 14657 2465 14691 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 2237 2397 2271 2431
rect 3617 2397 3651 2431
rect 5089 2397 5123 2431
rect 5733 2397 5767 2431
rect 7297 2397 7331 2431
rect 7941 2397 7975 2431
rect 9321 2397 9355 2431
rect 10793 2397 10827 2431
rect 10977 2397 11011 2431
rect 11897 2397 11931 2431
rect 13369 2397 13403 2431
rect 14105 2397 14139 2431
rect 9965 2329 9999 2363
rect 4537 2261 4571 2295
rect 8677 2261 8711 2295
rect 10333 2261 10367 2295
rect 17325 2261 17359 2295
rect 17877 2261 17911 2295
<< metal1 >>
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 5074 15416 5080 15428
rect 4120 15388 5080 15416
rect 4120 15376 4126 15388
rect 5074 15376 5080 15388
rect 5132 15376 5138 15428
rect 3694 15172 3700 15224
rect 3752 15212 3758 15224
rect 5902 15212 5908 15224
rect 3752 15184 5908 15212
rect 3752 15172 3758 15184
rect 5902 15172 5908 15184
rect 5960 15172 5966 15224
rect 3786 14832 3792 14884
rect 3844 14872 3850 14884
rect 10870 14872 10876 14884
rect 3844 14844 10876 14872
rect 3844 14832 3850 14844
rect 10870 14832 10876 14844
rect 10928 14832 10934 14884
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 17862 14804 17868 14816
rect 9456 14776 17868 14804
rect 9456 14764 9462 14776
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 2700 14504 3556 14532
rect 2038 14424 2044 14476
rect 2096 14464 2102 14476
rect 2133 14467 2191 14473
rect 2133 14464 2145 14467
rect 2096 14436 2145 14464
rect 2096 14424 2102 14436
rect 2133 14433 2145 14436
rect 2179 14433 2191 14467
rect 2133 14427 2191 14433
rect 2700 14408 2728 14504
rect 3050 14424 3056 14476
rect 3108 14464 3114 14476
rect 3329 14467 3387 14473
rect 3329 14464 3341 14467
rect 3108 14436 3341 14464
rect 3108 14424 3114 14436
rect 3329 14433 3341 14436
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 2222 14396 2228 14408
rect 2183 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2409 14399 2467 14405
rect 2409 14365 2421 14399
rect 2455 14396 2467 14399
rect 2682 14396 2688 14408
rect 2455 14368 2688 14396
rect 2455 14365 2467 14368
rect 2409 14359 2467 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3418 14396 3424 14408
rect 3379 14368 3424 14396
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 3528 14405 3556 14504
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 10318 14532 10324 14544
rect 3752 14504 10324 14532
rect 3752 14492 3758 14504
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 15933 14535 15991 14541
rect 15933 14532 15945 14535
rect 14424 14504 15945 14532
rect 14424 14492 14430 14504
rect 15933 14501 15945 14504
rect 15979 14501 15991 14535
rect 15933 14495 15991 14501
rect 16853 14535 16911 14541
rect 16853 14501 16865 14535
rect 16899 14532 16911 14535
rect 18782 14532 18788 14544
rect 16899 14504 18788 14532
rect 16899 14501 16911 14504
rect 16853 14495 16911 14501
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 4706 14424 4712 14476
rect 4764 14464 4770 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4764 14436 5089 14464
rect 4764 14424 4770 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 17494 14464 17500 14476
rect 17455 14436 17500 14464
rect 5077 14427 5135 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 17586 14424 17592 14476
rect 17644 14464 17650 14476
rect 17644 14436 17689 14464
rect 17644 14424 17650 14436
rect 3513 14399 3571 14405
rect 3513 14365 3525 14399
rect 3559 14365 3571 14399
rect 5166 14396 5172 14408
rect 5127 14368 5172 14396
rect 3513 14359 3571 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 5316 14368 5361 14396
rect 5316 14356 5322 14368
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 13354 14396 13360 14408
rect 10008 14368 13360 14396
rect 10008 14356 10014 14368
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 15102 14356 15108 14408
rect 15160 14396 15166 14408
rect 15562 14396 15568 14408
rect 15160 14368 15568 14396
rect 15160 14356 15166 14368
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 16114 14396 16120 14408
rect 15887 14368 16120 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17368 14368 17693 14396
rect 17368 14356 17374 14368
rect 17681 14365 17693 14368
rect 17727 14365 17739 14399
rect 17681 14359 17739 14365
rect 3326 14288 3332 14340
rect 3384 14328 3390 14340
rect 18046 14328 18052 14340
rect 3384 14300 18052 14328
rect 3384 14288 3390 14300
rect 18046 14288 18052 14300
rect 18104 14288 18110 14340
rect 1762 14260 1768 14272
rect 1723 14232 1768 14260
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 2866 14220 2872 14272
rect 2924 14260 2930 14272
rect 2961 14263 3019 14269
rect 2961 14260 2973 14263
rect 2924 14232 2973 14260
rect 2924 14220 2930 14232
rect 2961 14229 2973 14232
rect 3007 14229 3019 14263
rect 2961 14223 3019 14229
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4709 14263 4767 14269
rect 4709 14260 4721 14263
rect 4304 14232 4721 14260
rect 4304 14220 4310 14232
rect 4709 14229 4721 14232
rect 4755 14229 4767 14263
rect 4709 14223 4767 14229
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 10778 14260 10784 14272
rect 8168 14232 10784 14260
rect 8168 14220 8174 14232
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 15102 14260 15108 14272
rect 10928 14232 15108 14260
rect 10928 14220 10934 14232
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 15194 14220 15200 14272
rect 15252 14260 15258 14272
rect 17129 14263 17187 14269
rect 17129 14260 17141 14263
rect 15252 14232 17141 14260
rect 15252 14220 15258 14232
rect 17129 14229 17141 14232
rect 17175 14229 17187 14263
rect 17129 14223 17187 14229
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 2038 14056 2044 14068
rect 1999 14028 2044 14056
rect 2038 14016 2044 14028
rect 2096 14016 2102 14068
rect 3326 14056 3332 14068
rect 2700 14028 3332 14056
rect 2498 13880 2504 13932
rect 2556 13920 2562 13932
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 2556 13892 2605 13920
rect 2556 13880 2562 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 2700 13852 2728 14028
rect 3326 14016 3332 14028
rect 3384 14056 3390 14068
rect 3786 14056 3792 14068
rect 3384 14028 3792 14056
rect 3384 14016 3390 14028
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 4706 14056 4712 14068
rect 4667 14028 4712 14056
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 5408 14028 6837 14056
rect 5408 14016 5414 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 6825 14019 6883 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 10686 14056 10692 14068
rect 8496 14028 10692 14056
rect 3697 13991 3755 13997
rect 3697 13957 3709 13991
rect 3743 13988 3755 13991
rect 3743 13960 5488 13988
rect 3743 13957 3755 13960
rect 3697 13951 3755 13957
rect 3786 13880 3792 13932
rect 3844 13920 3850 13932
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 3844 13892 4261 13920
rect 3844 13880 3850 13892
rect 4249 13889 4261 13892
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13889 5411 13923
rect 5460 13920 5488 13960
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 5721 13991 5779 13997
rect 5721 13988 5733 13991
rect 5592 13960 5733 13988
rect 5592 13948 5598 13960
rect 5721 13957 5733 13960
rect 5767 13957 5779 13991
rect 8496 13988 8524 14028
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 16724 14028 17509 14056
rect 16724 14016 16730 14028
rect 17497 14025 17509 14028
rect 17543 14025 17555 14059
rect 17497 14019 17555 14025
rect 10137 13991 10195 13997
rect 10137 13988 10149 13991
rect 5721 13951 5779 13957
rect 6196 13960 8524 13988
rect 8588 13960 10149 13988
rect 6196 13920 6224 13960
rect 5460 13892 6224 13920
rect 6365 13923 6423 13929
rect 5353 13883 5411 13889
rect 6365 13889 6377 13923
rect 6411 13920 6423 13923
rect 6454 13920 6460 13932
rect 6411 13892 6460 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 2516 13824 2728 13852
rect 2516 13793 2544 13824
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 3016 13824 4169 13852
rect 3016 13812 3022 13824
rect 4157 13821 4169 13824
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 4798 13812 4804 13864
rect 4856 13852 4862 13864
rect 5169 13855 5227 13861
rect 5169 13852 5181 13855
rect 4856 13824 5181 13852
rect 4856 13812 4862 13824
rect 5169 13821 5181 13824
rect 5215 13821 5227 13855
rect 5368 13852 5396 13883
rect 6380 13852 6408 13883
rect 6454 13880 6460 13892
rect 6512 13880 6518 13932
rect 7466 13920 7472 13932
rect 7427 13892 7472 13920
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 8588 13929 8616 13960
rect 10137 13957 10149 13960
rect 10183 13957 10195 13991
rect 10137 13951 10195 13957
rect 14185 13991 14243 13997
rect 14185 13957 14197 13991
rect 14231 13988 14243 13991
rect 14366 13988 14372 14000
rect 14231 13960 14372 13988
rect 14231 13957 14243 13960
rect 14185 13951 14243 13957
rect 14366 13948 14372 13960
rect 14424 13948 14430 14000
rect 18233 13991 18291 13997
rect 14568 13960 15516 13988
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8754 13920 8760 13932
rect 8715 13892 8760 13920
rect 8573 13883 8631 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 9272 13892 9689 13920
rect 9272 13880 9278 13892
rect 9677 13889 9689 13892
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 11514 13920 11520 13932
rect 10827 13892 11520 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13920 13783 13923
rect 14274 13920 14280 13932
rect 13771 13892 14280 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14274 13880 14280 13892
rect 14332 13920 14338 13932
rect 14568 13920 14596 13960
rect 14734 13920 14740 13932
rect 14332 13892 14596 13920
rect 14695 13892 14740 13920
rect 14332 13880 14338 13892
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 5368 13824 6408 13852
rect 7285 13855 7343 13861
rect 5169 13815 5227 13821
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 8662 13852 8668 13864
rect 7331 13824 8668 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 8662 13812 8668 13824
rect 8720 13812 8726 13864
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9398 13852 9404 13864
rect 8904 13824 9404 13852
rect 8904 13812 8910 13824
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 10597 13855 10655 13861
rect 10597 13852 10609 13855
rect 9640 13824 10609 13852
rect 9640 13812 9646 13824
rect 10597 13821 10609 13824
rect 10643 13821 10655 13855
rect 10597 13815 10655 13821
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12768 13824 12817 13852
rect 12768 13812 12774 13824
rect 12805 13821 12817 13824
rect 12851 13852 12863 13855
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12851 13824 13001 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 12989 13821 13001 13824
rect 13035 13821 13047 13855
rect 13354 13852 13360 13864
rect 13315 13824 13360 13852
rect 12989 13815 13047 13821
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13852 14703 13855
rect 15378 13852 15384 13864
rect 14691 13824 15384 13852
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15488 13861 15516 13960
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18506 13988 18512 14000
rect 18279 13960 18512 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16574 13920 16580 13932
rect 16071 13892 16580 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17218 13920 17224 13932
rect 17083 13892 17224 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 15488 13855 15566 13861
rect 15488 13824 15520 13855
rect 15508 13821 15520 13824
rect 15554 13821 15566 13855
rect 15508 13815 15566 13821
rect 17313 13855 17371 13861
rect 17313 13821 17325 13855
rect 17359 13852 17371 13855
rect 17678 13852 17684 13864
rect 17359 13824 17684 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 2501 13787 2559 13793
rect 2501 13753 2513 13787
rect 2547 13753 2559 13787
rect 2501 13747 2559 13753
rect 4065 13787 4123 13793
rect 4065 13753 4077 13787
rect 4111 13784 4123 13787
rect 4246 13784 4252 13796
rect 4111 13756 4252 13784
rect 4111 13753 4123 13756
rect 4065 13747 4123 13753
rect 4246 13744 4252 13756
rect 4304 13744 4310 13796
rect 4706 13744 4712 13796
rect 4764 13784 4770 13796
rect 4764 13756 5764 13784
rect 4764 13744 4770 13756
rect 1394 13676 1400 13728
rect 1452 13716 1458 13728
rect 2409 13719 2467 13725
rect 2409 13716 2421 13719
rect 1452 13688 2421 13716
rect 1452 13676 1458 13688
rect 2409 13685 2421 13688
rect 2455 13685 2467 13719
rect 2409 13679 2467 13685
rect 5077 13719 5135 13725
rect 5077 13685 5089 13719
rect 5123 13716 5135 13719
rect 5626 13716 5632 13728
rect 5123 13688 5632 13716
rect 5123 13685 5135 13688
rect 5077 13679 5135 13685
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 5736 13716 5764 13756
rect 5810 13744 5816 13796
rect 5868 13784 5874 13796
rect 6730 13784 6736 13796
rect 5868 13756 6736 13784
rect 5868 13744 5874 13756
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 9306 13784 9312 13796
rect 6840 13756 9312 13784
rect 6086 13716 6092 13728
rect 5736 13688 6092 13716
rect 6086 13676 6092 13688
rect 6144 13676 6150 13728
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 6236 13688 6281 13716
rect 6236 13676 6242 13688
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6840 13716 6868 13756
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 6420 13688 6868 13716
rect 7193 13719 7251 13725
rect 6420 13676 6426 13688
rect 7193 13685 7205 13719
rect 7239 13716 7251 13719
rect 7834 13716 7840 13728
rect 7239 13688 7840 13716
rect 7239 13685 7251 13688
rect 7193 13679 7251 13685
rect 7834 13676 7840 13688
rect 7892 13676 7898 13728
rect 8478 13716 8484 13728
rect 8439 13688 8484 13716
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 9122 13716 9128 13728
rect 9083 13688 9128 13716
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9416 13716 9444 13812
rect 9493 13787 9551 13793
rect 9493 13753 9505 13787
rect 9539 13784 9551 13787
rect 9674 13784 9680 13796
rect 9539 13756 9680 13784
rect 9539 13753 9551 13756
rect 9493 13747 9551 13753
rect 9674 13744 9680 13756
rect 9732 13744 9738 13796
rect 16022 13784 16028 13796
rect 14108 13756 16028 13784
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 9416 13688 9597 13716
rect 9585 13685 9597 13688
rect 9631 13685 9643 13719
rect 10502 13716 10508 13728
rect 10463 13688 10508 13716
rect 9585 13679 9643 13685
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 12342 13676 12348 13728
rect 12400 13716 12406 13728
rect 14108 13716 14136 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 16117 13787 16175 13793
rect 16117 13753 16129 13787
rect 16163 13753 16175 13787
rect 16117 13747 16175 13753
rect 12400 13688 14136 13716
rect 12400 13676 12406 13688
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 14553 13719 14611 13725
rect 14553 13716 14565 13719
rect 14240 13688 14565 13716
rect 14240 13676 14246 13688
rect 14553 13685 14565 13688
rect 14599 13685 14611 13719
rect 14553 13679 14611 13685
rect 15611 13719 15669 13725
rect 15611 13685 15623 13719
rect 15657 13716 15669 13719
rect 16132 13716 16160 13747
rect 15657 13688 16160 13716
rect 15657 13685 15669 13688
rect 15611 13679 15669 13685
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 2222 13512 2228 13524
rect 1995 13484 2228 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 2774 13512 2780 13524
rect 2363 13484 2780 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2774 13472 2780 13484
rect 2832 13512 2838 13524
rect 2961 13515 3019 13521
rect 2832 13484 2925 13512
rect 2832 13472 2838 13484
rect 2884 13444 2912 13484
rect 2961 13481 2973 13515
rect 3007 13512 3019 13515
rect 3418 13512 3424 13524
rect 3007 13484 3424 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 5166 13512 5172 13524
rect 4847 13484 5172 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5813 13515 5871 13521
rect 5813 13481 5825 13515
rect 5859 13512 5871 13515
rect 6178 13512 6184 13524
rect 5859 13484 6184 13512
rect 5859 13481 5871 13484
rect 5813 13475 5871 13481
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 7466 13512 7472 13524
rect 6472 13484 7472 13512
rect 6270 13444 6276 13456
rect 2884 13416 6276 13444
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 6362 13404 6368 13456
rect 6420 13404 6426 13456
rect 1670 13336 1676 13388
rect 1728 13376 1734 13388
rect 2409 13379 2467 13385
rect 2409 13376 2421 13379
rect 1728 13348 2421 13376
rect 1728 13336 1734 13348
rect 2409 13345 2421 13348
rect 2455 13376 2467 13379
rect 2590 13376 2596 13388
rect 2455 13348 2596 13376
rect 2455 13345 2467 13348
rect 2409 13339 2467 13345
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 3142 13336 3148 13388
rect 3200 13376 3206 13388
rect 3329 13379 3387 13385
rect 3329 13376 3341 13379
rect 3200 13348 3341 13376
rect 3200 13336 3206 13348
rect 3329 13345 3341 13348
rect 3375 13345 3387 13379
rect 5166 13376 5172 13388
rect 5127 13348 5172 13376
rect 3329 13339 3387 13345
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 6380 13376 6408 13404
rect 6227 13348 6408 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 2556 13280 2601 13308
rect 2556 13268 2562 13280
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 2832 13280 3433 13308
rect 2832 13268 2838 13280
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 2516 13240 2544 13268
rect 3528 13240 3556 13271
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 5261 13311 5319 13317
rect 5261 13308 5273 13311
rect 4948 13280 5273 13308
rect 4948 13268 4954 13280
rect 5261 13277 5273 13280
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13277 5503 13311
rect 5445 13271 5503 13277
rect 2516 13212 3556 13240
rect 3694 13200 3700 13252
rect 3752 13240 3758 13252
rect 4706 13240 4712 13252
rect 3752 13212 4712 13240
rect 3752 13200 3758 13212
rect 4706 13200 4712 13212
rect 4764 13200 4770 13252
rect 5460 13240 5488 13271
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6472 13317 6500 13484
rect 7466 13472 7472 13484
rect 7524 13512 7530 13524
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 7524 13484 8217 13512
rect 7524 13472 7530 13484
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 8205 13475 8263 13481
rect 8941 13515 8999 13521
rect 8941 13481 8953 13515
rect 8987 13512 8999 13515
rect 9122 13512 9128 13524
rect 8987 13484 9128 13512
rect 8987 13481 8999 13484
rect 8941 13475 8999 13481
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 13262 13512 13268 13524
rect 9364 13484 13268 13512
rect 9364 13472 9370 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 14182 13512 14188 13524
rect 14143 13484 14188 13512
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 14553 13515 14611 13521
rect 14553 13481 14565 13515
rect 14599 13512 14611 13515
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 14599 13484 15301 13512
rect 14599 13481 14611 13484
rect 14553 13475 14611 13481
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15436 13484 16313 13512
rect 15436 13472 15442 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 17313 13515 17371 13521
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17586 13512 17592 13524
rect 17359 13484 17592 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17586 13472 17592 13484
rect 17644 13472 17650 13524
rect 6730 13404 6736 13456
rect 6788 13444 6794 13456
rect 7092 13447 7150 13453
rect 6788 13416 7052 13444
rect 6788 13404 6794 13416
rect 7024 13376 7052 13416
rect 7092 13413 7104 13447
rect 7138 13444 7150 13447
rect 7742 13444 7748 13456
rect 7138 13416 7748 13444
rect 7138 13413 7150 13416
rect 7092 13407 7150 13413
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 10134 13444 10140 13456
rect 8168 13416 10140 13444
rect 8168 13404 8174 13416
rect 10134 13404 10140 13416
rect 10192 13404 10198 13456
rect 10318 13444 10324 13456
rect 10279 13416 10324 13444
rect 10318 13404 10324 13416
rect 10376 13404 10382 13456
rect 10686 13404 10692 13456
rect 10744 13444 10750 13456
rect 10744 13416 12020 13444
rect 10744 13404 10750 13416
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 7024 13348 9413 13376
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 10244 13348 10732 13376
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6052 13280 6285 13308
rect 6052 13268 6058 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6696 13280 6837 13308
rect 6696 13268 6702 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 9030 13308 9036 13320
rect 8991 13280 9036 13308
rect 6825 13271 6883 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 9180 13280 9225 13308
rect 9180 13268 9186 13280
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 10244 13308 10272 13348
rect 10410 13308 10416 13320
rect 9548 13280 10272 13308
rect 10371 13280 10416 13308
rect 9548 13268 9554 13280
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 10594 13308 10600 13320
rect 10555 13280 10600 13308
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 10704 13308 10732 13348
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 10928 13348 11345 13376
rect 10928 13336 10934 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 11425 13379 11483 13385
rect 11425 13345 11437 13379
rect 11471 13376 11483 13379
rect 11606 13376 11612 13388
rect 11471 13348 11612 13376
rect 11471 13345 11483 13348
rect 11425 13339 11483 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 11992 13385 12020 13416
rect 12158 13404 12164 13456
rect 12216 13444 12222 13456
rect 12253 13447 12311 13453
rect 12253 13444 12265 13447
rect 12216 13416 12265 13444
rect 12216 13404 12222 13416
rect 12253 13413 12265 13416
rect 12299 13413 12311 13447
rect 12253 13407 12311 13413
rect 16022 13404 16028 13456
rect 16080 13444 16086 13456
rect 17770 13444 17776 13456
rect 16080 13416 17776 13444
rect 16080 13404 16086 13416
rect 17770 13404 17776 13416
rect 17828 13404 17834 13456
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13345 12035 13379
rect 11977 13339 12035 13345
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13376 13599 13379
rect 13998 13376 14004 13388
rect 13587 13348 14004 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14516 13348 15669 13376
rect 14516 13336 14522 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16298 13376 16304 13388
rect 15804 13348 16304 13376
rect 15804 13336 15810 13348
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 16669 13379 16727 13385
rect 16669 13376 16681 13379
rect 16632 13348 16681 13376
rect 16632 13336 16638 13348
rect 16669 13345 16681 13348
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 17586 13336 17592 13388
rect 17644 13376 17650 13388
rect 17681 13379 17739 13385
rect 17681 13376 17693 13379
rect 17644 13348 17693 13376
rect 17644 13336 17650 13348
rect 17681 13345 17693 13348
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 11514 13308 11520 13320
rect 10704 13280 11376 13308
rect 11475 13280 11520 13308
rect 5718 13240 5724 13252
rect 5460 13212 5724 13240
rect 5718 13200 5724 13212
rect 5776 13240 5782 13252
rect 9401 13243 9459 13249
rect 5776 13212 6500 13240
rect 5776 13200 5782 13212
rect 6472 13184 6500 13212
rect 9401 13209 9413 13243
rect 9447 13240 9459 13243
rect 11146 13240 11152 13252
rect 9447 13212 11152 13240
rect 9447 13209 9459 13212
rect 9401 13203 9459 13209
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 11348 13240 11376 13280
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 13630 13308 13636 13320
rect 13591 13280 13636 13308
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 14645 13311 14703 13317
rect 13780 13280 13825 13308
rect 13780 13268 13786 13280
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14826 13308 14832 13320
rect 14787 13280 14832 13308
rect 14645 13271 14703 13277
rect 14550 13240 14556 13252
rect 11348 13212 14556 13240
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 14660 13240 14688 13271
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16206 13308 16212 13320
rect 15979 13280 16212 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 15286 13240 15292 13252
rect 14660 13212 15292 13240
rect 15286 13200 15292 13212
rect 15344 13200 15350 13252
rect 16298 13200 16304 13252
rect 16356 13240 16362 13252
rect 16868 13240 16896 13271
rect 16356 13212 16896 13240
rect 16356 13200 16362 13212
rect 17586 13200 17592 13252
rect 17644 13240 17650 13252
rect 17880 13240 17908 13271
rect 17644 13212 17908 13240
rect 17644 13200 17650 13212
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 4614 13172 4620 13184
rect 2280 13144 4620 13172
rect 2280 13132 2286 13144
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 6454 13132 6460 13184
rect 6512 13172 6518 13184
rect 8202 13172 8208 13184
rect 6512 13144 8208 13172
rect 6512 13132 6518 13144
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 8573 13175 8631 13181
rect 8573 13172 8585 13175
rect 8352 13144 8585 13172
rect 8352 13132 8358 13144
rect 8573 13141 8585 13144
rect 8619 13141 8631 13175
rect 8573 13135 8631 13141
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9824 13144 9965 13172
rect 9824 13132 9830 13144
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 9953 13135 10011 13141
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10965 13175 11023 13181
rect 10965 13172 10977 13175
rect 10284 13144 10977 13172
rect 10284 13132 10290 13144
rect 10965 13141 10977 13144
rect 11011 13141 11023 13175
rect 10965 13135 11023 13141
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 16482 13172 16488 13184
rect 13219 13144 16488 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 3050 12968 3056 12980
rect 1903 12940 3056 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 3844 12940 4261 12968
rect 3844 12928 3850 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 4249 12931 4307 12937
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 11149 12971 11207 12977
rect 11149 12968 11161 12971
rect 10468 12940 11161 12968
rect 10468 12928 10474 12940
rect 11149 12937 11161 12940
rect 11195 12937 11207 12971
rect 14550 12968 14556 12980
rect 11149 12931 11207 12937
rect 12452 12940 14556 12968
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 6454 12900 6460 12912
rect 4672 12872 6460 12900
rect 4672 12860 4678 12872
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 8202 12900 8208 12912
rect 8163 12872 8208 12900
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 9490 12860 9496 12912
rect 9548 12900 9554 12912
rect 12452 12900 12480 12940
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 16298 12968 16304 12980
rect 14884 12940 16304 12968
rect 14884 12928 14890 12940
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 16574 12968 16580 12980
rect 16535 12940 16580 12968
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 9548 12872 12480 12900
rect 9548 12860 9554 12872
rect 13446 12860 13452 12912
rect 13504 12900 13510 12912
rect 13817 12903 13875 12909
rect 13817 12900 13829 12903
rect 13504 12872 13829 12900
rect 13504 12860 13510 12872
rect 13817 12869 13829 12872
rect 13863 12869 13875 12903
rect 13817 12863 13875 12869
rect 2406 12832 2412 12844
rect 2367 12804 2412 12832
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5442 12832 5448 12844
rect 5307 12804 5448 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5442 12792 5448 12804
rect 5500 12832 5506 12844
rect 5718 12832 5724 12844
rect 5500 12804 5724 12832
rect 5500 12792 5506 12804
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 10778 12832 10784 12844
rect 10691 12804 10784 12832
rect 6365 12795 6423 12801
rect 2222 12764 2228 12776
rect 2183 12736 2228 12764
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 3694 12764 3700 12776
rect 2915 12736 3700 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 5350 12764 5356 12776
rect 5215 12736 5356 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 3136 12699 3194 12705
rect 3136 12665 3148 12699
rect 3182 12696 3194 12699
rect 3602 12696 3608 12708
rect 3182 12668 3608 12696
rect 3182 12665 3194 12668
rect 3136 12659 3194 12665
rect 3602 12656 3608 12668
rect 3660 12696 3666 12708
rect 5077 12699 5135 12705
rect 3660 12668 4936 12696
rect 3660 12656 3666 12668
rect 2314 12588 2320 12640
rect 2372 12628 2378 12640
rect 4706 12628 4712 12640
rect 2372 12600 2417 12628
rect 4667 12600 4712 12628
rect 2372 12588 2378 12600
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 4908 12628 4936 12668
rect 5077 12665 5089 12699
rect 5123 12696 5135 12699
rect 6089 12699 6147 12705
rect 5123 12668 5764 12696
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 5258 12628 5264 12640
rect 4908 12600 5264 12628
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5736 12637 5764 12668
rect 6089 12665 6101 12699
rect 6135 12696 6147 12699
rect 6380 12696 6408 12795
rect 10778 12792 10784 12804
rect 10836 12832 10842 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 10836 12804 11713 12832
rect 10836 12792 10842 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 14458 12832 14464 12844
rect 14419 12804 14464 12832
rect 11701 12795 11759 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 16206 12832 16212 12844
rect 15988 12804 16212 12832
rect 15988 12792 15994 12804
rect 16206 12792 16212 12804
rect 16264 12832 16270 12844
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 16264 12804 17233 12832
rect 16264 12792 16270 12804
rect 17221 12801 17233 12804
rect 17267 12832 17279 12835
rect 17770 12832 17776 12844
rect 17267 12804 17776 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 6638 12724 6644 12776
rect 6696 12764 6702 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6696 12736 6837 12764
rect 6696 12724 6702 12736
rect 6825 12733 6837 12736
rect 6871 12764 6883 12767
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 6871 12736 8493 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 8481 12733 8493 12736
rect 8527 12733 8539 12767
rect 8481 12727 8539 12733
rect 8748 12767 8806 12773
rect 8748 12733 8760 12767
rect 8794 12764 8806 12767
rect 9214 12764 9220 12776
rect 8794 12736 9220 12764
rect 8794 12733 8806 12736
rect 8748 12727 8806 12733
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 10060 12736 10517 12764
rect 7092 12699 7150 12705
rect 7092 12696 7104 12699
rect 6135 12668 6316 12696
rect 6380 12668 7104 12696
rect 6135 12665 6147 12668
rect 6089 12659 6147 12665
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12597 5779 12631
rect 5721 12591 5779 12597
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 6181 12631 6239 12637
rect 6181 12628 6193 12631
rect 5868 12600 6193 12628
rect 5868 12588 5874 12600
rect 6181 12597 6193 12600
rect 6227 12597 6239 12631
rect 6288 12628 6316 12668
rect 7092 12665 7104 12668
rect 7138 12696 7150 12699
rect 7466 12696 7472 12708
rect 7138 12668 7472 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 10060 12696 10088 12736
rect 10505 12733 10517 12736
rect 10551 12764 10563 12767
rect 10962 12764 10968 12776
rect 10551 12736 10968 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 12342 12764 12348 12776
rect 11348 12736 12348 12764
rect 8128 12668 10088 12696
rect 8128 12628 8156 12668
rect 10318 12656 10324 12708
rect 10376 12696 10382 12708
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10376 12668 10609 12696
rect 10376 12656 10382 12668
rect 10597 12665 10609 12668
rect 10643 12665 10655 12699
rect 10597 12659 10655 12665
rect 6288 12600 8156 12628
rect 6181 12591 6239 12597
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 9122 12628 9128 12640
rect 8444 12600 9128 12628
rect 8444 12588 8450 12600
rect 9122 12588 9128 12600
rect 9180 12628 9186 12640
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 9180 12600 9873 12628
rect 9180 12588 9186 12600
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 10137 12631 10195 12637
rect 10137 12597 10149 12631
rect 10183 12628 10195 12631
rect 10226 12628 10232 12640
rect 10183 12600 10232 12628
rect 10183 12597 10195 12600
rect 10137 12591 10195 12597
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 10410 12588 10416 12640
rect 10468 12628 10474 12640
rect 11348 12628 11376 12736
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 12526 12764 12532 12776
rect 12483 12736 12532 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 12704 12767 12762 12773
rect 12704 12733 12716 12767
rect 12750 12764 12762 12767
rect 14642 12764 14648 12776
rect 12750 12736 14648 12764
rect 12750 12733 12762 12736
rect 12704 12727 12762 12733
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 14734 12724 14740 12776
rect 14792 12764 14798 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14792 12736 14933 12764
rect 14792 12724 14798 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 15188 12767 15246 12773
rect 15188 12733 15200 12767
rect 15234 12764 15246 12767
rect 15948 12764 15976 12792
rect 15234 12736 15976 12764
rect 15234 12733 15246 12736
rect 15188 12727 15246 12733
rect 11422 12656 11428 12708
rect 11480 12696 11486 12708
rect 11609 12699 11667 12705
rect 11609 12696 11621 12699
rect 11480 12668 11621 12696
rect 11480 12656 11486 12668
rect 11609 12665 11621 12668
rect 11655 12665 11667 12699
rect 11609 12659 11667 12665
rect 14274 12656 14280 12708
rect 14332 12696 14338 12708
rect 16850 12696 16856 12708
rect 14332 12668 16856 12696
rect 14332 12656 14338 12668
rect 16850 12656 16856 12668
rect 16908 12696 16914 12708
rect 16945 12699 17003 12705
rect 16945 12696 16957 12699
rect 16908 12668 16957 12696
rect 16908 12656 16914 12668
rect 16945 12665 16957 12668
rect 16991 12665 17003 12699
rect 16945 12659 17003 12665
rect 11514 12628 11520 12640
rect 10468 12600 11376 12628
rect 11475 12600 11520 12628
rect 10468 12588 10474 12600
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 17092 12600 17137 12628
rect 17092 12588 17098 12600
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2314 12424 2320 12436
rect 1995 12396 2320 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 2958 12424 2964 12436
rect 2919 12396 2964 12424
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3421 12427 3479 12433
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 4706 12424 4712 12436
rect 3467 12396 4712 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 5316 12396 5457 12424
rect 5316 12384 5322 12396
rect 5445 12393 5457 12396
rect 5491 12393 5503 12427
rect 5445 12387 5503 12393
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 5721 12427 5779 12433
rect 5721 12424 5733 12427
rect 5684 12396 5733 12424
rect 5684 12384 5690 12396
rect 5721 12393 5733 12396
rect 5767 12393 5779 12427
rect 5721 12387 5779 12393
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 8021 12427 8079 12433
rect 6512 12396 7604 12424
rect 6512 12384 6518 12396
rect 4154 12356 4160 12368
rect 2332 12328 4160 12356
rect 2332 12297 2360 12328
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 4332 12359 4390 12365
rect 4332 12325 4344 12359
rect 4378 12356 4390 12359
rect 5350 12356 5356 12368
rect 4378 12328 5356 12356
rect 4378 12325 4390 12328
rect 4332 12319 4390 12325
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 5902 12316 5908 12368
rect 5960 12356 5966 12368
rect 6086 12356 6092 12368
rect 5960 12328 6092 12356
rect 5960 12316 5966 12328
rect 6086 12316 6092 12328
rect 6144 12356 6150 12368
rect 7576 12356 7604 12396
rect 8021 12393 8033 12427
rect 8067 12424 8079 12427
rect 8481 12427 8539 12433
rect 8481 12424 8493 12427
rect 8067 12396 8493 12424
rect 8067 12393 8079 12396
rect 8021 12387 8079 12393
rect 8481 12393 8493 12396
rect 8527 12393 8539 12427
rect 8481 12387 8539 12393
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 9030 12424 9036 12436
rect 8619 12396 9036 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10594 12424 10600 12436
rect 9876 12396 10600 12424
rect 7650 12356 7656 12368
rect 6144 12328 7052 12356
rect 7576 12328 7656 12356
rect 6144 12316 6150 12328
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12257 2375 12291
rect 2317 12251 2375 12257
rect 2409 12291 2467 12297
rect 2409 12257 2421 12291
rect 2455 12288 2467 12291
rect 2498 12288 2504 12300
rect 2455 12260 2504 12288
rect 2455 12257 2467 12260
rect 2409 12251 2467 12257
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 5534 12288 5540 12300
rect 3375 12260 5540 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6472 12260 6929 12288
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3602 12220 3608 12232
rect 3563 12192 3608 12220
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3752 12192 4077 12220
rect 3752 12180 3758 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 6178 12084 6184 12096
rect 3476 12056 6184 12084
rect 3476 12044 3482 12056
rect 6178 12044 6184 12056
rect 6236 12084 6242 12096
rect 6472 12084 6500 12260
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 7024 12288 7052 12328
rect 7650 12316 7656 12328
rect 7708 12316 7714 12368
rect 7929 12359 7987 12365
rect 7929 12325 7941 12359
rect 7975 12356 7987 12359
rect 9766 12356 9772 12368
rect 7975 12328 9772 12356
rect 7975 12325 7987 12328
rect 7929 12319 7987 12325
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 8941 12291 8999 12297
rect 8941 12288 8953 12291
rect 7024 12260 8953 12288
rect 6917 12251 6975 12257
rect 8941 12257 8953 12260
rect 8987 12288 8999 12291
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 8987 12260 9413 12288
rect 8987 12257 8999 12260
rect 8941 12251 8999 12257
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 7006 12220 7012 12232
rect 6967 12192 7012 12220
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7282 12220 7288 12232
rect 7239 12192 7288 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 8110 12220 8116 12232
rect 8071 12192 8116 12220
rect 8110 12180 8116 12192
rect 8168 12220 8174 12232
rect 8386 12220 8392 12232
rect 8168 12192 8392 12220
rect 8168 12180 8174 12192
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 9030 12220 9036 12232
rect 8991 12192 9036 12220
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 9214 12220 9220 12232
rect 9127 12192 9220 12220
rect 9214 12180 9220 12192
rect 9272 12220 9278 12232
rect 9876 12220 9904 12396
rect 10594 12384 10600 12396
rect 10652 12424 10658 12436
rect 11609 12427 11667 12433
rect 11609 12424 11621 12427
rect 10652 12396 11621 12424
rect 10652 12384 10658 12396
rect 11609 12393 11621 12396
rect 11655 12393 11667 12427
rect 14458 12424 14464 12436
rect 11609 12387 11667 12393
rect 13096 12396 14464 12424
rect 10496 12359 10554 12365
rect 10496 12325 10508 12359
rect 10542 12356 10554 12359
rect 10778 12356 10784 12368
rect 10542 12328 10784 12356
rect 10542 12325 10554 12328
rect 10496 12319 10554 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 13096 12356 13124 12396
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 14642 12424 14648 12436
rect 14603 12396 14648 12424
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 12032 12328 13124 12356
rect 13532 12359 13590 12365
rect 12032 12316 12038 12328
rect 13532 12325 13544 12359
rect 13578 12356 13590 12359
rect 14734 12356 14740 12368
rect 13578 12328 14740 12356
rect 13578 12325 13590 12328
rect 13532 12319 13590 12325
rect 14734 12316 14740 12328
rect 14792 12316 14798 12368
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 16298 12356 16304 12368
rect 15804 12328 16304 12356
rect 15804 12316 15810 12328
rect 16298 12316 16304 12328
rect 16356 12316 16362 12368
rect 12158 12288 12164 12300
rect 9272 12192 9904 12220
rect 9968 12260 12164 12288
rect 9272 12180 9278 12192
rect 9401 12155 9459 12161
rect 9401 12121 9413 12155
rect 9447 12152 9459 12155
rect 9968 12152 9996 12260
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12288 12679 12291
rect 14090 12288 14096 12300
rect 12667 12260 14096 12288
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14274 12248 14280 12300
rect 14332 12288 14338 12300
rect 14550 12288 14556 12300
rect 14332 12260 14556 12288
rect 14332 12248 14338 12260
rect 14550 12248 14556 12260
rect 14608 12288 14614 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14608 12260 15669 12288
rect 14608 12248 14614 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15838 12288 15844 12300
rect 15657 12251 15715 12257
rect 15764 12260 15844 12288
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 12710 12220 12716 12232
rect 12671 12192 12716 12220
rect 10229 12183 10287 12189
rect 9447 12124 9996 12152
rect 9447 12121 9459 12124
rect 9401 12115 9459 12121
rect 6236 12056 6500 12084
rect 6549 12087 6607 12093
rect 6236 12044 6242 12056
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 7374 12084 7380 12096
rect 6595 12056 7380 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7561 12087 7619 12093
rect 7561 12053 7573 12087
rect 7607 12084 7619 12087
rect 8018 12084 8024 12096
rect 7607 12056 8024 12084
rect 7607 12053 7619 12056
rect 7561 12047 7619 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 9306 12084 9312 12096
rect 8527 12056 9312 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 10244 12084 10272 12183
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 10410 12084 10416 12096
rect 10244 12056 10416 12084
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 11756 12056 12265 12084
rect 11756 12044 11762 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12912 12084 12940 12183
rect 13170 12180 13176 12232
rect 13228 12220 13234 12232
rect 15764 12229 15792 12260
rect 15838 12248 15844 12260
rect 15896 12288 15902 12300
rect 16482 12288 16488 12300
rect 15896 12260 16488 12288
rect 15896 12248 15902 12260
rect 16482 12248 16488 12260
rect 16540 12248 16546 12300
rect 16660 12291 16718 12297
rect 16660 12257 16672 12291
rect 16706 12288 16718 12291
rect 16942 12288 16948 12300
rect 16706 12260 16948 12288
rect 16706 12257 16718 12260
rect 16660 12251 16718 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 13228 12192 13277 12220
rect 13228 12180 13234 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15930 12220 15936 12232
rect 15891 12192 15936 12220
rect 15749 12183 15807 12189
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 15286 12112 15292 12164
rect 15344 12152 15350 12164
rect 16408 12152 16436 12183
rect 15344 12124 16436 12152
rect 15344 12112 15350 12124
rect 13906 12084 13912 12096
rect 12912 12056 13912 12084
rect 12253 12047 12311 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 17770 12084 17776 12096
rect 17731 12056 17776 12084
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 2685 11883 2743 11889
rect 2685 11849 2697 11883
rect 2731 11880 2743 11883
rect 2774 11880 2780 11892
rect 2731 11852 2780 11880
rect 2731 11849 2743 11852
rect 2685 11843 2743 11849
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 3513 11883 3571 11889
rect 3513 11849 3525 11883
rect 3559 11880 3571 11883
rect 6454 11880 6460 11892
rect 3559 11852 6460 11880
rect 3559 11849 3571 11852
rect 3513 11843 3571 11849
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 9306 11880 9312 11892
rect 9267 11852 9312 11880
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 11606 11880 11612 11892
rect 9548 11852 11612 11880
rect 9548 11840 9554 11852
rect 11606 11840 11612 11852
rect 11664 11840 11670 11892
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 12768 11852 13093 11880
rect 12768 11840 12774 11852
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 13722 11880 13728 11892
rect 13081 11843 13139 11849
rect 13280 11852 13728 11880
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11812 1731 11815
rect 3142 11812 3148 11824
rect 1719 11784 3148 11812
rect 1719 11781 1731 11784
rect 1673 11775 1731 11781
rect 3142 11772 3148 11784
rect 3200 11772 3206 11824
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 7466 11812 7472 11824
rect 4764 11784 7472 11812
rect 4764 11772 4770 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 13280 11812 13308 11852
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 14090 11880 14096 11892
rect 14051 11852 14096 11880
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14458 11840 14464 11892
rect 14516 11880 14522 11892
rect 14516 11852 15332 11880
rect 14516 11840 14522 11852
rect 10980 11784 13308 11812
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2590 11744 2596 11756
rect 2363 11716 2596 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2590 11704 2596 11716
rect 2648 11744 2654 11756
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 2648 11716 3341 11744
rect 2648 11704 2654 11716
rect 3329 11713 3341 11716
rect 3375 11744 3387 11747
rect 3605 11747 3663 11753
rect 3605 11744 3617 11747
rect 3375 11716 3617 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3605 11713 3617 11716
rect 3651 11713 3663 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 3605 11707 3663 11713
rect 6288 11716 6377 11744
rect 6288 11688 6316 11716
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 10980 11753 11008 11784
rect 13354 11772 13360 11824
rect 13412 11812 13418 11824
rect 15194 11812 15200 11824
rect 13412 11784 15200 11812
rect 13412 11772 13418 11784
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 9861 11747 9919 11753
rect 9861 11744 9873 11747
rect 9272 11716 9873 11744
rect 9272 11704 9278 11716
rect 9861 11713 9873 11716
rect 9907 11713 9919 11747
rect 9861 11707 9919 11713
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 13446 11744 13452 11756
rect 12023 11716 13452 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 13538 11704 13544 11756
rect 13596 11744 13602 11756
rect 13725 11747 13783 11753
rect 13596 11716 13641 11744
rect 13596 11704 13602 11716
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 13814 11744 13820 11756
rect 13771 11716 13820 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 13814 11704 13820 11716
rect 13872 11744 13878 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 13872 11716 14657 11744
rect 13872 11704 13878 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 15304 11744 15332 11852
rect 15304 11716 15516 11744
rect 14645 11707 14703 11713
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11676 2099 11679
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 2087 11648 3525 11676
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3694 11676 3700 11688
rect 3655 11648 3700 11676
rect 3513 11639 3571 11645
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 3786 11636 3792 11688
rect 3844 11676 3850 11688
rect 3953 11679 4011 11685
rect 3953 11676 3965 11679
rect 3844 11648 3965 11676
rect 3844 11636 3850 11648
rect 3953 11645 3965 11648
rect 3999 11645 4011 11679
rect 3953 11639 4011 11645
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 6089 11679 6147 11685
rect 6089 11676 6101 11679
rect 4396 11648 6101 11676
rect 4396 11636 4402 11648
rect 6089 11645 6101 11648
rect 6135 11645 6147 11679
rect 6089 11639 6147 11645
rect 6270 11636 6276 11688
rect 6328 11636 6334 11688
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 7469 11679 7527 11685
rect 7469 11676 7481 11679
rect 7248 11648 7481 11676
rect 7248 11636 7254 11648
rect 7469 11645 7481 11648
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7828 11679 7886 11685
rect 7828 11645 7840 11679
rect 7874 11676 7886 11679
rect 8110 11676 8116 11688
rect 7874 11648 8116 11676
rect 7874 11645 7886 11648
rect 7828 11639 7886 11645
rect 3053 11611 3111 11617
rect 3053 11577 3065 11611
rect 3099 11608 3111 11611
rect 3418 11608 3424 11620
rect 3099 11580 3424 11608
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 6181 11611 6239 11617
rect 6181 11608 6193 11611
rect 4764 11580 6193 11608
rect 4764 11568 4770 11580
rect 6181 11577 6193 11580
rect 6227 11577 6239 11611
rect 6181 11571 6239 11577
rect 7583 11552 7611 11639
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10226 11676 10232 11688
rect 9723 11648 10232 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10318 11636 10324 11688
rect 10376 11636 10382 11688
rect 11698 11676 11704 11688
rect 11659 11648 11704 11676
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 14458 11676 14464 11688
rect 14419 11648 14464 11676
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 14553 11679 14611 11685
rect 14553 11645 14565 11679
rect 14599 11676 14611 11679
rect 15102 11676 15108 11688
rect 14599 11648 15108 11676
rect 14599 11645 14611 11648
rect 14553 11639 14611 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15344 11648 15393 11676
rect 15344 11636 15350 11648
rect 15381 11645 15393 11648
rect 15427 11645 15439 11679
rect 15488 11676 15516 11716
rect 15930 11676 15936 11688
rect 15488 11648 15936 11676
rect 15381 11639 15439 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 9306 11608 9312 11620
rect 7800 11580 9312 11608
rect 7800 11568 7806 11580
rect 9306 11568 9312 11580
rect 9364 11608 9370 11620
rect 10336 11608 10364 11636
rect 10781 11611 10839 11617
rect 10781 11608 10793 11611
rect 9364 11580 10793 11608
rect 9364 11568 9370 11580
rect 10781 11577 10793 11580
rect 10827 11577 10839 11611
rect 10781 11571 10839 11577
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 15626 11611 15684 11617
rect 15626 11608 15638 11611
rect 11020 11580 15638 11608
rect 11020 11568 11026 11580
rect 15626 11577 15638 11580
rect 15672 11608 15684 11611
rect 16666 11608 16672 11620
rect 15672 11580 16672 11608
rect 15672 11577 15684 11580
rect 15626 11571 15684 11577
rect 16666 11568 16672 11580
rect 16724 11568 16730 11620
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 2774 11540 2780 11552
rect 2179 11512 2780 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 2774 11500 2780 11512
rect 2832 11500 2838 11552
rect 3145 11543 3203 11549
rect 3145 11509 3157 11543
rect 3191 11540 3203 11543
rect 3510 11540 3516 11552
rect 3191 11512 3516 11540
rect 3191 11509 3203 11512
rect 3145 11503 3203 11509
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 3605 11543 3663 11549
rect 3605 11509 3617 11543
rect 3651 11540 3663 11543
rect 5074 11540 5080 11552
rect 3651 11512 5080 11540
rect 3651 11509 3663 11512
rect 3605 11503 3663 11509
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5721 11543 5779 11549
rect 5721 11509 5733 11543
rect 5767 11540 5779 11543
rect 5902 11540 5908 11552
rect 5767 11512 5908 11540
rect 5767 11509 5779 11512
rect 5721 11503 5779 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 7285 11543 7343 11549
rect 7285 11540 7297 11543
rect 6696 11512 7297 11540
rect 6696 11500 6702 11512
rect 7285 11509 7297 11512
rect 7331 11540 7343 11543
rect 7558 11540 7564 11552
rect 7331 11512 7564 11540
rect 7331 11509 7343 11512
rect 7285 11503 7343 11509
rect 7558 11500 7564 11512
rect 7616 11540 7622 11552
rect 8938 11540 8944 11552
rect 7616 11512 7709 11540
rect 8899 11512 8944 11540
rect 7616 11500 7622 11512
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10318 11540 10324 11552
rect 10279 11512 10324 11540
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 10652 11512 10701 11540
rect 10652 11500 10658 11512
rect 10689 11509 10701 11512
rect 10735 11540 10747 11543
rect 11054 11540 11060 11552
rect 10735 11512 11060 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11333 11543 11391 11549
rect 11333 11509 11345 11543
rect 11379 11540 11391 11543
rect 11606 11540 11612 11552
rect 11379 11512 11612 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11606 11500 11612 11512
rect 11664 11500 11670 11552
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 13170 11540 13176 11552
rect 11839 11512 13176 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 13449 11543 13507 11549
rect 13449 11540 13461 11543
rect 13320 11512 13461 11540
rect 13320 11500 13326 11512
rect 13449 11509 13461 11512
rect 13495 11509 13507 11543
rect 13449 11503 13507 11509
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 13780 11512 16773 11540
rect 13780 11500 13786 11512
rect 16761 11509 16773 11512
rect 16807 11540 16819 11543
rect 16942 11540 16948 11552
rect 16807 11512 16948 11540
rect 16807 11509 16819 11512
rect 16761 11503 16819 11509
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 2958 11336 2964 11348
rect 1719 11308 2964 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 2958 11296 2964 11308
rect 3016 11296 3022 11348
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 3878 11336 3884 11348
rect 3476 11308 3884 11336
rect 3476 11296 3482 11308
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 7742 11336 7748 11348
rect 5684 11308 7748 11336
rect 5684 11296 5690 11308
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 7834 11296 7840 11348
rect 7892 11336 7898 11348
rect 8573 11339 8631 11345
rect 7892 11308 8432 11336
rect 7892 11296 7898 11308
rect 3694 11268 3700 11280
rect 2056 11240 3700 11268
rect 1486 11200 1492 11212
rect 1447 11172 1492 11200
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 2056 11209 2084 11240
rect 3694 11228 3700 11240
rect 3752 11228 3758 11280
rect 4080 11240 5488 11268
rect 2314 11209 2320 11212
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11169 2099 11203
rect 2308 11200 2320 11209
rect 2227 11172 2320 11200
rect 2041 11163 2099 11169
rect 2308 11163 2320 11172
rect 2372 11200 2378 11212
rect 4080 11200 4108 11240
rect 2372 11172 4108 11200
rect 4332 11203 4390 11209
rect 2314 11160 2320 11163
rect 2372 11160 2378 11172
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 5074 11200 5080 11212
rect 4378 11172 5080 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3844 11104 4077 11132
rect 3844 11092 3850 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 5460 11073 5488 11240
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 7852 11268 7880 11296
rect 7524 11240 7880 11268
rect 7929 11271 7987 11277
rect 7524 11228 7530 11240
rect 7929 11237 7941 11271
rect 7975 11268 7987 11271
rect 8294 11268 8300 11280
rect 7975 11240 8300 11268
rect 7975 11237 7987 11240
rect 7929 11231 7987 11237
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 8404 11268 8432 11308
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 9766 11336 9772 11348
rect 8619 11308 9772 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10505 11339 10563 11345
rect 10505 11305 10517 11339
rect 10551 11336 10563 11339
rect 13354 11336 13360 11348
rect 10551 11308 13360 11336
rect 10551 11305 10563 11308
rect 10505 11299 10563 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 13504 11308 14197 11336
rect 13504 11296 13510 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14458 11336 14464 11348
rect 14419 11308 14464 11336
rect 14185 11299 14243 11305
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 16666 11336 16672 11348
rect 16627 11308 16672 11336
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 16758 11296 16764 11348
rect 16816 11336 16822 11348
rect 16945 11339 17003 11345
rect 16945 11336 16957 11339
rect 16816 11308 16957 11336
rect 16816 11296 16822 11308
rect 16945 11305 16957 11308
rect 16991 11305 17003 11339
rect 16945 11299 17003 11305
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 8404 11240 8953 11268
rect 8941 11237 8953 11240
rect 8987 11268 8999 11271
rect 11146 11268 11152 11280
rect 8987 11240 11152 11268
rect 8987 11237 8999 11240
rect 8941 11231 8999 11237
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 11416 11271 11474 11277
rect 11416 11237 11428 11271
rect 11462 11268 11474 11271
rect 13814 11268 13820 11280
rect 11462 11240 13820 11268
rect 11462 11237 11474 11240
rect 11416 11231 11474 11237
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 17313 11271 17371 11277
rect 17313 11268 17325 11271
rect 16264 11240 17325 11268
rect 16264 11228 16270 11240
rect 17313 11237 17325 11240
rect 17359 11237 17371 11271
rect 17313 11231 17371 11237
rect 6733 11203 6791 11209
rect 6733 11169 6745 11203
rect 6779 11200 6791 11203
rect 8018 11200 8024 11212
rect 6779 11172 7880 11200
rect 7979 11172 8024 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 6825 11135 6883 11141
rect 6825 11132 6837 11135
rect 5776 11104 6837 11132
rect 5776 11092 5782 11104
rect 6825 11101 6837 11104
rect 6871 11101 6883 11135
rect 7006 11132 7012 11144
rect 6967 11104 7012 11132
rect 6825 11095 6883 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 3421 11067 3479 11073
rect 3421 11064 3433 11067
rect 2976 11036 3433 11064
rect 2682 10956 2688 11008
rect 2740 10996 2746 11008
rect 2976 10996 3004 11036
rect 3421 11033 3433 11036
rect 3467 11033 3479 11067
rect 3421 11027 3479 11033
rect 5445 11067 5503 11073
rect 5445 11033 5457 11067
rect 5491 11033 5503 11067
rect 6362 11064 6368 11076
rect 6323 11036 6368 11064
rect 5445 11027 5503 11033
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 7561 11067 7619 11073
rect 7561 11033 7573 11067
rect 7607 11064 7619 11067
rect 7742 11064 7748 11076
rect 7607 11036 7748 11064
rect 7607 11033 7619 11036
rect 7561 11027 7619 11033
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 7852 11064 7880 11172
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 8662 11200 8668 11212
rect 8128 11172 8668 11200
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8128 11132 8156 11172
rect 8662 11160 8668 11172
rect 8720 11200 8726 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8720 11172 9045 11200
rect 8720 11160 8726 11172
rect 9033 11169 9045 11172
rect 9079 11200 9091 11203
rect 10134 11200 10140 11212
rect 9079 11172 10140 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10284 11172 10609 11200
rect 10284 11160 10290 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 13072 11203 13130 11209
rect 13072 11200 13084 11203
rect 10597 11163 10655 11169
rect 12728 11172 13084 11200
rect 7984 11104 8156 11132
rect 8205 11135 8263 11141
rect 7984 11092 7990 11104
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9766 11132 9772 11144
rect 9263 11104 9772 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 8018 11064 8024 11076
rect 7852 11036 8024 11064
rect 8018 11024 8024 11036
rect 8076 11024 8082 11076
rect 8220 11064 8248 11095
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 10962 11132 10968 11144
rect 10827 11104 10968 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 8938 11064 8944 11076
rect 8220 11036 8944 11064
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 10134 11064 10140 11076
rect 10095 11036 10140 11064
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10226 11024 10232 11076
rect 10284 11064 10290 11076
rect 10410 11064 10416 11076
rect 10284 11036 10416 11064
rect 10284 11024 10290 11036
rect 10410 11024 10416 11036
rect 10468 11064 10474 11076
rect 11164 11064 11192 11095
rect 10468 11036 11192 11064
rect 12529 11067 12587 11073
rect 10468 11024 10474 11036
rect 12529 11033 12541 11067
rect 12575 11064 12587 11067
rect 12728 11064 12756 11172
rect 13072 11169 13084 11172
rect 13118 11200 13130 11203
rect 13906 11200 13912 11212
rect 13118 11172 13912 11200
rect 13118 11169 13130 11172
rect 13072 11163 13130 11169
rect 13906 11160 13912 11172
rect 13964 11200 13970 11212
rect 14550 11200 14556 11212
rect 13964 11172 14556 11200
rect 13964 11160 13970 11172
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 15556 11203 15614 11209
rect 15556 11169 15568 11203
rect 15602 11200 15614 11203
rect 15602 11172 16528 11200
rect 15602 11169 15614 11172
rect 15556 11163 15614 11169
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 15286 11132 15292 11144
rect 12860 11104 12905 11132
rect 15247 11104 15292 11132
rect 12860 11092 12866 11104
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 16500 11132 16528 11172
rect 16574 11160 16580 11212
rect 16632 11200 16638 11212
rect 17405 11203 17463 11209
rect 17405 11200 17417 11203
rect 16632 11172 17417 11200
rect 16632 11160 16638 11172
rect 17405 11169 17417 11172
rect 17451 11169 17463 11203
rect 17405 11163 17463 11169
rect 17310 11132 17316 11144
rect 16500 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11132 17647 11135
rect 17770 11132 17776 11144
rect 17635 11104 17776 11132
rect 17635 11101 17647 11104
rect 17589 11095 17647 11101
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 12575 11036 12756 11064
rect 12575 11033 12587 11036
rect 12529 11027 12587 11033
rect 2740 10968 3004 10996
rect 2740 10956 2746 10968
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 8478 10996 8484 11008
rect 3752 10968 8484 10996
rect 3752 10956 3758 10968
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 12342 10996 12348 11008
rect 8720 10968 12348 10996
rect 8720 10956 8726 10968
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 16206 10996 16212 11008
rect 12676 10968 16212 10996
rect 12676 10956 12682 10968
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17770 10996 17776 11008
rect 17000 10968 17776 10996
rect 17000 10956 17006 10968
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 3694 10792 3700 10804
rect 3655 10764 3700 10792
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 4706 10792 4712 10804
rect 4667 10764 4712 10792
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 6822 10792 6828 10804
rect 6564 10764 6828 10792
rect 2866 10724 2872 10736
rect 2332 10696 2872 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 2332 10665 2360 10696
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 6564 10733 6592 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7064 10764 8217 10792
rect 7064 10752 7070 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 6549 10727 6607 10733
rect 6549 10724 6561 10727
rect 5092 10696 6561 10724
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2498 10656 2504 10668
rect 2459 10628 2504 10656
rect 2317 10619 2375 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 4341 10659 4399 10665
rect 3292 10628 4108 10656
rect 3292 10616 3298 10628
rect 4080 10600 4108 10628
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4982 10656 4988 10668
rect 4387 10628 4988 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 1762 10548 1768 10600
rect 1820 10588 1826 10600
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 1820 10560 2237 10588
rect 1820 10548 1826 10560
rect 2225 10557 2237 10560
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10588 2927 10591
rect 3326 10588 3332 10600
rect 2915 10560 3332 10588
rect 2915 10557 2927 10560
rect 2869 10551 2927 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 3602 10588 3608 10600
rect 3563 10560 3608 10588
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 4062 10588 4068 10600
rect 4023 10560 4068 10588
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 4890 10588 4896 10600
rect 4764 10560 4896 10588
rect 4764 10548 4770 10560
rect 4890 10548 4896 10560
rect 4948 10588 4954 10600
rect 5092 10588 5120 10696
rect 6549 10693 6561 10696
rect 6595 10693 6607 10727
rect 6549 10687 6607 10693
rect 5258 10656 5264 10668
rect 5219 10628 5264 10656
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5408 10628 6285 10656
rect 5408 10616 5414 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 6638 10616 6644 10668
rect 6696 10656 6702 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6696 10628 6837 10656
rect 6696 10616 6702 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 8220 10656 8248 10755
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 9861 10795 9919 10801
rect 9861 10792 9873 10795
rect 9824 10764 9873 10792
rect 9824 10752 9830 10764
rect 9861 10761 9873 10764
rect 9907 10792 9919 10795
rect 10778 10792 10784 10804
rect 9907 10764 10784 10792
rect 9907 10761 9919 10764
rect 9861 10755 9919 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11112 10764 11928 10792
rect 11112 10752 11118 10764
rect 11793 10727 11851 10733
rect 11793 10693 11805 10727
rect 11839 10693 11851 10727
rect 11793 10687 11851 10693
rect 8220 10628 8616 10656
rect 6825 10619 6883 10625
rect 4948 10560 5120 10588
rect 5169 10591 5227 10597
rect 4948 10548 4954 10560
rect 5169 10557 5181 10591
rect 5215 10588 5227 10591
rect 7834 10588 7840 10600
rect 5215 10560 7840 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 8018 10548 8024 10600
rect 8076 10588 8082 10600
rect 8294 10588 8300 10600
rect 8076 10560 8300 10588
rect 8076 10548 8082 10560
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10557 8539 10591
rect 8588 10588 8616 10628
rect 8737 10591 8795 10597
rect 8737 10588 8749 10591
rect 8588 10560 8749 10588
rect 8481 10551 8539 10557
rect 8737 10557 8749 10560
rect 8783 10557 8795 10591
rect 8737 10551 8795 10557
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 4203 10492 6684 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 1857 10455 1915 10461
rect 1857 10452 1869 10455
rect 1636 10424 1869 10452
rect 1636 10412 1642 10424
rect 1857 10421 1869 10424
rect 1903 10421 1915 10455
rect 3050 10452 3056 10464
rect 3011 10424 3056 10452
rect 1857 10415 1915 10421
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 3421 10455 3479 10461
rect 3421 10421 3433 10455
rect 3467 10452 3479 10455
rect 3786 10452 3792 10464
rect 3467 10424 3792 10452
rect 3467 10421 3479 10424
rect 3421 10415 3479 10421
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 5074 10452 5080 10464
rect 5035 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 5592 10424 5733 10452
rect 5592 10412 5598 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 6086 10452 6092 10464
rect 6047 10424 6092 10452
rect 5721 10415 5779 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6227 10424 6561 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 6656 10452 6684 10492
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7070 10523 7128 10529
rect 7070 10520 7082 10523
rect 6788 10492 7082 10520
rect 6788 10480 6794 10492
rect 7070 10489 7082 10492
rect 7116 10489 7128 10523
rect 7070 10483 7128 10489
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 8496 10520 8524 10551
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 9824 10560 10149 10588
rect 9824 10548 9830 10560
rect 10137 10557 10149 10560
rect 10183 10588 10195 10591
rect 10226 10588 10232 10600
rect 10183 10560 10232 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10226 10548 10232 10560
rect 10284 10588 10290 10600
rect 11808 10588 11836 10687
rect 11900 10656 11928 10764
rect 12342 10752 12348 10804
rect 12400 10792 12406 10804
rect 16390 10792 16396 10804
rect 12400 10764 16396 10792
rect 12400 10752 12406 10764
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 17310 10752 17316 10804
rect 17368 10792 17374 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17368 10764 17509 10792
rect 17368 10752 17374 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 17497 10755 17555 10761
rect 12526 10684 12532 10736
rect 12584 10724 12590 10736
rect 12584 10696 13032 10724
rect 12584 10684 12590 10696
rect 13004 10656 13032 10696
rect 15749 10659 15807 10665
rect 11900 10628 12940 10656
rect 13004 10628 13400 10656
rect 12912 10597 12940 10628
rect 10284 10560 11836 10588
rect 10284 10548 10290 10560
rect 7616 10492 8524 10520
rect 7616 10480 7622 10492
rect 8938 10480 8944 10532
rect 8996 10520 9002 10532
rect 10382 10523 10440 10529
rect 10382 10520 10394 10523
rect 8996 10492 10394 10520
rect 8996 10480 9002 10492
rect 10382 10489 10394 10492
rect 10428 10489 10440 10523
rect 11808 10520 11836 10560
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10588 12035 10591
rect 12897 10591 12955 10597
rect 12023 10560 12756 10588
rect 12023 10557 12035 10560
rect 11977 10551 12035 10557
rect 12618 10520 12624 10532
rect 11808 10492 12624 10520
rect 10382 10483 10440 10489
rect 12452 10464 12480 10492
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 9214 10452 9220 10464
rect 6656 10424 9220 10452
rect 6549 10415 6607 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 11020 10424 11529 10452
rect 11020 10412 11026 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 12728 10461 12756 10560
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 13262 10588 13268 10600
rect 13223 10560 13268 10588
rect 12897 10551 12955 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13372 10588 13400 10628
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 15795 10628 16252 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 15102 10588 15108 10600
rect 13372 10560 15108 10588
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15470 10588 15476 10600
rect 15344 10560 15476 10588
rect 15344 10548 15350 10560
rect 15470 10548 15476 10560
rect 15528 10588 15534 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15528 10560 16129 10588
rect 15528 10548 15534 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16224 10588 16252 10628
rect 16224 10560 16436 10588
rect 16117 10551 16175 10557
rect 13446 10480 13452 10532
rect 13504 10529 13510 10532
rect 16408 10529 16436 10560
rect 17586 10548 17592 10600
rect 17644 10548 17650 10600
rect 13504 10523 13568 10529
rect 13504 10489 13522 10523
rect 13556 10489 13568 10523
rect 16384 10523 16442 10529
rect 13504 10483 13568 10489
rect 15120 10492 16344 10520
rect 13504 10480 13510 10483
rect 12713 10455 12771 10461
rect 12713 10421 12725 10455
rect 12759 10452 12771 10455
rect 13722 10452 13728 10464
rect 12759 10424 13728 10452
rect 12759 10421 12771 10424
rect 12713 10415 12771 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 14642 10452 14648 10464
rect 14603 10424 14648 10452
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 15120 10461 15148 10492
rect 15105 10455 15163 10461
rect 15105 10421 15117 10455
rect 15151 10421 15163 10455
rect 15105 10415 15163 10421
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 15473 10455 15531 10461
rect 15473 10452 15485 10455
rect 15344 10424 15485 10452
rect 15344 10412 15350 10424
rect 15473 10421 15485 10424
rect 15519 10421 15531 10455
rect 15473 10415 15531 10421
rect 15565 10455 15623 10461
rect 15565 10421 15577 10455
rect 15611 10452 15623 10455
rect 16206 10452 16212 10464
rect 15611 10424 16212 10452
rect 15611 10421 15623 10424
rect 15565 10415 15623 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16316 10452 16344 10492
rect 16384 10489 16396 10523
rect 16430 10520 16442 10523
rect 17604 10520 17632 10548
rect 16430 10492 17632 10520
rect 16430 10489 16442 10492
rect 16384 10483 16442 10489
rect 16776 10464 16804 10492
rect 16574 10452 16580 10464
rect 16316 10424 16580 10452
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 16758 10412 16764 10464
rect 16816 10412 16822 10464
rect 17310 10412 17316 10464
rect 17368 10452 17374 10464
rect 17586 10452 17592 10464
rect 17368 10424 17592 10452
rect 17368 10412 17374 10424
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2556 10220 2789 10248
rect 2556 10208 2562 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 3602 10208 3608 10260
rect 3660 10248 3666 10260
rect 5442 10248 5448 10260
rect 3660 10220 5448 10248
rect 3660 10208 3666 10220
rect 5442 10208 5448 10220
rect 5500 10248 5506 10260
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 5500 10220 7113 10248
rect 5500 10208 5506 10220
rect 7101 10217 7113 10220
rect 7147 10217 7159 10251
rect 7101 10211 7159 10217
rect 7561 10251 7619 10257
rect 7561 10217 7573 10251
rect 7607 10248 7619 10251
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 7607 10220 9045 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 9033 10217 9045 10220
rect 9079 10217 9091 10251
rect 9033 10211 9091 10217
rect 11057 10251 11115 10257
rect 11057 10217 11069 10251
rect 11103 10248 11115 10251
rect 11238 10248 11244 10260
rect 11103 10220 11244 10248
rect 11103 10217 11115 10220
rect 11057 10211 11115 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 11977 10251 12035 10257
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12989 10251 13047 10257
rect 12023 10220 12940 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 1664 10183 1722 10189
rect 1664 10149 1676 10183
rect 1710 10180 1722 10183
rect 2682 10180 2688 10192
rect 1710 10152 2688 10180
rect 1710 10149 1722 10152
rect 1664 10143 1722 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 6638 10180 6644 10192
rect 4847 10152 6644 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 7466 10180 7472 10192
rect 7064 10152 7472 10180
rect 7064 10140 7070 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 7929 10183 7987 10189
rect 7929 10149 7941 10183
rect 7975 10180 7987 10183
rect 9490 10180 9496 10192
rect 7975 10152 9496 10180
rect 7975 10149 7987 10152
rect 7929 10143 7987 10149
rect 9490 10140 9496 10152
rect 9548 10140 9554 10192
rect 12345 10183 12403 10189
rect 12345 10149 12357 10183
rect 12391 10180 12403 10183
rect 12526 10180 12532 10192
rect 12391 10152 12532 10180
rect 12391 10149 12403 10152
rect 12345 10143 12403 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 12912 10180 12940 10220
rect 12989 10217 13001 10251
rect 13035 10248 13047 10251
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 13035 10220 14381 10248
rect 13035 10217 13047 10220
rect 12989 10211 13047 10217
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 14369 10211 14427 10217
rect 17034 10208 17040 10260
rect 17092 10248 17098 10260
rect 17129 10251 17187 10257
rect 17129 10248 17141 10251
rect 17092 10220 17141 10248
rect 17092 10208 17098 10220
rect 17129 10217 17141 10220
rect 17175 10217 17187 10251
rect 17129 10211 17187 10217
rect 13449 10183 13507 10189
rect 13449 10180 13461 10183
rect 12912 10152 13461 10180
rect 13449 10149 13461 10152
rect 13495 10149 13507 10183
rect 13630 10180 13636 10192
rect 13449 10143 13507 10149
rect 13556 10152 13636 10180
rect 3053 10115 3111 10121
rect 3053 10081 3065 10115
rect 3099 10081 3111 10115
rect 3053 10075 3111 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 3068 9976 3096 10075
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 3844 10084 5457 10112
rect 3844 10072 3850 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 5712 10115 5770 10121
rect 5712 10081 5724 10115
rect 5758 10112 5770 10115
rect 7190 10112 7196 10124
rect 5758 10084 7196 10112
rect 5758 10081 5770 10084
rect 5712 10075 5770 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10112 7343 10115
rect 7650 10112 7656 10124
rect 7331 10084 7656 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8202 10112 8208 10124
rect 8067 10084 8208 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8938 10112 8944 10124
rect 8899 10084 8944 10112
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9398 10112 9404 10124
rect 9088 10084 9404 10112
rect 9088 10072 9094 10084
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 9766 10112 9772 10124
rect 9723 10084 9772 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 9944 10115 10002 10121
rect 9944 10081 9956 10115
rect 9990 10112 10002 10115
rect 10962 10112 10968 10124
rect 9990 10084 10968 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 13354 10112 13360 10124
rect 13315 10084 13360 10112
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 4890 10044 4896 10056
rect 4851 10016 4896 10044
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5350 10044 5356 10056
rect 5123 10016 5356 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 7208 10044 7236 10072
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 7208 10016 8125 10044
rect 8113 10013 8125 10016
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 5442 9976 5448 9988
rect 3068 9948 5448 9976
rect 5442 9936 5448 9948
rect 5500 9936 5506 9988
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 6825 9979 6883 9985
rect 6825 9976 6837 9979
rect 6788 9948 6837 9976
rect 6788 9936 6794 9948
rect 6825 9945 6837 9948
rect 6871 9976 6883 9979
rect 9140 9976 9168 10007
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12032 10016 12449 10044
rect 12032 10004 12038 10016
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10044 12679 10047
rect 12710 10044 12716 10056
rect 12667 10016 12716 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 13556 10053 13584 10152
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 16390 10140 16396 10192
rect 16448 10180 16454 10192
rect 17497 10183 17555 10189
rect 17497 10180 17509 10183
rect 16448 10152 17509 10180
rect 16448 10140 16454 10152
rect 17497 10149 17509 10152
rect 17543 10149 17555 10183
rect 17497 10143 17555 10149
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 13780 10084 15669 10112
rect 13780 10072 13786 10084
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 15657 10075 15715 10081
rect 16485 10115 16543 10121
rect 16485 10081 16497 10115
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 17310 10112 17316 10124
rect 16623 10084 17316 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 13688 10016 14473 10044
rect 13688 10004 13694 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14550 10004 14556 10056
rect 14608 10044 14614 10056
rect 14608 10016 14653 10044
rect 14608 10004 14614 10016
rect 6871 9948 9168 9976
rect 6871 9945 6883 9948
rect 6825 9939 6883 9945
rect 13170 9936 13176 9988
rect 13228 9976 13234 9988
rect 14001 9979 14059 9985
rect 14001 9976 14013 9979
rect 13228 9948 14013 9976
rect 13228 9936 13234 9948
rect 14001 9945 14013 9948
rect 14047 9945 14059 9979
rect 14001 9939 14059 9945
rect 14090 9936 14096 9988
rect 14148 9976 14154 9988
rect 16500 9976 16528 10075
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 16758 10044 16764 10056
rect 16671 10016 16764 10044
rect 16758 10004 16764 10016
rect 16816 10044 16822 10056
rect 17034 10044 17040 10056
rect 16816 10016 17040 10044
rect 16816 10004 16822 10016
rect 17034 10004 17040 10016
rect 17092 10004 17098 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17770 10044 17776 10056
rect 17731 10016 17776 10044
rect 17589 10007 17647 10013
rect 14148 9948 16528 9976
rect 14148 9936 14154 9948
rect 16942 9936 16948 9988
rect 17000 9976 17006 9988
rect 17604 9976 17632 10007
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 18138 10044 18144 10056
rect 18099 10016 18144 10044
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 17000 9948 17632 9976
rect 17000 9936 17006 9948
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 4430 9908 4436 9920
rect 4391 9880 4436 9908
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4982 9868 4988 9920
rect 5040 9908 5046 9920
rect 7466 9908 7472 9920
rect 5040 9880 7472 9908
rect 5040 9868 5046 9880
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8352 9880 8585 9908
rect 8352 9868 8358 9880
rect 8573 9877 8585 9880
rect 8619 9877 8631 9911
rect 8573 9871 8631 9877
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 12342 9908 12348 9920
rect 8720 9880 12348 9908
rect 8720 9868 8726 9880
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 13722 9908 13728 9920
rect 13320 9880 13728 9908
rect 13320 9868 13326 9880
rect 13722 9868 13728 9880
rect 13780 9908 13786 9920
rect 15470 9908 15476 9920
rect 13780 9880 15476 9908
rect 13780 9868 13786 9880
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16758 9908 16764 9920
rect 16163 9880 16764 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 3786 9704 3792 9716
rect 1452 9676 3792 9704
rect 1452 9664 1458 9676
rect 2332 9577 2360 9676
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4709 9707 4767 9713
rect 4709 9673 4721 9707
rect 4755 9704 4767 9707
rect 5074 9704 5080 9716
rect 4755 9676 5080 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 6641 9707 6699 9713
rect 6641 9673 6653 9707
rect 6687 9704 6699 9707
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6687 9676 6837 9704
rect 6687 9673 6699 9676
rect 6641 9667 6699 9673
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8662 9704 8668 9716
rect 7616 9676 8668 9704
rect 7616 9664 7622 9676
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 11238 9704 11244 9716
rect 9272 9676 9720 9704
rect 9272 9664 9278 9676
rect 3510 9596 3516 9648
rect 3568 9636 3574 9648
rect 5166 9636 5172 9648
rect 3568 9608 5172 9636
rect 3568 9596 3574 9608
rect 5166 9596 5172 9608
rect 5224 9636 5230 9648
rect 5718 9636 5724 9648
rect 5224 9608 5308 9636
rect 5679 9608 5724 9636
rect 5224 9596 5230 9608
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 6178 9596 6184 9648
rect 6236 9636 6242 9648
rect 7745 9639 7803 9645
rect 7745 9636 7757 9639
rect 6236 9608 7757 9636
rect 6236 9596 6242 9608
rect 7745 9605 7757 9608
rect 7791 9605 7803 9639
rect 7745 9599 7803 9605
rect 7837 9639 7895 9645
rect 7837 9605 7849 9639
rect 7883 9636 7895 9639
rect 8938 9636 8944 9648
rect 7883 9608 8944 9636
rect 7883 9605 7895 9608
rect 7837 9599 7895 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 9493 9639 9551 9645
rect 9493 9605 9505 9639
rect 9539 9636 9551 9639
rect 9582 9636 9588 9648
rect 9539 9608 9588 9636
rect 9539 9605 9551 9608
rect 9493 9599 9551 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 9692 9636 9720 9676
rect 11164 9676 11244 9704
rect 10321 9639 10379 9645
rect 10321 9636 10333 9639
rect 9692 9608 10333 9636
rect 10321 9605 10333 9608
rect 10367 9605 10379 9639
rect 10321 9599 10379 9605
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 4338 9568 4344 9580
rect 2317 9531 2375 9537
rect 3896 9540 4344 9568
rect 1670 9500 1676 9512
rect 1631 9472 1676 9500
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 3896 9500 3924 9540
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4798 9568 4804 9580
rect 4540 9540 4804 9568
rect 4540 9512 4568 9540
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 5175 9512 5203 9596
rect 11164 9580 11192 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 11333 9707 11391 9713
rect 11333 9673 11345 9707
rect 11379 9704 11391 9707
rect 13630 9704 13636 9716
rect 11379 9676 13636 9704
rect 11379 9673 11391 9676
rect 11333 9667 11391 9673
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 14274 9704 14280 9716
rect 14056 9676 14280 9704
rect 14056 9664 14062 9676
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 16206 9704 16212 9716
rect 14516 9676 16212 9704
rect 14516 9664 14522 9676
rect 15856 9648 15884 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 16942 9664 16948 9716
rect 17000 9704 17006 9716
rect 17954 9704 17960 9716
rect 17000 9676 17960 9704
rect 17000 9664 17006 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 13538 9636 13544 9648
rect 13451 9608 13544 9636
rect 5350 9568 5356 9580
rect 5311 9540 5356 9568
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 6730 9568 6736 9580
rect 6411 9540 6736 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7248 9540 7389 9568
rect 7248 9528 7254 9540
rect 7377 9537 7389 9540
rect 7423 9568 7435 9571
rect 8202 9568 8208 9580
rect 7423 9540 8208 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 8202 9528 8208 9540
rect 8260 9568 8266 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8260 9540 8401 9568
rect 8260 9528 8266 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 8536 9540 9965 9568
rect 8536 9528 8542 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 10962 9568 10968 9580
rect 10183 9540 10968 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11146 9528 11152 9580
rect 11204 9528 11210 9580
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12023 9540 12296 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 2424 9472 3924 9500
rect 3973 9503 4031 9509
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 2424 9432 2452 9472
rect 3973 9469 3985 9503
rect 4019 9500 4031 9503
rect 4522 9500 4528 9512
rect 4019 9472 4528 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 4522 9460 4528 9472
rect 4580 9460 4586 9512
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 5077 9503 5135 9509
rect 5077 9500 5089 9503
rect 4672 9472 5089 9500
rect 4672 9460 4678 9472
rect 5077 9469 5089 9472
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 5166 9460 5172 9512
rect 5224 9460 5230 9512
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8297 9503 8355 9509
rect 8297 9500 8309 9503
rect 8168 9472 8309 9500
rect 8168 9460 8174 9472
rect 8297 9469 8309 9472
rect 8343 9469 8355 9503
rect 8297 9463 8355 9469
rect 8570 9460 8576 9512
rect 8628 9500 8634 9512
rect 9214 9500 9220 9512
rect 8628 9472 9220 9500
rect 8628 9460 8634 9472
rect 9214 9460 9220 9472
rect 9272 9500 9278 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 9272 9472 10793 9500
rect 9272 9460 9278 9472
rect 10781 9469 10793 9472
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 2004 9404 2452 9432
rect 2004 9392 2010 9404
rect 2498 9392 2504 9444
rect 2556 9441 2562 9444
rect 2556 9435 2620 9441
rect 2556 9401 2574 9435
rect 2608 9401 2620 9435
rect 2556 9395 2620 9401
rect 2556 9392 2562 9395
rect 2682 9392 2688 9444
rect 2740 9432 2746 9444
rect 5718 9432 5724 9444
rect 2740 9404 5724 9432
rect 2740 9392 2746 9404
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 6641 9435 6699 9441
rect 6641 9432 6653 9435
rect 6135 9404 6653 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 6641 9401 6653 9404
rect 6687 9401 6699 9435
rect 6641 9395 6699 9401
rect 7193 9435 7251 9441
rect 7193 9401 7205 9435
rect 7239 9432 7251 9435
rect 7558 9432 7564 9444
rect 7239 9404 7564 9432
rect 7239 9401 7251 9404
rect 7193 9395 7251 9401
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 8849 9435 8907 9441
rect 8849 9432 8861 9435
rect 8251 9404 8861 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 8849 9401 8861 9404
rect 8895 9401 8907 9435
rect 8849 9395 8907 9401
rect 9306 9392 9312 9444
rect 9364 9432 9370 9444
rect 9766 9432 9772 9444
rect 9364 9404 9772 9432
rect 9364 9392 9370 9404
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 12268 9432 12296 9540
rect 12360 9540 12449 9568
rect 12360 9512 12388 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12342 9460 12348 9512
rect 12400 9460 12406 9512
rect 13464 9500 13492 9608
rect 13538 9596 13544 9608
rect 13596 9636 13602 9648
rect 13814 9636 13820 9648
rect 13596 9608 13820 9636
rect 13596 9596 13602 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 15838 9596 15844 9648
rect 15896 9596 15902 9648
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 17770 9636 17776 9648
rect 17460 9608 17776 9636
rect 17460 9596 17466 9608
rect 17770 9596 17776 9608
rect 17828 9596 17834 9648
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 16022 9568 16028 9580
rect 15528 9540 16028 9568
rect 15528 9528 15534 9540
rect 16022 9528 16028 9540
rect 16080 9568 16086 9580
rect 16301 9571 16359 9577
rect 16301 9568 16313 9571
rect 16080 9540 16313 9568
rect 16080 9528 16086 9540
rect 16301 9537 16313 9540
rect 16347 9537 16359 9571
rect 16301 9531 16359 9537
rect 12544 9472 13492 9500
rect 12544 9432 12572 9472
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 13872 9472 14105 9500
rect 13872 9460 13878 9472
rect 14093 9469 14105 9472
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14360 9503 14418 9509
rect 14360 9469 14372 9503
rect 14406 9500 14418 9503
rect 14642 9500 14648 9512
rect 14406 9472 14648 9500
rect 14406 9469 14418 9472
rect 14360 9463 14418 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 15102 9460 15108 9512
rect 15160 9500 15166 9512
rect 15378 9500 15384 9512
rect 15160 9472 15384 9500
rect 15160 9460 15166 9472
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 12710 9441 12716 9444
rect 12704 9432 12716 9441
rect 12268 9404 12572 9432
rect 12671 9404 12716 9432
rect 12704 9395 12716 9404
rect 12710 9392 12716 9395
rect 12768 9392 12774 9444
rect 16568 9435 16626 9441
rect 16568 9401 16580 9435
rect 16614 9432 16626 9435
rect 17402 9432 17408 9444
rect 16614 9404 17408 9432
rect 16614 9401 16626 9404
rect 16568 9395 16626 9401
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 1857 9367 1915 9373
rect 1857 9333 1869 9367
rect 1903 9364 1915 9367
rect 3510 9364 3516 9376
rect 1903 9336 3516 9364
rect 1903 9333 1915 9336
rect 1857 9327 1915 9333
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3697 9367 3755 9373
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 4062 9364 4068 9376
rect 3743 9336 4068 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4338 9364 4344 9376
rect 4203 9336 4344 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 4856 9336 5181 9364
rect 4856 9324 4862 9336
rect 5169 9333 5181 9336
rect 5215 9364 5227 9367
rect 5626 9364 5632 9376
rect 5215 9336 5632 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 6730 9364 6736 9376
rect 6512 9336 6736 9364
rect 6512 9324 6518 9336
rect 6730 9324 6736 9336
rect 6788 9364 6794 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6788 9336 7297 9364
rect 6788 9324 6794 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 7745 9367 7803 9373
rect 7745 9333 7757 9367
rect 7791 9364 7803 9367
rect 9858 9364 9864 9376
rect 7791 9336 9864 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 10376 9336 10701 9364
rect 10376 9324 10382 9336
rect 10689 9333 10701 9336
rect 10735 9333 10747 9367
rect 11698 9364 11704 9376
rect 11659 9336 11704 9364
rect 10689 9327 10747 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 11793 9367 11851 9373
rect 11793 9333 11805 9367
rect 11839 9364 11851 9367
rect 12526 9364 12532 9376
rect 11839 9336 12532 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 14458 9364 14464 9376
rect 12676 9336 14464 9364
rect 12676 9324 12682 9336
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 15473 9367 15531 9373
rect 15473 9364 15485 9367
rect 14700 9336 15485 9364
rect 14700 9324 14706 9336
rect 15473 9333 15485 9336
rect 15519 9333 15531 9367
rect 15473 9327 15531 9333
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 17092 9336 17693 9364
rect 17092 9324 17098 9336
rect 17681 9333 17693 9336
rect 17727 9364 17739 9367
rect 17954 9364 17960 9376
rect 17727 9336 17960 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 4430 9160 4436 9172
rect 2363 9132 4436 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7282 9160 7288 9172
rect 7147 9132 7288 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8260 9132 8769 9160
rect 8260 9120 8266 9132
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 8757 9123 8815 9129
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10502 9160 10508 9172
rect 10183 9132 10508 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11756 9132 12081 9160
rect 11756 9120 11762 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12434 9160 12440 9172
rect 12395 9132 12440 9160
rect 12069 9123 12127 9129
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12584 9132 13093 9160
rect 12584 9120 12590 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 13320 9132 13461 9160
rect 13320 9120 13326 9132
rect 13449 9129 13461 9132
rect 13495 9129 13507 9163
rect 13449 9123 13507 9129
rect 13541 9163 13599 9169
rect 13541 9129 13553 9163
rect 13587 9160 13599 9163
rect 13998 9160 14004 9172
rect 13587 9132 14004 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 15105 9163 15163 9169
rect 15105 9129 15117 9163
rect 15151 9160 15163 9163
rect 16482 9160 16488 9172
rect 15151 9132 16488 9160
rect 15151 9129 15163 9132
rect 15105 9123 15163 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 2455 9064 3832 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1443 8996 3280 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 2774 8888 2780 8900
rect 1627 8860 2780 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 3252 8888 3280 8996
rect 3326 8984 3332 9036
rect 3384 9024 3390 9036
rect 3804 9024 3832 9064
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 4246 9092 4252 9104
rect 4120 9064 4252 9092
rect 4120 9052 4126 9064
rect 4246 9052 4252 9064
rect 4304 9101 4310 9104
rect 4304 9095 4368 9101
rect 4304 9061 4322 9095
rect 4356 9061 4368 9095
rect 4304 9055 4368 9061
rect 5988 9095 6046 9101
rect 5988 9061 6000 9095
rect 6034 9092 6046 9095
rect 6270 9092 6276 9104
rect 6034 9064 6276 9092
rect 6034 9061 6046 9064
rect 5988 9055 6046 9061
rect 4304 9052 4310 9055
rect 6270 9052 6276 9064
rect 6328 9052 6334 9104
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 7300 9092 7328 9120
rect 7622 9095 7680 9101
rect 7622 9092 7634 9095
rect 6788 9064 6868 9092
rect 7300 9064 7634 9092
rect 6788 9052 6794 9064
rect 5534 9024 5540 9036
rect 3384 8996 3429 9024
rect 3804 8996 5540 9024
rect 3384 8984 3390 8996
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 6546 9024 6552 9036
rect 5767 8996 6552 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 6546 8984 6552 8996
rect 6604 9024 6610 9036
rect 6840 9024 6868 9064
rect 7622 9061 7634 9064
rect 7668 9061 7680 9095
rect 7622 9055 7680 9061
rect 10597 9095 10655 9101
rect 10597 9061 10609 9095
rect 10643 9092 10655 9095
rect 11885 9095 11943 9101
rect 10643 9064 11836 9092
rect 10643 9061 10655 9064
rect 10597 9055 10655 9061
rect 10410 9024 10416 9036
rect 6604 8996 6776 9024
rect 6840 8996 10416 9024
rect 6604 8984 6610 8996
rect 6748 8968 6776 8996
rect 10410 8984 10416 8996
rect 10468 9024 10474 9036
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 10468 8996 10517 9024
rect 10468 8984 10474 8996
rect 10505 8993 10517 8996
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3326 8888 3332 8900
rect 3252 8860 3332 8888
rect 3326 8848 3332 8860
rect 3384 8848 3390 8900
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2464 8792 2973 8820
rect 2464 8780 2470 8792
rect 2961 8789 2973 8792
rect 3007 8789 3019 8823
rect 3620 8820 3648 8919
rect 3786 8916 3792 8968
rect 3844 8956 3850 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3844 8928 4077 8956
rect 3844 8916 3850 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 6788 8928 7389 8956
rect 6788 8916 6794 8928
rect 7377 8925 7389 8928
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 4706 8820 4712 8832
rect 3620 8792 4712 8820
rect 2961 8783 3019 8789
rect 4706 8780 4712 8792
rect 4764 8820 4770 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 4764 8792 5457 8820
rect 4764 8780 4770 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 5445 8783 5503 8789
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 7098 8820 7104 8832
rect 5776 8792 7104 8820
rect 5776 8780 5782 8792
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 8018 8820 8024 8832
rect 7616 8792 8024 8820
rect 7616 8780 7622 8792
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 10612 8820 10640 9055
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 11808 9024 11836 9064
rect 11885 9061 11897 9095
rect 11931 9092 11943 9095
rect 15381 9095 15439 9101
rect 11931 9064 15240 9092
rect 11931 9061 11943 9064
rect 11885 9055 11943 9061
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 11471 8996 11652 9024
rect 11808 8996 12541 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10962 8956 10968 8968
rect 10827 8928 10968 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 8168 8792 10640 8820
rect 8168 8780 8174 8792
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 11020 8792 11069 8820
rect 11020 8780 11026 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11532 8820 11560 8919
rect 11624 8888 11652 8996
rect 12529 8993 12541 8996
rect 12575 9024 12587 9027
rect 14090 9024 14096 9036
rect 12575 8996 14096 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 14550 9024 14556 9036
rect 14463 8996 14556 9024
rect 14550 8984 14556 8996
rect 14608 9024 14614 9036
rect 15105 9027 15163 9033
rect 15105 9024 15117 9027
rect 14608 8996 15117 9024
rect 14608 8984 14614 8996
rect 15105 8993 15117 8996
rect 15151 8993 15163 9027
rect 15212 9024 15240 9064
rect 15381 9061 15393 9095
rect 15427 9092 15439 9095
rect 16666 9092 16672 9104
rect 15427 9064 16672 9092
rect 15427 9061 15439 9064
rect 15381 9055 15439 9061
rect 16666 9052 16672 9064
rect 16724 9052 16730 9104
rect 16298 9033 16304 9036
rect 16281 9027 16304 9033
rect 16281 9024 16293 9027
rect 15212 8996 16293 9024
rect 15105 8987 15163 8993
rect 16281 8993 16293 8996
rect 16356 9024 16362 9036
rect 16356 8996 16429 9024
rect 16281 8987 16304 8993
rect 16298 8984 16304 8987
rect 16356 8984 16362 8996
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 17865 9027 17923 9033
rect 17865 9024 17877 9027
rect 17828 8996 17877 9024
rect 17828 8984 17834 8996
rect 17865 8993 17877 8996
rect 17911 8993 17923 9027
rect 17865 8987 17923 8993
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11747 8928 11897 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 12710 8956 12716 8968
rect 12671 8928 12716 8956
rect 11885 8919 11943 8925
rect 12710 8916 12716 8928
rect 12768 8956 12774 8968
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 12768 8928 13645 8956
rect 12768 8916 12774 8928
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 14516 8928 14657 8956
rect 14516 8916 14522 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14645 8919 14703 8925
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 16022 8956 16028 8968
rect 14792 8928 14837 8956
rect 15983 8928 16028 8956
rect 14792 8916 14798 8928
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 12986 8888 12992 8900
rect 11624 8860 12992 8888
rect 12986 8848 12992 8860
rect 13044 8848 13050 8900
rect 14108 8860 16068 8888
rect 14108 8820 14136 8860
rect 11532 8792 14136 8820
rect 14185 8823 14243 8829
rect 11057 8783 11115 8789
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 14550 8820 14556 8832
rect 14231 8792 14556 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 15102 8820 15108 8832
rect 15063 8792 15108 8820
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16040 8820 16068 8860
rect 16206 8820 16212 8832
rect 16040 8792 16212 8820
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 17402 8820 17408 8832
rect 17315 8792 17408 8820
rect 17402 8780 17408 8792
rect 17460 8820 17466 8832
rect 17862 8820 17868 8832
rect 17460 8792 17868 8820
rect 17460 8780 17466 8792
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3476 8588 3525 8616
rect 3476 8576 3482 8588
rect 3513 8585 3525 8588
rect 3559 8585 3571 8619
rect 3513 8579 3571 8585
rect 3786 8576 3792 8628
rect 3844 8616 3850 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 3844 8588 4353 8616
rect 3844 8576 3850 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 5258 8616 5264 8628
rect 4341 8579 4399 8585
rect 4908 8588 5264 8616
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 4908 8548 4936 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6236 8588 6837 8616
rect 6236 8576 6242 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 7708 8588 8493 8616
rect 7708 8576 7714 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 11054 8616 11060 8628
rect 11015 8588 11060 8616
rect 8481 8579 8539 8585
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8616 11391 8619
rect 14093 8619 14151 8625
rect 11379 8588 13308 8616
rect 11379 8585 11391 8588
rect 11333 8579 11391 8585
rect 2648 8520 4936 8548
rect 2648 8508 2654 8520
rect 6270 8508 6276 8560
rect 6328 8548 6334 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 6328 8520 6377 8548
rect 6328 8508 6334 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 7837 8551 7895 8557
rect 7837 8548 7849 8551
rect 6365 8511 6423 8517
rect 6472 8520 7849 8548
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 3418 8480 3424 8492
rect 2924 8452 3424 8480
rect 2924 8440 2930 8452
rect 3418 8440 3424 8452
rect 3476 8440 3482 8492
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3660 8452 3985 8480
rect 3660 8440 3666 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4246 8480 4252 8492
rect 4203 8452 4252 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4387 8452 4997 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 1664 8415 1722 8421
rect 1664 8381 1676 8415
rect 1710 8412 1722 8415
rect 4614 8412 4620 8424
rect 1710 8384 4620 8412
rect 1710 8381 1722 8384
rect 1664 8375 1722 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 6472 8412 6500 8520
rect 7837 8517 7849 8520
rect 7883 8517 7895 8551
rect 11072 8548 11100 8576
rect 11514 8548 11520 8560
rect 11072 8520 11520 8548
rect 7837 8511 7895 8517
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 11624 8520 12449 8548
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 8202 8480 8208 8492
rect 7515 8452 8208 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 11624 8480 11652 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 13280 8548 13308 8588
rect 14093 8585 14105 8619
rect 14139 8616 14151 8619
rect 14139 8588 17264 8616
rect 14139 8585 14151 8588
rect 14093 8579 14151 8585
rect 14182 8548 14188 8560
rect 13280 8520 14188 8548
rect 12437 8511 12495 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 16206 8508 16212 8560
rect 16264 8548 16270 8560
rect 16761 8551 16819 8557
rect 16761 8548 16773 8551
rect 16264 8520 16773 8548
rect 16264 8508 16270 8520
rect 16761 8517 16773 8520
rect 16807 8517 16819 8551
rect 16761 8511 16819 8517
rect 11348 8452 11652 8480
rect 5092 8384 6500 8412
rect 2498 8304 2504 8356
rect 2556 8344 2562 8356
rect 3881 8347 3939 8353
rect 3881 8344 3893 8347
rect 2556 8316 3893 8344
rect 2556 8304 2562 8316
rect 3881 8313 3893 8316
rect 3927 8313 3939 8347
rect 5092 8344 5120 8384
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 7653 8415 7711 8421
rect 6696 8384 7512 8412
rect 6696 8372 6702 8384
rect 5258 8353 5264 8356
rect 5252 8344 5264 8353
rect 3881 8307 3939 8313
rect 4172 8316 5120 8344
rect 5219 8316 5264 8344
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 2866 8276 2872 8288
rect 2823 8248 2872 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4172 8276 4200 8316
rect 5252 8307 5264 8316
rect 5258 8304 5264 8307
rect 5316 8304 5322 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7193 8347 7251 8353
rect 7193 8344 7205 8347
rect 6972 8316 7205 8344
rect 6972 8304 6978 8316
rect 7193 8313 7205 8316
rect 7239 8313 7251 8347
rect 7193 8307 7251 8313
rect 7285 8347 7343 8353
rect 7285 8313 7297 8347
rect 7331 8344 7343 8347
rect 7374 8344 7380 8356
rect 7331 8316 7380 8344
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 7484 8344 7512 8384
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 7834 8412 7840 8424
rect 7699 8384 7840 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 8711 8384 10517 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 10505 8381 10517 8384
rect 10551 8412 10563 8415
rect 11241 8415 11299 8421
rect 11241 8412 11253 8415
rect 10551 8384 11253 8412
rect 10551 8381 10563 8384
rect 10505 8375 10563 8381
rect 11241 8381 11253 8384
rect 11287 8381 11299 8415
rect 11241 8375 11299 8381
rect 8021 8347 8079 8353
rect 8021 8344 8033 8347
rect 7484 8316 8033 8344
rect 8021 8313 8033 8316
rect 8067 8313 8079 8347
rect 8021 8307 8079 8313
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 8168 8316 8953 8344
rect 8168 8304 8174 8316
rect 8941 8313 8953 8316
rect 8987 8313 8999 8347
rect 11348 8344 11376 8452
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 11940 8452 11985 8480
rect 11940 8440 11946 8452
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12584 8452 13001 8480
rect 12584 8440 12590 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 14550 8480 14556 8492
rect 14511 8452 14556 8480
rect 12989 8443 13047 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 17236 8489 17264 8588
rect 18230 8548 18236 8560
rect 18191 8520 18236 8548
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 17221 8483 17279 8489
rect 14700 8452 14745 8480
rect 14700 8440 14706 8452
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 15010 8412 15016 8424
rect 12360 8384 15016 8412
rect 11701 8347 11759 8353
rect 11701 8344 11713 8347
rect 11348 8316 11713 8344
rect 8941 8307 8999 8313
rect 11701 8313 11713 8316
rect 11747 8313 11759 8347
rect 11701 8307 11759 8313
rect 11793 8347 11851 8353
rect 11793 8313 11805 8347
rect 11839 8344 11851 8347
rect 12066 8344 12072 8356
rect 11839 8316 12072 8344
rect 11839 8313 11851 8316
rect 11793 8307 11851 8313
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 4522 8276 4528 8288
rect 4120 8248 4200 8276
rect 4483 8248 4528 8276
rect 4120 8236 4126 8248
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 8386 8276 8392 8288
rect 7524 8248 8392 8276
rect 7524 8236 7530 8248
rect 8386 8236 8392 8248
rect 8444 8276 8450 8288
rect 11146 8276 11152 8288
rect 8444 8248 11152 8276
rect 8444 8236 8450 8248
rect 11146 8236 11152 8248
rect 11204 8276 11210 8288
rect 12360 8276 12388 8384
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 15105 8415 15163 8421
rect 15105 8381 15117 8415
rect 15151 8381 15163 8415
rect 15105 8375 15163 8381
rect 12434 8304 12440 8356
rect 12492 8344 12498 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12492 8316 12909 8344
rect 12492 8304 12498 8316
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 13722 8344 13728 8356
rect 13635 8316 13728 8344
rect 12897 8307 12955 8313
rect 13722 8304 13728 8316
rect 13780 8344 13786 8356
rect 15120 8344 15148 8375
rect 15194 8372 15200 8424
rect 15252 8412 15258 8424
rect 15372 8415 15430 8421
rect 15372 8412 15384 8415
rect 15252 8384 15384 8412
rect 15252 8372 15258 8384
rect 15372 8381 15384 8384
rect 15418 8412 15430 8415
rect 16482 8412 16488 8424
rect 15418 8384 16488 8412
rect 15418 8381 15430 8384
rect 15372 8375 15430 8381
rect 16482 8372 16488 8384
rect 16540 8412 16546 8424
rect 17328 8412 17356 8443
rect 16540 8384 17356 8412
rect 18049 8415 18107 8421
rect 16540 8372 16546 8384
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 13780 8316 15148 8344
rect 13780 8304 13786 8316
rect 16298 8304 16304 8356
rect 16356 8344 16362 8356
rect 16356 8316 16528 8344
rect 16356 8304 16362 8316
rect 11204 8248 12388 8276
rect 12805 8279 12863 8285
rect 11204 8236 11210 8248
rect 12805 8245 12817 8279
rect 12851 8276 12863 8279
rect 13446 8276 13452 8288
rect 12851 8248 13452 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 13740 8276 13768 8304
rect 13596 8248 13768 8276
rect 14461 8279 14519 8285
rect 13596 8236 13602 8248
rect 14461 8245 14473 8279
rect 14507 8276 14519 8279
rect 14734 8276 14740 8288
rect 14507 8248 14740 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 15286 8276 15292 8288
rect 14884 8248 15292 8276
rect 14884 8236 14890 8248
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 16500 8285 16528 8316
rect 17034 8304 17040 8356
rect 17092 8344 17098 8356
rect 18064 8344 18092 8375
rect 17092 8316 18092 8344
rect 17092 8304 17098 8316
rect 16485 8279 16543 8285
rect 16485 8245 16497 8279
rect 16531 8245 16543 8279
rect 17126 8276 17132 8288
rect 17087 8248 17132 8276
rect 16485 8239 16543 8245
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2317 8075 2375 8081
rect 2317 8041 2329 8075
rect 2363 8072 2375 8075
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2363 8044 2973 8072
rect 2363 8041 2375 8044
rect 2317 8035 2375 8041
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 3200 8044 3341 8072
rect 3200 8032 3206 8044
rect 3329 8041 3341 8044
rect 3375 8072 3387 8075
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3375 8044 3801 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 4111 8044 5549 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 6595 8044 7297 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 10226 8072 10232 8084
rect 7791 8044 10232 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10870 8072 10876 8084
rect 10831 8044 10876 8072
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11790 8072 11796 8084
rect 11072 8044 11796 8072
rect 2406 8004 2412 8016
rect 2367 7976 2412 8004
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 3421 8007 3479 8013
rect 3421 7973 3433 8007
rect 3467 8004 3479 8007
rect 3602 8004 3608 8016
rect 3467 7976 3608 8004
rect 3467 7973 3479 7976
rect 3421 7967 3479 7973
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 4893 8007 4951 8013
rect 4893 8004 4905 8007
rect 4724 7976 4905 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1486 7936 1492 7948
rect 1443 7908 1492 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 4430 7936 4436 7948
rect 4391 7908 4436 7936
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 4724 7936 4752 7976
rect 4893 7973 4905 7976
rect 4939 7973 4951 8007
rect 4893 7967 4951 7973
rect 7653 8007 7711 8013
rect 7653 7973 7665 8007
rect 7699 8004 7711 8007
rect 8570 8004 8576 8016
rect 7699 7976 8576 8004
rect 7699 7973 7711 7976
rect 7653 7967 7711 7973
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 8662 7964 8668 8016
rect 8720 8004 8726 8016
rect 11072 8004 11100 8044
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12710 8072 12716 8084
rect 12671 8044 12716 8072
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13630 8072 13636 8084
rect 13035 8044 13636 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14829 8075 14887 8081
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 15194 8072 15200 8084
rect 14875 8044 15200 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 16850 8072 16856 8084
rect 16500 8044 16856 8072
rect 8720 7976 11100 8004
rect 11600 8007 11658 8013
rect 8720 7964 8726 7976
rect 11600 7973 11612 8007
rect 11646 8004 11658 8007
rect 11882 8004 11888 8016
rect 11646 7976 11888 8004
rect 11646 7973 11658 7976
rect 11600 7967 11658 7973
rect 11882 7964 11888 7976
rect 11940 7964 11946 8016
rect 13716 8007 13774 8013
rect 13716 7973 13728 8007
rect 13762 8004 13774 8007
rect 14642 8004 14648 8016
rect 13762 7976 14648 8004
rect 13762 7973 13774 7976
rect 13716 7967 13774 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15657 8007 15715 8013
rect 15657 7973 15669 8007
rect 15703 8004 15715 8007
rect 15703 7976 16252 8004
rect 15703 7973 15715 7976
rect 15657 7967 15715 7973
rect 4571 7908 4752 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 4856 7908 5457 7936
rect 4856 7896 4862 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 6730 7896 6736 7948
rect 6788 7936 6794 7948
rect 8386 7945 8392 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 6788 7908 8125 7936
rect 6788 7896 6794 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8380 7936 8392 7945
rect 8347 7908 8392 7936
rect 8113 7899 8171 7905
rect 8380 7899 8392 7908
rect 8386 7896 8392 7899
rect 8444 7896 8450 7948
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 9490 7936 9496 7948
rect 8812 7908 9496 7936
rect 8812 7896 8818 7908
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 10042 7896 10048 7948
rect 10100 7936 10106 7948
rect 13449 7939 13507 7945
rect 10100 7908 10145 7936
rect 10100 7896 10106 7908
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 13538 7936 13544 7948
rect 13495 7908 13544 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 14660 7936 14688 7964
rect 16224 7936 16252 7976
rect 16500 7936 16528 8044
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 17310 8072 17316 8084
rect 17271 8044 17316 8072
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 18322 8072 18328 8084
rect 17727 8044 18328 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 16666 8004 16672 8016
rect 16627 7976 16672 8004
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 16761 8007 16819 8013
rect 16761 7973 16773 8007
rect 16807 8004 16819 8007
rect 17770 8004 17776 8016
rect 16807 7976 17776 8004
rect 16807 7973 16819 7976
rect 16761 7967 16819 7973
rect 17770 7964 17776 7976
rect 17828 7964 17834 8016
rect 17402 7936 17408 7948
rect 14660 7908 15884 7936
rect 16224 7908 17408 7936
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2866 7868 2872 7880
rect 2639 7840 2872 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2866 7828 2872 7840
rect 2924 7868 2930 7880
rect 3605 7871 3663 7877
rect 2924 7840 3372 7868
rect 2924 7828 2930 7840
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 3344 7800 3372 7840
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 4614 7868 4620 7880
rect 3651 7840 4620 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 4724 7840 5641 7868
rect 4724 7800 4752 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 6638 7868 6644 7880
rect 6599 7840 6644 7868
rect 5629 7831 5687 7837
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7282 7868 7288 7880
rect 6871 7840 7288 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7524 7840 7849 7868
rect 7524 7828 7530 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9364 7840 10149 7868
rect 9364 7828 9370 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 8018 7800 8024 7812
rect 1627 7772 3004 7800
rect 3344 7772 4752 7800
rect 4816 7772 8024 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2866 7732 2872 7744
rect 1995 7704 2872 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 2976 7732 3004 7772
rect 3602 7732 3608 7744
rect 2976 7704 3608 7732
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 3789 7735 3847 7741
rect 3789 7701 3801 7735
rect 3835 7732 3847 7735
rect 4816 7732 4844 7772
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 9677 7803 9735 7809
rect 9677 7800 9689 7803
rect 9048 7772 9689 7800
rect 3835 7704 4844 7732
rect 3835 7701 3847 7704
rect 3789 7695 3847 7701
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 5074 7732 5080 7744
rect 4948 7704 4993 7732
rect 5035 7704 5080 7732
rect 4948 7692 4954 7704
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 5592 7704 6193 7732
rect 5592 7692 5598 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 6181 7695 6239 7701
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 9048 7732 9076 7772
rect 9677 7769 9689 7772
rect 9723 7769 9735 7803
rect 9677 7763 9735 7769
rect 9490 7732 9496 7744
rect 7984 7704 9076 7732
rect 9451 7704 9496 7732
rect 7984 7692 7990 7704
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 10244 7732 10272 7831
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 10560 7840 11345 7868
rect 10560 7828 10566 7840
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 15856 7877 15884 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 15712 7840 15761 7868
rect 15712 7828 15718 7840
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7868 15899 7871
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 15887 7840 16221 7868
rect 15887 7837 15899 7840
rect 15841 7831 15899 7837
rect 16209 7837 16221 7840
rect 16255 7868 16267 7871
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 16255 7840 16865 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 16853 7837 16865 7840
rect 16899 7837 16911 7871
rect 17770 7868 17776 7880
rect 17731 7840 17776 7868
rect 16853 7831 16911 7837
rect 17770 7828 17776 7840
rect 17828 7828 17834 7880
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 17920 7840 17965 7868
rect 17920 7828 17926 7840
rect 15289 7803 15347 7809
rect 15289 7769 15301 7803
rect 15335 7800 15347 7803
rect 17126 7800 17132 7812
rect 15335 7772 17132 7800
rect 15335 7769 15347 7772
rect 15289 7763 15347 7769
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 16206 7732 16212 7744
rect 9640 7704 10272 7732
rect 16167 7704 16212 7732
rect 9640 7692 9646 7704
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 16301 7735 16359 7741
rect 16301 7701 16313 7735
rect 16347 7732 16359 7735
rect 16850 7732 16856 7744
rect 16347 7704 16856 7732
rect 16347 7701 16359 7704
rect 16301 7695 16359 7701
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7528 3847 7531
rect 4706 7528 4712 7540
rect 3835 7500 4712 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 6273 7531 6331 7537
rect 6273 7528 6285 7531
rect 5316 7500 6285 7528
rect 5316 7488 5322 7500
rect 6273 7497 6285 7500
rect 6319 7497 6331 7531
rect 6273 7491 6331 7497
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 9306 7528 9312 7540
rect 7239 7500 9312 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 11882 7528 11888 7540
rect 9456 7500 11560 7528
rect 11843 7500 11888 7528
rect 9456 7488 9462 7500
rect 4890 7460 4896 7472
rect 3344 7432 4896 7460
rect 1394 7352 1400 7404
rect 1452 7392 1458 7404
rect 3344 7401 3372 7432
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 8662 7460 8668 7472
rect 6236 7432 8668 7460
rect 6236 7420 6242 7432
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1452 7364 1685 7392
rect 1452 7352 1458 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 1940 7327 1998 7333
rect 1940 7293 1952 7327
rect 1986 7324 1998 7327
rect 2958 7324 2964 7336
rect 1986 7296 2964 7324
rect 1986 7293 1998 7296
rect 1940 7287 1998 7293
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 4154 7324 4160 7336
rect 4115 7296 4160 7324
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4448 7324 4476 7355
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 7558 7392 7564 7404
rect 6604 7364 7564 7392
rect 6604 7352 6610 7364
rect 7558 7352 7564 7364
rect 7616 7392 7622 7404
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 7616 7364 7665 7392
rect 7616 7352 7622 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8202 7392 8208 7404
rect 7883 7364 8208 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 10502 7392 10508 7404
rect 10463 7364 10508 7392
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 11532 7392 11560 7500
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12710 7528 12716 7540
rect 12492 7500 12537 7528
rect 12636 7500 12716 7528
rect 12492 7488 12498 7500
rect 12250 7420 12256 7472
rect 12308 7460 12314 7472
rect 12636 7460 12664 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 16485 7531 16543 7537
rect 16485 7497 16497 7531
rect 16531 7497 16543 7531
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 16485 7491 16543 7497
rect 12308 7432 12664 7460
rect 12308 7420 12314 7432
rect 13170 7420 13176 7472
rect 13228 7460 13234 7472
rect 16500 7460 16528 7491
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 13228 7432 16528 7460
rect 13228 7420 13234 7432
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 11532 7364 12909 7392
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13998 7392 14004 7404
rect 13127 7364 14004 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 15102 7392 15108 7404
rect 15063 7364 15108 7392
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 16117 7395 16175 7401
rect 15344 7364 15884 7392
rect 15344 7352 15350 7364
rect 15856 7336 15884 7364
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16206 7392 16212 7404
rect 16163 7364 16212 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16540 7364 17049 7392
rect 16540 7352 16546 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 4614 7324 4620 7336
rect 4448 7296 4620 7324
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 4062 7216 4068 7268
rect 4120 7256 4126 7268
rect 4908 7256 4936 7287
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 7432 7296 8677 7324
rect 7432 7284 7438 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 8921 7327 8979 7333
rect 8921 7324 8933 7327
rect 8812 7296 8933 7324
rect 8812 7284 8818 7296
rect 8921 7293 8933 7296
rect 8967 7293 8979 7327
rect 8921 7287 8979 7293
rect 10772 7327 10830 7333
rect 10772 7293 10784 7327
rect 10818 7324 10830 7327
rect 12526 7324 12532 7336
rect 10818 7296 12532 7324
rect 10818 7293 10830 7296
rect 10772 7287 10830 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 13170 7324 13176 7336
rect 12636 7296 13176 7324
rect 4120 7228 4936 7256
rect 5160 7259 5218 7265
rect 4120 7216 4126 7228
rect 5160 7225 5172 7259
rect 5206 7256 5218 7259
rect 5350 7256 5356 7268
rect 5206 7228 5356 7256
rect 5206 7225 5218 7228
rect 5160 7219 5218 7225
rect 5350 7216 5356 7228
rect 5408 7256 5414 7268
rect 8294 7256 8300 7268
rect 5408 7228 8300 7256
rect 5408 7216 5414 7228
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 12636 7256 12664 7296
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 13630 7284 13636 7336
rect 13688 7324 13694 7336
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 13688 7296 13829 7324
rect 13688 7284 13694 7296
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14829 7327 14887 7333
rect 13964 7296 14009 7324
rect 13964 7284 13970 7296
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 15654 7324 15660 7336
rect 14875 7296 15660 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 14844 7256 14872 7287
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 15838 7324 15844 7336
rect 15751 7296 15844 7324
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 15933 7327 15991 7333
rect 15933 7293 15945 7327
rect 15979 7324 15991 7327
rect 16390 7324 16396 7336
rect 15979 7296 16396 7324
rect 15979 7293 15991 7296
rect 15933 7287 15991 7293
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 16850 7324 16856 7336
rect 16811 7296 16856 7324
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 16945 7259 17003 7265
rect 16945 7256 16957 7259
rect 8404 7228 12664 7256
rect 12728 7228 14872 7256
rect 15488 7228 16957 7256
rect 3050 7188 3056 7200
rect 3011 7160 3056 7188
rect 3050 7148 3056 7160
rect 3108 7148 3114 7200
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 4249 7191 4307 7197
rect 4249 7188 4261 7191
rect 3384 7160 4261 7188
rect 3384 7148 3390 7160
rect 4249 7157 4261 7160
rect 4295 7188 4307 7191
rect 6178 7188 6184 7200
rect 4295 7160 6184 7188
rect 4295 7157 4307 7160
rect 4249 7151 4307 7157
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 6730 7148 6736 7200
rect 6788 7188 6794 7200
rect 7561 7191 7619 7197
rect 7561 7188 7573 7191
rect 6788 7160 7573 7188
rect 6788 7148 6794 7160
rect 7561 7157 7573 7160
rect 7607 7157 7619 7191
rect 7561 7151 7619 7157
rect 8018 7148 8024 7200
rect 8076 7188 8082 7200
rect 8404 7188 8432 7228
rect 8076 7160 8432 7188
rect 8076 7148 8082 7160
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 9824 7160 10057 7188
rect 9824 7148 9830 7160
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 10045 7151 10103 7157
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12728 7188 12756 7228
rect 12032 7160 12756 7188
rect 12805 7191 12863 7197
rect 12032 7148 12038 7160
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 13814 7188 13820 7200
rect 12851 7160 13820 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 14918 7188 14924 7200
rect 14792 7160 14924 7188
rect 14792 7148 14798 7160
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 15488 7197 15516 7228
rect 16945 7225 16957 7228
rect 16991 7225 17003 7259
rect 16945 7219 17003 7225
rect 15473 7191 15531 7197
rect 15473 7157 15485 7191
rect 15519 7157 15531 7191
rect 15473 7151 15531 7157
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 18064 7188 18092 7287
rect 15896 7160 18092 7188
rect 15896 7148 15902 7160
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 1104 7024 18860 7046
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 4982 6984 4988 6996
rect 4396 6956 4988 6984
rect 4396 6944 4402 6956
rect 4982 6944 4988 6956
rect 5040 6984 5046 6996
rect 5258 6984 5264 6996
rect 5040 6956 5264 6984
rect 5040 6944 5046 6956
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 6638 6984 6644 6996
rect 6411 6956 6644 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8757 6987 8815 6993
rect 8757 6984 8769 6987
rect 8352 6956 8769 6984
rect 8352 6944 8358 6956
rect 8757 6953 8769 6956
rect 8803 6984 8815 6987
rect 9582 6984 9588 6996
rect 8803 6956 9588 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6953 9919 6987
rect 9861 6947 9919 6953
rect 3142 6876 3148 6928
rect 3200 6916 3206 6928
rect 3881 6919 3939 6925
rect 3881 6916 3893 6919
rect 3200 6888 3893 6916
rect 3200 6876 3206 6888
rect 3881 6885 3893 6888
rect 3927 6885 3939 6919
rect 8846 6916 8852 6928
rect 3881 6879 3939 6885
rect 6840 6888 8852 6916
rect 1670 6848 1676 6860
rect 1631 6820 1676 6848
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 2584 6851 2642 6857
rect 2584 6817 2596 6851
rect 2630 6848 2642 6851
rect 3050 6848 3056 6860
rect 2630 6820 3056 6848
rect 2630 6817 2642 6820
rect 2584 6811 2642 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 4332 6851 4390 6857
rect 4332 6848 4344 6851
rect 3712 6820 4344 6848
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 2314 6780 2320 6792
rect 1452 6752 2320 6780
rect 1452 6740 1458 6752
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 3712 6721 3740 6820
rect 4332 6817 4344 6820
rect 4378 6848 4390 6851
rect 5350 6848 5356 6860
rect 4378 6820 5356 6848
rect 4378 6817 4390 6820
rect 4332 6811 4390 6817
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 6733 6851 6791 6857
rect 6733 6817 6745 6851
rect 6779 6848 6791 6851
rect 6840 6848 6868 6888
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 9876 6916 9904 6947
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 11701 6987 11759 6993
rect 10652 6956 11008 6984
rect 10652 6944 10658 6956
rect 10980 6928 11008 6956
rect 11701 6953 11713 6987
rect 11747 6984 11759 6987
rect 12342 6984 12348 6996
rect 11747 6956 12348 6984
rect 11747 6953 11759 6956
rect 11701 6947 11759 6953
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12710 6984 12716 6996
rect 12623 6956 12716 6984
rect 12710 6944 12716 6956
rect 12768 6984 12774 6996
rect 13262 6984 13268 6996
rect 12768 6956 13268 6984
rect 12768 6944 12774 6956
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 14458 6984 14464 6996
rect 13771 6956 14464 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 15252 6956 15669 6984
rect 15252 6944 15258 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 16758 6984 16764 6996
rect 16719 6956 16764 6984
rect 15657 6947 15715 6953
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 17865 6987 17923 6993
rect 17865 6953 17877 6987
rect 17911 6984 17923 6987
rect 18138 6984 18144 6996
rect 17911 6956 18144 6984
rect 17911 6953 17923 6956
rect 17865 6947 17923 6953
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 10502 6916 10508 6928
rect 9876 6888 10508 6916
rect 7466 6848 7472 6860
rect 6779 6820 6868 6848
rect 7024 6820 7472 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 4062 6780 4068 6792
rect 3927 6752 4068 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 3697 6715 3755 6721
rect 3697 6681 3709 6715
rect 3743 6681 3755 6715
rect 5736 6712 5764 6811
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 5994 6780 6000 6792
rect 5868 6752 6000 6780
rect 5868 6740 5874 6752
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6822 6780 6828 6792
rect 6783 6752 6828 6780
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7024 6789 7052 6820
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7644 6851 7702 6857
rect 7644 6817 7656 6851
rect 7690 6848 7702 6851
rect 8202 6848 8208 6860
rect 7690 6820 8208 6848
rect 7690 6817 7702 6820
rect 7644 6811 7702 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10336 6857 10364 6888
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 10962 6876 10968 6928
rect 11020 6916 11026 6928
rect 11974 6916 11980 6928
rect 11020 6888 11980 6916
rect 11020 6876 11026 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 12084 6888 13032 6916
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 10588 6851 10646 6857
rect 10588 6817 10600 6851
rect 10634 6848 10646 6851
rect 12084 6848 12112 6888
rect 10634 6820 12112 6848
rect 12161 6851 12219 6857
rect 10634 6817 10646 6820
rect 10588 6811 10646 6817
rect 12161 6817 12173 6851
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 13004 6848 13032 6888
rect 15562 6876 15568 6928
rect 15620 6916 15626 6928
rect 15620 6888 15792 6916
rect 15620 6876 15626 6888
rect 13004 6820 14044 6848
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7374 6780 7380 6792
rect 7335 6752 7380 6780
rect 7009 6743 7067 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 12176 6780 12204 6811
rect 11572 6752 12204 6780
rect 11572 6740 11578 6752
rect 12250 6740 12256 6792
rect 12308 6780 12314 6792
rect 12802 6780 12808 6792
rect 12308 6752 12664 6780
rect 12763 6752 12808 6780
rect 12308 6740 12314 6752
rect 12636 6712 12664 6752
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 13004 6789 13032 6820
rect 14016 6792 14044 6820
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 15764 6848 15792 6888
rect 16574 6876 16580 6928
rect 16632 6916 16638 6928
rect 16669 6919 16727 6925
rect 16669 6916 16681 6919
rect 16632 6888 16681 6916
rect 16632 6876 16638 6888
rect 16669 6885 16681 6888
rect 16715 6885 16727 6919
rect 16669 6879 16727 6885
rect 14792 6820 15516 6848
rect 15764 6820 16344 6848
rect 14792 6808 14798 6820
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13722 6780 13728 6792
rect 13136 6752 13728 6780
rect 13136 6740 13142 6752
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13817 6743 13875 6749
rect 13832 6712 13860 6743
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 15102 6780 15108 6792
rect 14516 6752 15108 6780
rect 14516 6740 14522 6752
rect 15102 6740 15108 6752
rect 15160 6780 15166 6792
rect 15488 6780 15516 6820
rect 15749 6783 15807 6789
rect 15749 6780 15761 6783
rect 15160 6752 15424 6780
rect 15488 6752 15761 6780
rect 15160 6740 15166 6752
rect 15289 6715 15347 6721
rect 15289 6712 15301 6715
rect 3697 6675 3755 6681
rect 5000 6684 5580 6712
rect 5736 6684 7420 6712
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 2958 6644 2964 6656
rect 1903 6616 2964 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3786 6604 3792 6656
rect 3844 6644 3850 6656
rect 5000 6644 5028 6684
rect 3844 6616 5028 6644
rect 3844 6604 3850 6616
rect 5166 6604 5172 6656
rect 5224 6644 5230 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5224 6616 5457 6644
rect 5224 6604 5230 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5552 6644 5580 6684
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5552 6616 5917 6644
rect 5445 6607 5503 6613
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 7392 6644 7420 6684
rect 8680 6684 10364 6712
rect 8680 6644 8708 6684
rect 7392 6616 8708 6644
rect 10336 6644 10364 6684
rect 11256 6684 12572 6712
rect 12636 6684 13768 6712
rect 13832 6684 15301 6712
rect 11256 6644 11284 6684
rect 11974 6644 11980 6656
rect 10336 6616 11284 6644
rect 11935 6616 11980 6644
rect 5905 6607 5963 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12342 6644 12348 6656
rect 12303 6616 12348 6644
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12544 6644 12572 6684
rect 13078 6644 13084 6656
rect 12544 6616 13084 6644
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13354 6644 13360 6656
rect 13315 6616 13360 6644
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13740 6644 13768 6684
rect 15289 6681 15301 6684
rect 15335 6681 15347 6715
rect 15396 6712 15424 6752
rect 15749 6749 15761 6752
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 15856 6712 15884 6743
rect 16316 6721 16344 6820
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17957 6851 18015 6857
rect 17957 6848 17969 6851
rect 17000 6820 17969 6848
rect 17000 6808 17006 6820
rect 17957 6817 17969 6820
rect 18003 6817 18015 6851
rect 17957 6811 18015 6817
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6780 16911 6783
rect 17586 6780 17592 6792
rect 16899 6752 17592 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 17862 6740 17868 6792
rect 17920 6780 17926 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17920 6752 18061 6780
rect 17920 6740 17926 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 15396 6684 15884 6712
rect 16301 6715 16359 6721
rect 15289 6675 15347 6681
rect 16301 6681 16313 6715
rect 16347 6681 16359 6715
rect 17494 6712 17500 6724
rect 17455 6684 17500 6712
rect 16301 6675 16359 6681
rect 17494 6672 17500 6684
rect 17552 6672 17558 6724
rect 15654 6644 15660 6656
rect 13740 6616 15660 6644
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 3142 6440 3148 6452
rect 2372 6412 3148 6440
rect 2372 6400 2378 6412
rect 3142 6400 3148 6412
rect 3200 6440 3206 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3200 6412 3433 6440
rect 3200 6400 3206 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 3421 6403 3479 6409
rect 4430 6400 4436 6452
rect 4488 6440 4494 6452
rect 5074 6440 5080 6452
rect 4488 6412 5080 6440
rect 4488 6400 4494 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 6730 6440 6736 6452
rect 5316 6412 6736 6440
rect 5316 6400 5322 6412
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 8202 6440 8208 6452
rect 6880 6412 8064 6440
rect 8163 6412 8208 6440
rect 6880 6400 6886 6412
rect 3329 6375 3387 6381
rect 3329 6341 3341 6375
rect 3375 6372 3387 6375
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3375 6344 3801 6372
rect 3375 6341 3387 6344
rect 3329 6335 3387 6341
rect 3789 6341 3801 6344
rect 3835 6341 3847 6375
rect 3789 6335 3847 6341
rect 4246 6332 4252 6384
rect 4304 6372 4310 6384
rect 5997 6375 6055 6381
rect 5997 6372 6009 6375
rect 4304 6344 6009 6372
rect 4304 6332 4310 6344
rect 5997 6341 6009 6344
rect 6043 6341 6055 6375
rect 8036 6372 8064 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9398 6440 9404 6452
rect 9140 6412 9404 6440
rect 8662 6372 8668 6384
rect 8036 6344 8668 6372
rect 5997 6335 6055 6341
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2590 6304 2596 6316
rect 2087 6276 2596 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3053 6307 3111 6313
rect 2924 6276 2969 6304
rect 2924 6264 2930 6276
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3142 6304 3148 6316
rect 3099 6276 3148 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3476 6276 3709 6304
rect 3476 6264 3482 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 4430 6304 4436 6316
rect 4391 6276 4436 6304
rect 3697 6267 3755 6273
rect 4430 6264 4436 6276
rect 4488 6304 4494 6316
rect 5166 6304 5172 6316
rect 4488 6276 5172 6304
rect 4488 6264 4494 6276
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 5350 6304 5356 6316
rect 5311 6276 5356 6304
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5828 6276 6960 6304
rect 2774 6236 2780 6248
rect 2735 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 3605 6239 3663 6245
rect 3605 6205 3617 6239
rect 3651 6236 3663 6239
rect 5261 6239 5319 6245
rect 3651 6208 5212 6236
rect 3651 6205 3663 6208
rect 3605 6199 3663 6205
rect 1857 6171 1915 6177
rect 1857 6137 1869 6171
rect 1903 6168 1915 6171
rect 3329 6171 3387 6177
rect 3329 6168 3341 6171
rect 1903 6140 3341 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 3329 6137 3341 6140
rect 3375 6137 3387 6171
rect 5184 6168 5212 6208
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5626 6236 5632 6248
rect 5307 6208 5632 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 5828 6245 5856 6276
rect 5813 6239 5871 6245
rect 5813 6205 5825 6239
rect 5859 6205 5871 6239
rect 5813 6199 5871 6205
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6205 6883 6239
rect 6932 6236 6960 6276
rect 9140 6236 9168 6412
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 12066 6440 12072 6452
rect 11379 6412 12072 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 13081 6443 13139 6449
rect 13081 6440 13093 6443
rect 12860 6412 13093 6440
rect 12860 6400 12866 6412
rect 13081 6409 13093 6412
rect 13127 6409 13139 6443
rect 13081 6403 13139 6409
rect 13998 6400 14004 6452
rect 14056 6440 14062 6452
rect 15473 6443 15531 6449
rect 15473 6440 15485 6443
rect 14056 6412 15485 6440
rect 14056 6400 14062 6412
rect 15473 6409 15485 6412
rect 15519 6409 15531 6443
rect 17586 6440 17592 6452
rect 17547 6412 17592 6440
rect 15473 6403 15531 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 18230 6440 18236 6452
rect 18191 6412 18236 6440
rect 18230 6400 18236 6412
rect 18288 6400 18294 6452
rect 13354 6372 13360 6384
rect 11808 6344 13360 6372
rect 11808 6313 11836 6344
rect 13354 6332 13360 6344
rect 13412 6332 13418 6384
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12434 6304 12440 6316
rect 12023 6276 12440 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 13998 6304 14004 6316
rect 13771 6276 14004 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 15160 6276 16313 6304
rect 15160 6264 15166 6276
rect 16301 6273 16313 6276
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 16408 6276 18092 6304
rect 6932 6208 9168 6236
rect 9217 6239 9275 6245
rect 6825 6199 6883 6205
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 10502 6236 10508 6248
rect 9263 6208 10508 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 5350 6168 5356 6180
rect 5184 6140 5356 6168
rect 3329 6131 3387 6137
rect 5350 6128 5356 6140
rect 5408 6168 5414 6180
rect 6656 6168 6684 6199
rect 5408 6140 6684 6168
rect 5408 6128 5414 6140
rect 1397 6103 1455 6109
rect 1397 6069 1409 6103
rect 1443 6100 1455 6103
rect 1486 6100 1492 6112
rect 1443 6072 1492 6100
rect 1443 6069 1455 6072
rect 1397 6063 1455 6069
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 1762 6100 1768 6112
rect 1723 6072 1768 6100
rect 1762 6060 1768 6072
rect 1820 6060 1826 6112
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2409 6103 2467 6109
rect 2409 6100 2421 6103
rect 2096 6072 2421 6100
rect 2096 6060 2102 6072
rect 2409 6069 2421 6072
rect 2455 6069 2467 6103
rect 2409 6063 2467 6069
rect 3697 6103 3755 6109
rect 3697 6069 3709 6103
rect 3743 6100 3755 6103
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 3743 6072 4169 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 4157 6069 4169 6072
rect 4203 6069 4215 6103
rect 4157 6063 4215 6069
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4295 6072 4813 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5810 6100 5816 6112
rect 5215 6072 5816 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5810 6060 5816 6072
rect 5868 6100 5874 6112
rect 6086 6100 6092 6112
rect 5868 6072 6092 6100
rect 5868 6060 5874 6072
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 6546 6100 6552 6112
rect 6503 6072 6552 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 6546 6060 6552 6072
rect 6604 6100 6610 6112
rect 6840 6100 6868 6199
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6236 11759 6239
rect 12342 6236 12348 6248
rect 11747 6208 12348 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13688 6208 14105 6236
rect 13688 6196 13694 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 16408 6236 16436 6276
rect 14093 6199 14151 6205
rect 14200 6208 16436 6236
rect 6914 6128 6920 6180
rect 6972 6128 6978 6180
rect 7092 6171 7150 6177
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 7282 6168 7288 6180
rect 7138 6140 7288 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 7282 6128 7288 6140
rect 7340 6128 7346 6180
rect 7926 6128 7932 6180
rect 7984 6168 7990 6180
rect 8294 6168 8300 6180
rect 7984 6140 8300 6168
rect 7984 6128 7990 6140
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 9484 6171 9542 6177
rect 9484 6137 9496 6171
rect 9530 6168 9542 6171
rect 9766 6168 9772 6180
rect 9530 6140 9772 6168
rect 9530 6137 9542 6140
rect 9484 6131 9542 6137
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 11790 6128 11796 6180
rect 11848 6168 11854 6180
rect 12066 6168 12072 6180
rect 11848 6140 12072 6168
rect 11848 6128 11854 6140
rect 12066 6128 12072 6140
rect 12124 6128 12130 6180
rect 13449 6171 13507 6177
rect 13449 6168 13461 6171
rect 12176 6140 13461 6168
rect 6604 6072 6868 6100
rect 6932 6100 6960 6128
rect 12176 6112 12204 6140
rect 13449 6137 13461 6140
rect 13495 6137 13507 6171
rect 13449 6131 13507 6137
rect 13814 6128 13820 6180
rect 13872 6168 13878 6180
rect 14200 6168 14228 6208
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 18064 6245 18092 6276
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 16632 6208 17417 6236
rect 16632 6196 16638 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 13872 6140 14228 6168
rect 14360 6171 14418 6177
rect 13872 6128 13878 6140
rect 14360 6137 14372 6171
rect 14406 6168 14418 6171
rect 14458 6168 14464 6180
rect 14406 6140 14464 6168
rect 14406 6137 14418 6140
rect 14360 6131 14418 6137
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 16117 6171 16175 6177
rect 14568 6140 15884 6168
rect 8202 6100 8208 6112
rect 6932 6072 8208 6100
rect 6604 6060 6610 6072
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8757 6103 8815 6109
rect 8757 6069 8769 6103
rect 8803 6100 8815 6103
rect 8938 6100 8944 6112
rect 8803 6072 8944 6100
rect 8803 6069 8815 6072
rect 8757 6063 8815 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 11238 6100 11244 6112
rect 10643 6072 11244 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 12158 6060 12164 6112
rect 12216 6060 12222 6112
rect 13170 6060 13176 6112
rect 13228 6100 13234 6112
rect 13538 6100 13544 6112
rect 13228 6072 13544 6100
rect 13228 6060 13234 6072
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14568 6100 14596 6140
rect 13780 6072 14596 6100
rect 13780 6060 13786 6072
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 15252 6072 15761 6100
rect 15252 6060 15258 6072
rect 15749 6069 15761 6072
rect 15795 6069 15807 6103
rect 15856 6100 15884 6140
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 17034 6168 17040 6180
rect 16163 6140 17040 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 17034 6128 17040 6140
rect 17092 6128 17098 6180
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 15856 6072 16221 6100
rect 15749 6063 15807 6069
rect 16209 6069 16221 6072
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 4157 5899 4215 5905
rect 4157 5896 4169 5899
rect 1820 5868 4169 5896
rect 1820 5856 1826 5868
rect 4157 5865 4169 5868
rect 4203 5865 4215 5899
rect 4614 5896 4620 5908
rect 4575 5868 4620 5896
rect 4157 5859 4215 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5258 5896 5264 5908
rect 5219 5868 5264 5896
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7282 5896 7288 5908
rect 6963 5868 7288 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 7524 5868 9229 5896
rect 7524 5856 7530 5868
rect 9217 5865 9229 5868
rect 9263 5865 9275 5899
rect 11882 5896 11888 5908
rect 9217 5859 9275 5865
rect 10060 5868 11888 5896
rect 5804 5831 5862 5837
rect 5804 5797 5816 5831
rect 5850 5828 5862 5831
rect 7484 5828 7512 5856
rect 10060 5828 10088 5868
rect 11882 5856 11888 5868
rect 11940 5896 11946 5908
rect 12250 5896 12256 5908
rect 11940 5868 12256 5896
rect 11940 5856 11946 5868
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 13998 5896 14004 5908
rect 13504 5868 13768 5896
rect 13911 5868 14004 5896
rect 13504 5856 13510 5868
rect 10502 5828 10508 5840
rect 5850 5800 7512 5828
rect 8036 5800 10088 5828
rect 10152 5800 10508 5828
rect 5850 5797 5862 5800
rect 5804 5791 5862 5797
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1581 5763 1639 5769
rect 1581 5760 1593 5763
rect 1452 5732 1593 5760
rect 1452 5720 1458 5732
rect 1581 5729 1593 5732
rect 1627 5729 1639 5763
rect 1581 5723 1639 5729
rect 1848 5763 1906 5769
rect 1848 5729 1860 5763
rect 1894 5760 1906 5763
rect 3237 5763 3295 5769
rect 1894 5732 3188 5760
rect 1894 5729 1906 5732
rect 1848 5723 1906 5729
rect 3160 5624 3188 5732
rect 3237 5729 3249 5763
rect 3283 5729 3295 5763
rect 3237 5723 3295 5729
rect 3252 5692 3280 5723
rect 3694 5720 3700 5772
rect 3752 5760 3758 5772
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 3752 5732 4537 5760
rect 3752 5720 3758 5732
rect 4525 5729 4537 5732
rect 4571 5760 4583 5763
rect 5258 5760 5264 5772
rect 4571 5732 5264 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 6546 5760 6552 5772
rect 5583 5732 6552 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 4338 5692 4344 5704
rect 3252 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4522 5624 4528 5636
rect 3160 5596 4528 5624
rect 4522 5584 4528 5596
rect 4580 5624 4586 5636
rect 4724 5624 4752 5655
rect 4580 5596 4752 5624
rect 4580 5584 4586 5596
rect 2590 5516 2596 5568
rect 2648 5556 2654 5568
rect 2961 5559 3019 5565
rect 2961 5556 2973 5559
rect 2648 5528 2973 5556
rect 2648 5516 2654 5528
rect 2961 5525 2973 5528
rect 3007 5525 3019 5559
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 2961 5519 3019 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5258 5556 5264 5568
rect 4948 5528 5264 5556
rect 4948 5516 4954 5528
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 5460 5556 5488 5723
rect 6546 5720 6552 5732
rect 6604 5760 6610 5772
rect 7190 5760 7196 5772
rect 6604 5732 7052 5760
rect 7151 5732 7196 5760
rect 6604 5720 6610 5732
rect 7024 5692 7052 5732
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 8036 5760 8064 5800
rect 7340 5732 8064 5760
rect 8104 5763 8162 5769
rect 7340 5720 7346 5732
rect 8104 5729 8116 5763
rect 8150 5760 8162 5763
rect 9582 5760 9588 5772
rect 8150 5732 9588 5760
rect 8150 5729 8162 5732
rect 8104 5723 8162 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 10152 5769 10180 5800
rect 10502 5788 10508 5800
rect 10560 5788 10566 5840
rect 13740 5828 13768 5868
rect 13998 5856 14004 5868
rect 14056 5896 14062 5908
rect 14458 5896 14464 5908
rect 14056 5868 14464 5896
rect 14056 5856 14062 5868
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 18046 5896 18052 5908
rect 18007 5868 18052 5896
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 13740 5800 17356 5828
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10404 5763 10462 5769
rect 10404 5729 10416 5763
rect 10450 5760 10462 5763
rect 11238 5760 11244 5772
rect 10450 5732 11244 5760
rect 10450 5729 10462 5732
rect 10404 5723 10462 5729
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 12888 5763 12946 5769
rect 12888 5729 12900 5763
rect 12934 5760 12946 5763
rect 13722 5760 13728 5772
rect 12934 5732 13728 5760
rect 12934 5729 12946 5732
rect 12888 5723 12946 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5760 14795 5763
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 14783 5732 15669 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 15657 5729 15669 5732
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 16666 5720 16672 5772
rect 16724 5760 16730 5772
rect 17328 5769 17356 5800
rect 16761 5763 16819 5769
rect 16761 5760 16773 5763
rect 16724 5732 16773 5760
rect 16724 5720 16730 5732
rect 16761 5729 16773 5732
rect 16807 5729 16819 5763
rect 16761 5723 16819 5729
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5729 17371 5763
rect 17313 5723 17371 5729
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 7374 5692 7380 5704
rect 7024 5664 7380 5692
rect 7374 5652 7380 5664
rect 7432 5692 7438 5704
rect 7834 5692 7840 5704
rect 7432 5664 7840 5692
rect 7432 5652 7438 5664
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 12492 5664 12633 5692
rect 12492 5652 12498 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 12621 5655 12679 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 16206 5692 16212 5704
rect 15979 5664 16212 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 17880 5692 17908 5723
rect 16356 5664 17908 5692
rect 16356 5652 16362 5664
rect 7650 5624 7656 5636
rect 7208 5596 7656 5624
rect 7208 5556 7236 5596
rect 7650 5584 7656 5596
rect 7708 5584 7714 5636
rect 11698 5624 11704 5636
rect 11440 5596 11704 5624
rect 7374 5556 7380 5568
rect 5460 5528 7236 5556
rect 7335 5528 7380 5556
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 11440 5556 11468 5596
rect 11698 5584 11704 5596
rect 11756 5624 11762 5636
rect 12158 5624 12164 5636
rect 11756 5596 12164 5624
rect 11756 5584 11762 5596
rect 12158 5584 12164 5596
rect 12216 5584 12222 5636
rect 17494 5624 17500 5636
rect 17455 5596 17500 5624
rect 17494 5584 17500 5596
rect 17552 5584 17558 5636
rect 8260 5528 11468 5556
rect 11517 5559 11575 5565
rect 8260 5516 8266 5528
rect 11517 5525 11529 5559
rect 11563 5556 11575 5559
rect 11882 5556 11888 5568
rect 11563 5528 11888 5556
rect 11563 5525 11575 5528
rect 11517 5519 11575 5525
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 16942 5556 16948 5568
rect 16903 5528 16948 5556
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 4246 5352 4252 5364
rect 3752 5324 4252 5352
rect 3752 5312 3758 5324
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 6089 5355 6147 5361
rect 6089 5352 6101 5355
rect 5224 5324 6101 5352
rect 5224 5312 5230 5324
rect 6089 5321 6101 5324
rect 6135 5321 6147 5355
rect 6089 5315 6147 5321
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 7837 5355 7895 5361
rect 6328 5324 7420 5352
rect 6328 5312 6334 5324
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5176 1458 5228
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 4430 5216 4436 5228
rect 2648 5188 4436 5216
rect 2648 5176 2654 5188
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4522 5176 4528 5228
rect 4580 5216 4586 5228
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 4580 5188 5457 5216
rect 4580 5176 4586 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 6730 5216 6736 5228
rect 5445 5179 5503 5185
rect 5644 5188 6736 5216
rect 1664 5151 1722 5157
rect 1664 5117 1676 5151
rect 1710 5148 1722 5151
rect 2608 5148 2636 5176
rect 3050 5148 3056 5160
rect 1710 5120 2636 5148
rect 3011 5120 3056 5148
rect 1710 5117 1722 5120
rect 1664 5111 1722 5117
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 5644 5148 5672 5188
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7392 5225 7420 5324
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 7883 5324 8677 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 8665 5321 8677 5324
rect 8711 5321 8723 5355
rect 8846 5352 8852 5364
rect 8807 5324 8852 5352
rect 8665 5315 8723 5321
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10226 5352 10232 5364
rect 9907 5324 10232 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 11808 5324 13676 5352
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 11422 5284 11428 5296
rect 7524 5256 11428 5284
rect 7524 5244 7530 5256
rect 11422 5244 11428 5256
rect 11480 5244 11486 5296
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5185 7435 5219
rect 8294 5216 8300 5228
rect 8255 5188 8300 5216
rect 7377 5179 7435 5185
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 3896 5120 5672 5148
rect 5905 5151 5963 5157
rect 3142 5040 3148 5092
rect 3200 5080 3206 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 3200 5052 3341 5080
rect 3200 5040 3206 5052
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 3329 5043 3387 5049
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 3896 5021 3924 5120
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 6454 5148 6460 5160
rect 5951 5120 6460 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 6564 5120 7205 5148
rect 4246 5080 4252 5092
rect 4207 5052 4252 5080
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 6564 5080 6592 5120
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 8202 5148 8208 5160
rect 7616 5120 8208 5148
rect 7616 5108 7622 5120
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 4908 5052 6592 5080
rect 3881 5015 3939 5021
rect 2832 4984 2877 5012
rect 2832 4972 2838 4984
rect 3881 4981 3893 5015
rect 3927 4981 3939 5015
rect 3881 4975 3939 4981
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4522 5012 4528 5024
rect 4387 4984 4528 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4522 4972 4528 4984
rect 4580 4972 4586 5024
rect 4908 5021 4936 5052
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 6972 5052 7297 5080
rect 6972 5040 6978 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 7285 5043 7343 5049
rect 4893 5015 4951 5021
rect 4893 4981 4905 5015
rect 4939 4981 4951 5015
rect 5258 5012 5264 5024
rect 5219 4984 5264 5012
rect 4893 4975 4951 4981
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 5353 5015 5411 5021
rect 5353 4981 5365 5015
rect 5399 5012 5411 5015
rect 5442 5012 5448 5024
rect 5399 4984 5448 5012
rect 5399 4981 5411 4984
rect 5353 4975 5411 4981
rect 5442 4972 5448 4984
rect 5500 5012 5506 5024
rect 6270 5012 6276 5024
rect 5500 4984 6276 5012
rect 5500 4972 5506 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 6825 5015 6883 5021
rect 6825 5012 6837 5015
rect 6604 4984 6837 5012
rect 6604 4972 6610 4984
rect 6825 4981 6837 4984
rect 6871 4981 6883 5015
rect 6825 4975 6883 4981
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8404 5012 8432 5179
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 9493 5219 9551 5225
rect 8812 5188 9352 5216
rect 8812 5176 8818 5188
rect 9214 5148 9220 5160
rect 9175 5120 9220 5148
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9324 5148 9352 5188
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9582 5216 9588 5228
rect 9539 5188 9588 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9582 5176 9588 5188
rect 9640 5216 9646 5228
rect 11808 5225 11836 5324
rect 13648 5284 13676 5324
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13780 5324 13829 5352
rect 13780 5312 13786 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 13817 5315 13875 5321
rect 13924 5324 16037 5352
rect 13924 5284 13952 5324
rect 16025 5321 16037 5324
rect 16071 5321 16083 5355
rect 16025 5315 16083 5321
rect 13648 5256 13952 5284
rect 15470 5244 15476 5296
rect 15528 5284 15534 5296
rect 15528 5256 18092 5284
rect 15528 5244 15534 5256
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 9640 5188 10425 5216
rect 9640 5176 9646 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12023 5188 12572 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9324 5120 10241 5148
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 10778 5148 10784 5160
rect 10275 5120 10784 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 12434 5148 12440 5160
rect 11348 5120 12204 5148
rect 12395 5120 12440 5148
rect 8665 5083 8723 5089
rect 8665 5049 8677 5083
rect 8711 5080 8723 5083
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 8711 5052 9321 5080
rect 8711 5049 8723 5052
rect 8665 5043 8723 5049
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9309 5043 9367 5049
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 9456 5052 10272 5080
rect 9456 5040 9462 5052
rect 10244 5024 10272 5052
rect 8352 4984 8432 5012
rect 8352 4972 8358 4984
rect 10226 4972 10232 5024
rect 10284 4972 10290 5024
rect 10318 4972 10324 5024
rect 10376 5012 10382 5024
rect 10870 5012 10876 5024
rect 10376 4984 10421 5012
rect 10831 4984 10876 5012
rect 10376 4972 10382 4984
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 11348 5021 11376 5120
rect 11701 5083 11759 5089
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 12176 5080 12204 5120
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12544 5148 12572 5188
rect 16206 5176 16212 5228
rect 16264 5216 16270 5228
rect 16577 5219 16635 5225
rect 16577 5216 16589 5219
rect 16264 5188 16589 5216
rect 16264 5176 16270 5188
rect 16577 5185 16589 5188
rect 16623 5185 16635 5219
rect 16577 5179 16635 5185
rect 12544 5120 12747 5148
rect 12526 5080 12532 5092
rect 11747 5052 12112 5080
rect 12176 5052 12532 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 11333 5015 11391 5021
rect 11333 4981 11345 5015
rect 11379 4981 11391 5015
rect 12084 5012 12112 5052
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 12719 5089 12747 5120
rect 13630 5108 13636 5160
rect 13688 5148 13694 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 13688 5120 14381 5148
rect 13688 5108 13694 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 14636 5151 14694 5157
rect 14636 5148 14648 5151
rect 14516 5120 14648 5148
rect 14516 5108 14522 5120
rect 14636 5117 14648 5120
rect 14682 5148 14694 5151
rect 16224 5148 16252 5176
rect 17402 5148 17408 5160
rect 14682 5120 16252 5148
rect 17363 5120 17408 5148
rect 14682 5117 14694 5120
rect 14636 5111 14694 5117
rect 17402 5108 17408 5120
rect 17460 5108 17466 5160
rect 18064 5157 18092 5256
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 12704 5083 12762 5089
rect 12704 5049 12716 5083
rect 12750 5080 12762 5083
rect 13262 5080 13268 5092
rect 12750 5052 13268 5080
rect 12750 5049 12762 5052
rect 12704 5043 12762 5049
rect 13262 5040 13268 5052
rect 13320 5080 13326 5092
rect 16393 5083 16451 5089
rect 13320 5052 15792 5080
rect 13320 5040 13326 5052
rect 15286 5012 15292 5024
rect 12084 4984 15292 5012
rect 11333 4975 11391 4981
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 15764 5021 15792 5052
rect 16393 5049 16405 5083
rect 16439 5080 16451 5083
rect 16574 5080 16580 5092
rect 16439 5052 16580 5080
rect 16439 5049 16451 5052
rect 16393 5043 16451 5049
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 15749 5015 15807 5021
rect 15749 4981 15761 5015
rect 15795 4981 15807 5015
rect 16482 5012 16488 5024
rect 16443 4984 16488 5012
rect 15749 4975 15807 4981
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 17586 5012 17592 5024
rect 17547 4984 17592 5012
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 6178 4808 6184 4820
rect 6139 4780 6184 4808
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 6270 4768 6276 4820
rect 6328 4808 6334 4820
rect 9030 4808 9036 4820
rect 6328 4780 9036 4808
rect 6328 4768 6334 4780
rect 9030 4768 9036 4780
rect 9088 4808 9094 4820
rect 10594 4808 10600 4820
rect 9088 4780 10600 4808
rect 9088 4768 9094 4780
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 10870 4768 10876 4820
rect 10928 4808 10934 4820
rect 11701 4811 11759 4817
rect 11701 4808 11713 4811
rect 10928 4780 11713 4808
rect 10928 4768 10934 4780
rect 11701 4777 11713 4780
rect 11747 4777 11759 4811
rect 12066 4808 12072 4820
rect 11701 4771 11759 4777
rect 11808 4780 12072 4808
rect 4246 4740 4252 4752
rect 1504 4712 4252 4740
rect 1504 4681 1532 4712
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 4430 4700 4436 4752
rect 4488 4740 4494 4752
rect 6089 4743 6147 4749
rect 6089 4740 6101 4743
rect 4488 4712 6101 4740
rect 4488 4700 4494 4712
rect 6089 4709 6101 4712
rect 6135 4709 6147 4743
rect 6089 4703 6147 4709
rect 7193 4743 7251 4749
rect 7193 4709 7205 4743
rect 7239 4740 7251 4743
rect 7466 4740 7472 4752
rect 7239 4712 7472 4740
rect 7239 4709 7251 4712
rect 7193 4703 7251 4709
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 8104 4743 8162 4749
rect 8104 4709 8116 4743
rect 8150 4740 8162 4743
rect 8294 4740 8300 4752
rect 8150 4712 8300 4740
rect 8150 4709 8162 4712
rect 8104 4703 8162 4709
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 10502 4740 10508 4752
rect 9692 4712 10508 4740
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 2308 4675 2366 4681
rect 2308 4641 2320 4675
rect 2354 4672 2366 4675
rect 2774 4672 2780 4684
rect 2354 4644 2780 4672
rect 2354 4641 2366 4644
rect 2308 4635 2366 4641
rect 2774 4632 2780 4644
rect 2832 4672 2838 4684
rect 3234 4672 3240 4684
rect 2832 4644 3240 4672
rect 2832 4632 2838 4644
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 4338 4681 4344 4684
rect 4332 4672 4344 4681
rect 4251 4644 4344 4672
rect 4332 4635 4344 4644
rect 4396 4672 4402 4684
rect 9692 4681 9720 4712
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 11808 4749 11836 4780
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 13081 4811 13139 4817
rect 13081 4777 13093 4811
rect 13127 4808 13139 4811
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13127 4780 13645 4808
rect 13127 4777 13139 4780
rect 13081 4771 13139 4777
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 14274 4808 14280 4820
rect 14047 4780 14280 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 14274 4768 14280 4780
rect 14332 4808 14338 4820
rect 15010 4808 15016 4820
rect 14332 4780 15016 4808
rect 14332 4768 14338 4780
rect 15010 4768 15016 4780
rect 15068 4768 15074 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4777 15347 4811
rect 15654 4808 15660 4820
rect 15615 4780 15660 4808
rect 15289 4771 15347 4777
rect 11793 4743 11851 4749
rect 11793 4709 11805 4743
rect 11839 4709 11851 4743
rect 11793 4703 11851 4709
rect 12253 4743 12311 4749
rect 12253 4709 12265 4743
rect 12299 4740 12311 4743
rect 12989 4743 13047 4749
rect 12299 4712 12940 4740
rect 12299 4709 12311 4712
rect 12253 4703 12311 4709
rect 7101 4675 7159 4681
rect 4396 4644 6224 4672
rect 4338 4632 4344 4635
rect 4396 4632 4402 4644
rect 6196 4616 6224 4644
rect 7101 4641 7113 4675
rect 7147 4672 7159 4675
rect 9677 4675 9735 4681
rect 7147 4644 7420 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 1394 4564 1400 4616
rect 1452 4604 1458 4616
rect 1946 4604 1952 4616
rect 1452 4576 1952 4604
rect 1452 4564 1458 4576
rect 1946 4564 1952 4576
rect 2004 4604 2010 4616
rect 2041 4607 2099 4613
rect 2041 4604 2053 4607
rect 2004 4576 2053 4604
rect 2004 4564 2010 4576
rect 2041 4573 2053 4576
rect 2087 4573 2099 4607
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 2041 4567 2099 4573
rect 3068 4576 4077 4604
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 2056 4468 2084 4567
rect 3068 4468 3096 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6365 4607 6423 4613
rect 6365 4604 6377 4607
rect 6236 4576 6377 4604
rect 6236 4564 6242 4576
rect 6365 4573 6377 4576
rect 6411 4604 6423 4607
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 6411 4576 7297 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 7285 4573 7297 4576
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 5074 4496 5080 4548
rect 5132 4536 5138 4548
rect 7392 4536 7420 4644
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 9944 4675 10002 4681
rect 9944 4641 9956 4675
rect 9990 4672 10002 4675
rect 10870 4672 10876 4684
rect 9990 4644 10876 4672
rect 9990 4641 10002 4644
rect 9944 4635 10002 4641
rect 10870 4632 10876 4644
rect 10928 4672 10934 4684
rect 10928 4644 11928 4672
rect 10928 4632 10934 4644
rect 11900 4616 11928 4644
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12032 4644 12541 4672
rect 12032 4632 12038 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12912 4672 12940 4712
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 13446 4740 13452 4752
rect 13035 4712 13452 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 13446 4700 13452 4712
rect 13504 4700 13510 4752
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 14093 4743 14151 4749
rect 14093 4740 14105 4743
rect 13872 4712 14105 4740
rect 13872 4700 13878 4712
rect 14093 4709 14105 4712
rect 14139 4709 14151 4743
rect 14093 4703 14151 4709
rect 14550 4700 14556 4752
rect 14608 4740 14614 4752
rect 15304 4740 15332 4771
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 15746 4768 15752 4820
rect 15804 4808 15810 4820
rect 15804 4780 15849 4808
rect 15804 4768 15810 4780
rect 16574 4740 16580 4752
rect 14608 4712 15332 4740
rect 15580 4712 16580 4740
rect 14608 4700 14614 4712
rect 15580 4672 15608 4712
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 17862 4672 17868 4684
rect 12912 4644 15608 4672
rect 17823 4644 17868 4672
rect 12529 4635 12587 4641
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 7834 4604 7840 4616
rect 7795 4576 7840 4604
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 11698 4604 11704 4616
rect 10704 4576 11704 4604
rect 5132 4508 7420 4536
rect 5132 4496 5138 4508
rect 2056 4440 3096 4468
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 3602 4468 3608 4480
rect 3467 4440 3608 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 5442 4468 5448 4480
rect 5403 4440 5448 4468
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5718 4468 5724 4480
rect 5679 4440 5724 4468
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 7392 4468 7420 4508
rect 9217 4539 9275 4545
rect 9217 4505 9229 4539
rect 9263 4536 9275 4539
rect 9306 4536 9312 4548
rect 9263 4508 9312 4536
rect 9263 4505 9275 4508
rect 9217 4499 9275 4505
rect 9306 4496 9312 4508
rect 9364 4536 9370 4548
rect 9582 4536 9588 4548
rect 9364 4508 9588 4536
rect 9364 4496 9370 4508
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 10704 4468 10732 4576
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11882 4604 11888 4616
rect 11843 4576 11888 4604
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 12253 4607 12311 4613
rect 12253 4604 12265 4607
rect 11992 4576 12265 4604
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 11992 4536 12020 4576
rect 12253 4573 12265 4576
rect 12299 4573 12311 4607
rect 13262 4604 13268 4616
rect 13223 4576 13268 4604
rect 12253 4567 12311 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14458 4604 14464 4616
rect 14323 4576 14464 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16206 4604 16212 4616
rect 15979 4576 16212 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 10836 4508 12020 4536
rect 10836 4496 10842 4508
rect 11054 4468 11060 4480
rect 7392 4440 10732 4468
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11330 4468 11336 4480
rect 11291 4440 11336 4468
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 12158 4428 12164 4480
rect 12216 4468 12222 4480
rect 12345 4471 12403 4477
rect 12345 4468 12357 4471
rect 12216 4440 12357 4468
rect 12216 4428 12222 4440
rect 12345 4437 12357 4440
rect 12391 4468 12403 4471
rect 12434 4468 12440 4480
rect 12391 4440 12440 4468
rect 12391 4437 12403 4440
rect 12345 4431 12403 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 12618 4468 12624 4480
rect 12579 4440 12624 4468
rect 12618 4428 12624 4440
rect 12676 4428 12682 4480
rect 13538 4428 13544 4480
rect 13596 4468 13602 4480
rect 13998 4468 14004 4480
rect 13596 4440 14004 4468
rect 13596 4428 13602 4440
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 17920 4440 18061 4468
rect 17920 4428 17926 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18049 4431 18107 4437
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 3973 4267 4031 4273
rect 3973 4233 3985 4267
rect 4019 4264 4031 4267
rect 4338 4264 4344 4276
rect 4019 4236 4344 4264
rect 4019 4233 4031 4236
rect 3973 4227 4031 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 10410 4264 10416 4276
rect 4580 4236 10416 4264
rect 4580 4224 4586 4236
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 15013 4267 15071 4273
rect 15013 4233 15025 4267
rect 15059 4264 15071 4267
rect 16206 4264 16212 4276
rect 15059 4236 16212 4264
rect 15059 4233 15071 4236
rect 15013 4227 15071 4233
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 10318 4196 10324 4208
rect 4304 4168 10324 4196
rect 4304 4156 4310 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 13630 4196 13636 4208
rect 12544 4168 13216 4196
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2004 4100 2605 4128
rect 2004 4088 2010 4100
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 5442 4128 5448 4140
rect 5403 4100 5448 4128
rect 2593 4091 2651 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 8018 4128 8024 4140
rect 6512 4100 8024 4128
rect 6512 4088 6518 4100
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8294 4128 8300 4140
rect 8255 4100 8300 4128
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 9306 4128 9312 4140
rect 9267 4100 9312 4128
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9456 4100 9965 4128
rect 9456 4088 9462 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 12544 4128 12572 4168
rect 9953 4091 10011 4097
rect 12176 4100 12572 4128
rect 12176 4072 12204 4100
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 12676 4100 13093 4128
rect 12676 4088 12682 4100
rect 13081 4097 13093 4100
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 1578 4060 1584 4072
rect 1539 4032 1584 4060
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4060 4307 4063
rect 5261 4063 5319 4069
rect 4295 4032 4568 4060
rect 4295 4029 4307 4032
rect 4249 4023 4307 4029
rect 1210 3952 1216 4004
rect 1268 3992 1274 4004
rect 2866 4001 2872 4004
rect 1857 3995 1915 4001
rect 1857 3992 1869 3995
rect 1268 3964 1869 3992
rect 1268 3952 1274 3964
rect 1857 3961 1869 3964
rect 1903 3961 1915 3995
rect 2860 3992 2872 4001
rect 2827 3964 2872 3992
rect 1857 3955 1915 3961
rect 2860 3955 2872 3964
rect 2866 3952 2872 3955
rect 2924 3952 2930 4004
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 4540 3992 4568 4032
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5718 4060 5724 4072
rect 5307 4032 5724 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 5902 4060 5908 4072
rect 5863 4032 5908 4060
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6420 4032 6837 4060
rect 6420 4020 6426 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 7984 4032 8217 4060
rect 7984 4020 7990 4032
rect 8205 4029 8217 4032
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4060 10747 4063
rect 12158 4060 12164 4072
rect 10735 4032 12164 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 5626 3992 5632 4004
rect 3568 3964 4476 3992
rect 4540 3964 5632 3992
rect 3568 3952 3574 3964
rect 4448 3933 4476 3964
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 5810 3952 5816 4004
rect 5868 3992 5874 4004
rect 6181 3995 6239 4001
rect 6181 3992 6193 3995
rect 5868 3964 6193 3992
rect 5868 3952 5874 3964
rect 6181 3961 6193 3964
rect 6227 3961 6239 3995
rect 6181 3955 6239 3961
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 7101 3995 7159 4001
rect 7101 3992 7113 3995
rect 6696 3964 7113 3992
rect 6696 3952 6702 3964
rect 7101 3961 7113 3964
rect 7147 3961 7159 3995
rect 9125 3995 9183 4001
rect 9125 3992 9137 3995
rect 7101 3955 7159 3961
rect 7944 3964 9137 3992
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 4893 3927 4951 3933
rect 4893 3924 4905 3927
rect 4672 3896 4905 3924
rect 4672 3884 4678 3896
rect 4893 3893 4905 3896
rect 4939 3893 4951 3927
rect 4893 3887 4951 3893
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 6730 3924 6736 3936
rect 5399 3896 6736 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 7944 3924 7972 3964
rect 9125 3961 9137 3964
rect 9171 3961 9183 3995
rect 9125 3955 9183 3961
rect 7791 3896 7972 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8113 3927 8171 3933
rect 8113 3924 8125 3927
rect 8076 3896 8125 3924
rect 8076 3884 8082 3896
rect 8113 3893 8125 3896
rect 8159 3893 8171 3927
rect 8113 3887 8171 3893
rect 8662 3884 8668 3936
rect 8720 3924 8726 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 8720 3896 8769 3924
rect 8720 3884 8726 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 9214 3924 9220 3936
rect 9175 3896 9220 3924
rect 8757 3887 8815 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9784 3924 9812 4023
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12492 4032 12664 4060
rect 12492 4020 12498 4032
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 10934 3995 10992 4001
rect 10934 3992 10946 3995
rect 10652 3964 10946 3992
rect 10652 3952 10658 3964
rect 10934 3961 10946 3964
rect 10980 3961 10992 3995
rect 12636 3992 12664 4032
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12768 4032 13001 4060
rect 12768 4020 12774 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 13188 4060 13216 4168
rect 13280 4168 13636 4196
rect 13280 4137 13308 4168
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 17218 4128 17224 4140
rect 16724 4100 17224 4128
rect 16724 4088 16730 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 13538 4060 13544 4072
rect 13188 4032 13544 4060
rect 12989 4023 13047 4029
rect 13538 4020 13544 4032
rect 13596 4060 13602 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 13596 4032 13645 4060
rect 13596 4020 13602 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 17405 4063 17463 4069
rect 17405 4060 17417 4063
rect 13633 4023 13691 4029
rect 13740 4032 17417 4060
rect 13740 3992 13768 4032
rect 17405 4029 17417 4032
rect 17451 4029 17463 4063
rect 17405 4023 17463 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 13906 4001 13912 4004
rect 13900 3992 13912 4001
rect 10934 3955 10992 3961
rect 11072 3964 12572 3992
rect 12636 3964 13768 3992
rect 13867 3964 13912 3992
rect 11072 3924 11100 3964
rect 12544 3936 12572 3964
rect 13900 3955 13912 3964
rect 13906 3952 13912 3955
rect 13964 3952 13970 4004
rect 13998 3952 14004 4004
rect 14056 3992 14062 4004
rect 18064 3992 18092 4023
rect 14056 3964 18092 3992
rect 14056 3952 14062 3964
rect 12066 3924 12072 3936
rect 9784 3896 11100 3924
rect 12027 3896 12072 3924
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 12526 3884 12532 3936
rect 12584 3884 12590 3936
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 14642 3924 14648 3936
rect 12667 3896 14648 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 17586 3924 17592 3936
rect 17547 3896 17592 3924
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17920 3896 18245 3924
rect 17920 3884 17926 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 1995 3692 3433 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 4614 3720 4620 3732
rect 4575 3692 4620 3720
rect 3421 3683 3479 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 5215 3692 6837 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 6825 3689 6837 3692
rect 6871 3720 6883 3723
rect 7834 3720 7840 3732
rect 6871 3692 7840 3720
rect 6871 3689 6883 3692
rect 6825 3683 6883 3689
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8570 3720 8576 3732
rect 8531 3692 8576 3720
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 9030 3720 9036 3732
rect 8991 3692 9036 3720
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 9677 3723 9735 3729
rect 9677 3720 9689 3723
rect 9640 3692 9689 3720
rect 9640 3680 9646 3692
rect 9677 3689 9689 3692
rect 9723 3689 9735 3723
rect 9677 3683 9735 3689
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 9916 3692 10057 3720
rect 9916 3680 9922 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 10045 3683 10103 3689
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10560 3692 10701 3720
rect 10560 3680 10566 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 10962 3720 10968 3732
rect 10836 3692 10968 3720
rect 10836 3680 10842 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12069 3723 12127 3729
rect 12069 3689 12081 3723
rect 12115 3720 12127 3723
rect 14090 3720 14096 3732
rect 12115 3692 14096 3720
rect 12115 3689 12127 3692
rect 12069 3683 12127 3689
rect 14090 3680 14096 3692
rect 14148 3720 14154 3732
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14148 3692 14289 3720
rect 14148 3680 14154 3692
rect 14277 3689 14289 3692
rect 14323 3720 14335 3723
rect 17770 3720 17776 3732
rect 14323 3692 17776 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 5350 3652 5356 3664
rect 1412 3624 5356 3652
rect 1412 3593 1440 3624
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 5442 3612 5448 3664
rect 5500 3661 5506 3664
rect 5500 3655 5564 3661
rect 5500 3621 5518 3655
rect 5552 3621 5564 3655
rect 8938 3652 8944 3664
rect 8899 3624 8944 3652
rect 5500 3615 5564 3621
rect 5500 3612 5506 3615
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 10137 3655 10195 3661
rect 10137 3621 10149 3655
rect 10183 3652 10195 3655
rect 15194 3652 15200 3664
rect 10183 3624 15200 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3584 2375 3587
rect 2498 3584 2504 3596
rect 2363 3556 2504 3584
rect 2363 3553 2375 3556
rect 2317 3547 2375 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 2958 3544 2964 3596
rect 3016 3584 3022 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 3016 3556 3341 3584
rect 3016 3544 3022 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 7173 3587 7231 3593
rect 7173 3584 7185 3587
rect 3329 3547 3387 3553
rect 6656 3556 7185 3584
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 2280 3488 2421 3516
rect 2280 3476 2286 3488
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 4338 3516 4344 3528
rect 3559 3488 4344 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 2608 3448 2636 3479
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4706 3516 4712 3528
rect 4667 3488 4712 3516
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 5215 3488 5273 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 2866 3448 2872 3460
rect 2608 3420 2872 3448
rect 2866 3408 2872 3420
rect 2924 3448 2930 3460
rect 3602 3448 3608 3460
rect 2924 3420 3608 3448
rect 2924 3408 2930 3420
rect 3602 3408 3608 3420
rect 3660 3408 3666 3460
rect 2961 3383 3019 3389
rect 2961 3349 2973 3383
rect 3007 3380 3019 3383
rect 3786 3380 3792 3392
rect 3007 3352 3792 3380
rect 3007 3349 3019 3352
rect 2961 3343 3019 3349
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4908 3380 4936 3479
rect 6656 3389 6684 3556
rect 7173 3553 7185 3556
rect 7219 3553 7231 3587
rect 7173 3547 7231 3553
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 10505 3587 10563 3593
rect 7708 3556 10364 3584
rect 7708 3544 7714 3556
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6871 3488 6929 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8938 3516 8944 3528
rect 8536 3488 8944 3516
rect 8536 3476 8542 3488
rect 8938 3476 8944 3488
rect 8996 3516 9002 3528
rect 9217 3519 9275 3525
rect 8996 3488 9168 3516
rect 8996 3476 9002 3488
rect 9140 3448 9168 3488
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9306 3516 9312 3528
rect 9263 3488 9312 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9548 3488 10241 3516
rect 9548 3476 9554 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10336 3516 10364 3556
rect 10505 3553 10517 3587
rect 10551 3584 10563 3587
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 10551 3556 11069 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 11057 3553 11069 3556
rect 11103 3553 11115 3587
rect 11974 3584 11980 3596
rect 11057 3547 11115 3553
rect 11164 3556 11980 3584
rect 11164 3525 11192 3556
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 12066 3544 12072 3596
rect 12124 3584 12130 3596
rect 12428 3587 12486 3593
rect 12428 3584 12440 3587
rect 12124 3556 12440 3584
rect 12124 3544 12130 3556
rect 12428 3553 12440 3556
rect 12474 3584 12486 3587
rect 13998 3584 14004 3596
rect 12474 3556 14004 3584
rect 12474 3553 12486 3556
rect 12428 3547 12486 3553
rect 13998 3544 14004 3556
rect 14056 3544 14062 3596
rect 14185 3587 14243 3593
rect 14185 3553 14197 3587
rect 14231 3584 14243 3587
rect 14826 3584 14832 3596
rect 14231 3556 14832 3584
rect 14231 3553 14243 3556
rect 14185 3547 14243 3553
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 17788 3593 17816 3680
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 15712 3556 17233 3584
rect 15712 3544 15718 3556
rect 17221 3553 17233 3556
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 17773 3587 17831 3593
rect 17773 3553 17785 3587
rect 17819 3553 17831 3587
rect 17773 3547 17831 3553
rect 11149 3519 11207 3525
rect 11149 3516 11161 3519
rect 10336 3488 11161 3516
rect 10229 3479 10287 3485
rect 11149 3485 11161 3488
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 12158 3516 12164 3528
rect 11296 3488 11341 3516
rect 12119 3488 12164 3516
rect 11296 3476 11302 3488
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 12069 3451 12127 3457
rect 12069 3448 12081 3451
rect 8119 3420 8423 3448
rect 9140 3420 12081 3448
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 4908 3352 6653 3380
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 6641 3343 6699 3349
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 8119 3380 8147 3420
rect 8294 3380 8300 3392
rect 7340 3352 8147 3380
rect 8255 3352 8300 3380
rect 7340 3340 7346 3352
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 8395 3380 8423 3420
rect 12069 3417 12081 3420
rect 12115 3417 12127 3451
rect 12069 3411 12127 3417
rect 13541 3451 13599 3457
rect 13541 3417 13553 3451
rect 13587 3448 13599 3451
rect 13906 3448 13912 3460
rect 13587 3420 13912 3448
rect 13587 3417 13599 3420
rect 13541 3411 13599 3417
rect 13906 3408 13912 3420
rect 13964 3448 13970 3460
rect 14384 3448 14412 3479
rect 13964 3420 14412 3448
rect 13964 3408 13970 3420
rect 14734 3408 14740 3460
rect 14792 3448 14798 3460
rect 18046 3448 18052 3460
rect 14792 3420 18052 3448
rect 14792 3408 14798 3420
rect 18046 3408 18052 3420
rect 18104 3408 18110 3460
rect 10505 3383 10563 3389
rect 10505 3380 10517 3383
rect 8395 3352 10517 3380
rect 10505 3349 10517 3352
rect 10551 3349 10563 3383
rect 10505 3343 10563 3349
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 13630 3380 13636 3392
rect 11204 3352 13636 3380
rect 11204 3340 11210 3352
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13814 3380 13820 3392
rect 13775 3352 13820 3380
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 17402 3380 17408 3392
rect 17363 3352 17408 3380
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17954 3380 17960 3392
rect 17915 3352 17960 3380
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 3050 3176 3056 3188
rect 2731 3148 3056 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4706 3176 4712 3188
rect 4663 3148 4712 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 7466 3176 7472 3188
rect 5408 3148 7472 3176
rect 5408 3136 5414 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 8481 3179 8539 3185
rect 8481 3145 8493 3179
rect 8527 3176 8539 3179
rect 9214 3176 9220 3188
rect 8527 3148 9220 3176
rect 8527 3145 8539 3148
rect 8481 3139 8539 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 11146 3176 11152 3188
rect 9324 3148 11152 3176
rect 382 3068 388 3120
rect 440 3108 446 3120
rect 9324 3108 9352 3148
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 11256 3148 12265 3176
rect 440 3080 9352 3108
rect 10505 3111 10563 3117
rect 440 3068 446 3080
rect 10505 3077 10517 3111
rect 10551 3108 10563 3111
rect 11256 3108 11284 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 12676 3148 13461 3176
rect 12676 3136 12682 3148
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 13449 3139 13507 3145
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 16301 3179 16359 3185
rect 16301 3176 16313 3179
rect 13688 3148 16313 3176
rect 13688 3136 13694 3148
rect 16301 3145 16313 3148
rect 16347 3145 16359 3179
rect 16301 3139 16359 3145
rect 12066 3108 12072 3120
rect 10551 3080 11284 3108
rect 11440 3080 12072 3108
rect 10551 3077 10563 3080
rect 10505 3071 10563 3077
rect 3234 3040 3240 3052
rect 3195 3012 3240 3040
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 5077 3043 5135 3049
rect 5077 3040 5089 3043
rect 3844 3012 5089 3040
rect 3844 3000 3850 3012
rect 5077 3009 5089 3012
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 5442 3040 5448 3052
rect 5307 3012 5448 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 6086 3040 6092 3052
rect 6047 3012 6092 3040
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6178 3000 6184 3052
rect 6236 3040 6242 3052
rect 8021 3043 8079 3049
rect 6236 3012 6281 3040
rect 6236 3000 6242 3012
rect 8021 3009 8033 3043
rect 8067 3040 8079 3043
rect 8110 3040 8116 3052
rect 8067 3012 8116 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8294 3000 8300 3052
rect 8352 3040 8358 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8352 3012 9045 3040
rect 8352 3000 8358 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9824 3012 10057 3040
rect 9824 3000 9830 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 11054 3040 11060 3052
rect 11015 3012 11060 3040
rect 10045 3003 10103 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2972 1639 2975
rect 3881 2975 3939 2981
rect 1627 2944 3740 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 1857 2907 1915 2913
rect 1857 2873 1869 2907
rect 1903 2904 1915 2907
rect 2774 2904 2780 2916
rect 1903 2876 2780 2904
rect 1903 2873 1915 2876
rect 1857 2867 1915 2873
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 3145 2907 3203 2913
rect 3145 2904 3157 2907
rect 2875 2876 3157 2904
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 2875 2836 2903 2876
rect 3145 2873 3157 2876
rect 3191 2873 3203 2907
rect 3145 2867 3203 2873
rect 3050 2836 3056 2848
rect 1544 2808 2903 2836
rect 3011 2808 3056 2836
rect 1544 2796 1550 2808
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 3712 2836 3740 2944
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 4246 2972 4252 2984
rect 3927 2944 4252 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 7193 2975 7251 2981
rect 7193 2972 7205 2975
rect 4908 2944 7205 2972
rect 3786 2864 3792 2916
rect 3844 2904 3850 2916
rect 4157 2907 4215 2913
rect 4157 2904 4169 2907
rect 3844 2876 4169 2904
rect 3844 2864 3850 2876
rect 4157 2873 4169 2876
rect 4203 2873 4215 2907
rect 4157 2867 4215 2873
rect 4908 2836 4936 2944
rect 7193 2941 7205 2944
rect 7239 2972 7251 2975
rect 7239 2944 7328 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 4985 2907 5043 2913
rect 4985 2873 4997 2907
rect 5031 2904 5043 2907
rect 5031 2876 5672 2904
rect 5031 2873 5043 2876
rect 4985 2867 5043 2873
rect 5644 2845 5672 2876
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 7300 2904 7328 2944
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 8996 2944 9041 2972
rect 8996 2932 9002 2944
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9640 2944 9873 2972
rect 9640 2932 9646 2944
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10873 2975 10931 2981
rect 10873 2941 10885 2975
rect 10919 2972 10931 2975
rect 11440 2972 11468 3080
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3108 12495 3111
rect 12483 3080 13952 3108
rect 12483 3077 12495 3080
rect 12437 3071 12495 3077
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13924 3049 13952 3080
rect 13909 3043 13967 3049
rect 13136 3012 13181 3040
rect 13136 3000 13142 3012
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14918 3040 14924 3052
rect 14056 3012 14101 3040
rect 14200 3012 14924 3040
rect 14056 3000 14062 3012
rect 11606 2972 11612 2984
rect 10919 2944 11468 2972
rect 11567 2944 11612 2972
rect 10919 2941 10931 2944
rect 10873 2935 10931 2941
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 14200 2972 14228 3012
rect 14918 3000 14924 3012
rect 14976 3040 14982 3052
rect 14976 3012 17448 3040
rect 14976 3000 14982 3012
rect 12124 2944 14228 2972
rect 12124 2932 12130 2944
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14424 2944 14473 2972
rect 14424 2932 14430 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 15378 2972 15384 2984
rect 15243 2944 15384 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 16117 2975 16175 2981
rect 15519 2944 15608 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 10226 2904 10232 2916
rect 5776 2876 7236 2904
rect 7300 2876 10232 2904
rect 5776 2864 5782 2876
rect 3712 2808 4936 2836
rect 5629 2839 5687 2845
rect 5629 2805 5641 2839
rect 5675 2805 5687 2839
rect 5629 2799 5687 2805
rect 5997 2839 6055 2845
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6270 2836 6276 2848
rect 6043 2808 6276 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6270 2796 6276 2808
rect 6328 2796 6334 2848
rect 7208 2836 7236 2876
rect 10226 2864 10232 2876
rect 10284 2864 10290 2916
rect 10686 2904 10692 2916
rect 10336 2876 10692 2904
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 7208 2808 8861 2836
rect 8849 2805 8861 2808
rect 8895 2805 8907 2839
rect 8849 2799 8907 2805
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 8996 2808 9505 2836
rect 8996 2796 9002 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9493 2799 9551 2805
rect 9953 2839 10011 2845
rect 9953 2805 9965 2839
rect 9999 2836 10011 2839
rect 10336 2836 10364 2876
rect 10686 2864 10692 2876
rect 10744 2864 10750 2916
rect 11885 2907 11943 2913
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 12158 2904 12164 2916
rect 11931 2876 12164 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 12802 2904 12808 2916
rect 12763 2876 12808 2904
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 14737 2907 14795 2913
rect 14737 2873 14749 2907
rect 14783 2904 14795 2907
rect 14826 2904 14832 2916
rect 14783 2876 14832 2904
rect 14783 2873 14795 2876
rect 14737 2867 14795 2873
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 9999 2808 10364 2836
rect 9999 2805 10011 2808
rect 9953 2799 10011 2805
rect 10502 2796 10508 2848
rect 10560 2836 10566 2848
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 10560 2808 10977 2836
rect 10560 2796 10566 2808
rect 10965 2805 10977 2808
rect 11011 2805 11023 2839
rect 10965 2799 11023 2805
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12299 2808 12909 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 13814 2836 13820 2848
rect 13775 2808 13820 2836
rect 12897 2799 12955 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 15580 2836 15608 2944
rect 16117 2941 16129 2975
rect 16163 2972 16175 2975
rect 16666 2972 16672 2984
rect 16163 2944 16672 2972
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 16850 2972 16856 2984
rect 16811 2944 16856 2972
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 17420 2981 17448 3012
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2941 17463 2975
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 17405 2935 17463 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 17034 2836 17040 2848
rect 13964 2808 15608 2836
rect 16995 2808 17040 2836
rect 13964 2796 13970 2808
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 17589 2839 17647 2845
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 17770 2836 17776 2848
rect 17635 2808 17776 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18230 2836 18236 2848
rect 18191 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 1670 2632 1676 2644
rect 1631 2604 1676 2632
rect 1670 2592 1676 2604
rect 1728 2592 1734 2644
rect 2958 2632 2964 2644
rect 2919 2604 2964 2632
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 4430 2632 4436 2644
rect 4111 2604 4436 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 4982 2632 4988 2644
rect 4943 2604 4988 2632
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 5132 2604 6469 2632
rect 5132 2592 5138 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 8938 2632 8944 2644
rect 6963 2604 8944 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 11333 2635 11391 2641
rect 11333 2632 11345 2635
rect 9171 2604 11345 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 11333 2601 11345 2604
rect 11379 2601 11391 2635
rect 11790 2632 11796 2644
rect 11751 2604 11796 2632
rect 11333 2595 11391 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 16298 2632 16304 2644
rect 11992 2604 16304 2632
rect 4522 2564 4528 2576
rect 1504 2536 4528 2564
rect 1504 2505 1532 2536
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 4890 2564 4896 2576
rect 4851 2536 4896 2564
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 7558 2564 7564 2576
rect 6288 2536 7564 2564
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2465 1547 2499
rect 2038 2496 2044 2508
rect 1999 2468 2044 2496
rect 1489 2459 1547 2465
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 3326 2496 3332 2508
rect 3287 2468 3332 2496
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6288 2505 6316 2536
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 11238 2564 11244 2576
rect 9048 2536 11244 2564
rect 6273 2499 6331 2505
rect 6273 2465 6285 2499
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 6963 2468 7021 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7742 2496 7748 2508
rect 7703 2468 7748 2496
rect 7009 2459 7067 2465
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 9048 2505 9076 2536
rect 11238 2524 11244 2536
rect 11296 2524 11302 2576
rect 11698 2564 11704 2576
rect 11611 2536 11704 2564
rect 11698 2524 11704 2536
rect 11756 2564 11762 2576
rect 11992 2564 12020 2604
rect 16298 2592 16304 2604
rect 16356 2592 16362 2644
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 11756 2536 12020 2564
rect 12084 2536 14933 2564
rect 11756 2524 11762 2536
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2465 9091 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 9033 2459 9091 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 10686 2496 10692 2508
rect 10647 2468 10692 2496
rect 10686 2456 10692 2468
rect 10744 2456 10750 2508
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 12084 2496 12112 2536
rect 14921 2533 14933 2536
rect 14967 2533 14979 2567
rect 14921 2527 14979 2533
rect 10928 2468 12112 2496
rect 10928 2456 10934 2468
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12308 2468 13185 2496
rect 12308 2456 12314 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2496 13967 2499
rect 14182 2496 14188 2508
rect 13955 2468 14188 2496
rect 13955 2465 13967 2468
rect 13909 2459 13967 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 14642 2496 14648 2508
rect 14603 2468 14648 2496
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 15010 2456 15016 2508
rect 15068 2496 15074 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 15068 2468 17141 2496
rect 15068 2456 15074 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17678 2496 17684 2508
rect 17639 2468 17684 2496
rect 17129 2459 17187 2465
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 2130 2388 2136 2440
rect 2188 2428 2194 2440
rect 2225 2431 2283 2437
rect 2225 2428 2237 2431
rect 2188 2400 2237 2428
rect 2188 2388 2194 2400
rect 2225 2397 2237 2400
rect 2271 2397 2283 2431
rect 3602 2428 3608 2440
rect 3515 2400 3608 2428
rect 2225 2391 2283 2397
rect 3602 2388 3608 2400
rect 3660 2428 3666 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 3660 2400 5089 2428
rect 3660 2388 3666 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 4890 2320 4896 2372
rect 4948 2360 4954 2372
rect 5736 2360 5764 2391
rect 4948 2332 5764 2360
rect 7300 2360 7328 2391
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7616 2400 7941 2428
rect 7616 2388 7622 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 10594 2428 10600 2440
rect 9355 2400 10600 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10778 2428 10784 2440
rect 10691 2400 10784 2428
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 10962 2428 10968 2440
rect 10923 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2428 11026 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11020 2400 11897 2428
rect 11020 2388 11026 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 13136 2400 13369 2428
rect 13136 2388 13142 2400
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 8478 2360 8484 2372
rect 7300 2332 8484 2360
rect 4948 2320 4954 2332
rect 8478 2320 8484 2332
rect 8536 2320 8542 2372
rect 8570 2320 8576 2372
rect 8628 2360 8634 2372
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 8628 2332 9965 2360
rect 8628 2320 8634 2332
rect 9953 2329 9965 2332
rect 9999 2329 10011 2363
rect 10796 2360 10824 2388
rect 9953 2323 10011 2329
rect 10244 2332 10824 2360
rect 4525 2295 4583 2301
rect 4525 2261 4537 2295
rect 4571 2292 4583 2295
rect 6086 2292 6092 2304
rect 4571 2264 6092 2292
rect 4571 2261 4583 2264
rect 4525 2255 4583 2261
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 8662 2292 8668 2304
rect 8623 2264 8668 2292
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 9766 2252 9772 2304
rect 9824 2292 9830 2304
rect 10244 2292 10272 2332
rect 11238 2320 11244 2372
rect 11296 2360 11302 2372
rect 14108 2360 14136 2391
rect 11296 2332 14136 2360
rect 11296 2320 11302 2332
rect 9824 2264 10272 2292
rect 10321 2295 10379 2301
rect 9824 2252 9830 2264
rect 10321 2261 10333 2295
rect 10367 2292 10379 2295
rect 12342 2292 12348 2304
rect 10367 2264 12348 2292
rect 10367 2261 10379 2264
rect 10321 2255 10379 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 17310 2292 17316 2304
rect 17271 2264 17316 2292
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17862 2292 17868 2304
rect 17823 2264 17868 2292
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 3326 2048 3332 2100
rect 3384 2088 3390 2100
rect 9766 2088 9772 2100
rect 3384 2060 9772 2088
rect 3384 2048 3390 2060
rect 9766 2048 9772 2060
rect 9824 2048 9830 2100
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 13354 2088 13360 2100
rect 10744 2060 13360 2088
rect 10744 2048 10750 2060
rect 13354 2048 13360 2060
rect 13412 2048 13418 2100
rect 8662 1980 8668 2032
rect 8720 2020 8726 2032
rect 13814 2020 13820 2032
rect 8720 1992 13820 2020
rect 8720 1980 8726 1992
rect 13814 1980 13820 1992
rect 13872 1980 13878 2032
rect 3234 1844 3240 1896
rect 3292 1884 3298 1896
rect 5166 1884 5172 1896
rect 3292 1856 5172 1884
rect 3292 1844 3298 1856
rect 5166 1844 5172 1856
rect 5224 1844 5230 1896
rect 10226 1436 10232 1488
rect 10284 1476 10290 1488
rect 19426 1476 19432 1488
rect 10284 1448 19432 1476
rect 10284 1436 10290 1448
rect 19426 1436 19432 1448
rect 19484 1436 19490 1488
<< via1 >>
rect 4068 15376 4120 15428
rect 5080 15376 5132 15428
rect 3700 15172 3752 15224
rect 5908 15172 5960 15224
rect 3792 14832 3844 14884
rect 10876 14832 10928 14884
rect 9404 14764 9456 14816
rect 17868 14764 17920 14816
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 2044 14424 2096 14476
rect 3056 14424 3108 14476
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 2688 14356 2740 14408
rect 3424 14399 3476 14408
rect 3424 14365 3433 14399
rect 3433 14365 3467 14399
rect 3467 14365 3476 14399
rect 3424 14356 3476 14365
rect 3700 14492 3752 14544
rect 10324 14492 10376 14544
rect 14372 14492 14424 14544
rect 18788 14492 18840 14544
rect 4712 14424 4764 14476
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 17592 14467 17644 14476
rect 17592 14433 17601 14467
rect 17601 14433 17635 14467
rect 17635 14433 17644 14467
rect 17592 14424 17644 14433
rect 5172 14399 5224 14408
rect 5172 14365 5181 14399
rect 5181 14365 5215 14399
rect 5215 14365 5224 14399
rect 5172 14356 5224 14365
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 5264 14356 5316 14365
rect 9956 14356 10008 14408
rect 13360 14356 13412 14408
rect 15108 14356 15160 14408
rect 15568 14356 15620 14408
rect 16120 14356 16172 14408
rect 17316 14356 17368 14408
rect 3332 14288 3384 14340
rect 18052 14288 18104 14340
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 2872 14220 2924 14272
rect 4252 14220 4304 14272
rect 8116 14220 8168 14272
rect 10784 14220 10836 14272
rect 10876 14220 10928 14272
rect 15108 14220 15160 14272
rect 15200 14220 15252 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 2044 14059 2096 14068
rect 2044 14025 2053 14059
rect 2053 14025 2087 14059
rect 2087 14025 2096 14059
rect 2044 14016 2096 14025
rect 2504 13880 2556 13932
rect 3332 14016 3384 14068
rect 3792 14016 3844 14068
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 5356 14016 5408 14068
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 3792 13880 3844 13932
rect 5540 13948 5592 14000
rect 10692 14016 10744 14068
rect 16672 14016 16724 14068
rect 2964 13812 3016 13864
rect 4804 13812 4856 13864
rect 6460 13880 6512 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 14372 13948 14424 14000
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9220 13880 9272 13932
rect 11520 13880 11572 13932
rect 14280 13880 14332 13932
rect 14740 13923 14792 13932
rect 14740 13889 14749 13923
rect 14749 13889 14783 13923
rect 14783 13889 14792 13923
rect 14740 13880 14792 13889
rect 8668 13812 8720 13864
rect 8852 13812 8904 13864
rect 9404 13812 9456 13864
rect 9588 13812 9640 13864
rect 12716 13812 12768 13864
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 15384 13812 15436 13864
rect 18512 13948 18564 14000
rect 16580 13880 16632 13932
rect 17224 13880 17276 13932
rect 17684 13812 17736 13864
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 4252 13744 4304 13796
rect 4712 13744 4764 13796
rect 1400 13676 1452 13728
rect 5632 13676 5684 13728
rect 5816 13744 5868 13796
rect 6736 13744 6788 13796
rect 6092 13719 6144 13728
rect 6092 13685 6101 13719
rect 6101 13685 6135 13719
rect 6135 13685 6144 13719
rect 6092 13676 6144 13685
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 6368 13676 6420 13728
rect 9312 13744 9364 13796
rect 7840 13676 7892 13728
rect 8484 13719 8536 13728
rect 8484 13685 8493 13719
rect 8493 13685 8527 13719
rect 8527 13685 8536 13719
rect 8484 13676 8536 13685
rect 9128 13719 9180 13728
rect 9128 13685 9137 13719
rect 9137 13685 9171 13719
rect 9171 13685 9180 13719
rect 9128 13676 9180 13685
rect 9680 13744 9732 13796
rect 10508 13719 10560 13728
rect 10508 13685 10517 13719
rect 10517 13685 10551 13719
rect 10551 13685 10560 13719
rect 10508 13676 10560 13685
rect 12348 13676 12400 13728
rect 16028 13744 16080 13796
rect 14188 13676 14240 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 2228 13472 2280 13524
rect 2780 13472 2832 13524
rect 3424 13472 3476 13524
rect 5172 13472 5224 13524
rect 6184 13472 6236 13524
rect 6276 13404 6328 13456
rect 6368 13404 6420 13456
rect 1676 13336 1728 13388
rect 2596 13336 2648 13388
rect 3148 13336 3200 13388
rect 5172 13379 5224 13388
rect 5172 13345 5181 13379
rect 5181 13345 5215 13379
rect 5215 13345 5224 13379
rect 5172 13336 5224 13345
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 2780 13268 2832 13320
rect 4896 13268 4948 13320
rect 3700 13200 3752 13252
rect 4712 13200 4764 13252
rect 6000 13268 6052 13320
rect 7472 13472 7524 13524
rect 9128 13472 9180 13524
rect 9312 13472 9364 13524
rect 13268 13472 13320 13524
rect 14188 13515 14240 13524
rect 14188 13481 14197 13515
rect 14197 13481 14231 13515
rect 14231 13481 14240 13515
rect 14188 13472 14240 13481
rect 15384 13472 15436 13524
rect 17592 13472 17644 13524
rect 6736 13404 6788 13456
rect 7748 13404 7800 13456
rect 8116 13404 8168 13456
rect 10140 13404 10192 13456
rect 10324 13447 10376 13456
rect 10324 13413 10333 13447
rect 10333 13413 10367 13447
rect 10367 13413 10376 13447
rect 10324 13404 10376 13413
rect 10692 13404 10744 13456
rect 6644 13268 6696 13320
rect 9036 13311 9088 13320
rect 9036 13277 9045 13311
rect 9045 13277 9079 13311
rect 9079 13277 9088 13311
rect 9036 13268 9088 13277
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9496 13268 9548 13320
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 10876 13336 10928 13388
rect 11612 13336 11664 13388
rect 12164 13404 12216 13456
rect 16028 13404 16080 13456
rect 17776 13447 17828 13456
rect 17776 13413 17785 13447
rect 17785 13413 17819 13447
rect 17819 13413 17828 13447
rect 17776 13404 17828 13413
rect 14004 13336 14056 13388
rect 14464 13336 14516 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 16304 13336 16356 13388
rect 16580 13336 16632 13388
rect 17592 13336 17644 13388
rect 11520 13311 11572 13320
rect 5724 13200 5776 13252
rect 11152 13200 11204 13252
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 14832 13311 14884 13320
rect 14556 13200 14608 13252
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 16212 13268 16264 13320
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 15292 13200 15344 13252
rect 16304 13200 16356 13252
rect 17592 13200 17644 13252
rect 2228 13132 2280 13184
rect 4620 13132 4672 13184
rect 6460 13132 6512 13184
rect 8208 13132 8260 13184
rect 8300 13132 8352 13184
rect 9772 13132 9824 13184
rect 10232 13132 10284 13184
rect 16488 13132 16540 13184
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 3056 12928 3108 12980
rect 3792 12928 3844 12980
rect 10416 12928 10468 12980
rect 4620 12860 4672 12912
rect 6460 12860 6512 12912
rect 8208 12903 8260 12912
rect 8208 12869 8217 12903
rect 8217 12869 8251 12903
rect 8251 12869 8260 12903
rect 8208 12860 8260 12869
rect 9496 12860 9548 12912
rect 14556 12928 14608 12980
rect 14832 12928 14884 12980
rect 16304 12971 16356 12980
rect 16304 12937 16313 12971
rect 16313 12937 16347 12971
rect 16347 12937 16356 12971
rect 16304 12928 16356 12937
rect 16580 12971 16632 12980
rect 16580 12937 16589 12971
rect 16589 12937 16623 12971
rect 16623 12937 16632 12971
rect 16580 12928 16632 12937
rect 13452 12860 13504 12912
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 5448 12792 5500 12844
rect 5724 12792 5776 12844
rect 10784 12835 10836 12844
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 3700 12724 3752 12776
rect 5356 12724 5408 12776
rect 3608 12656 3660 12708
rect 2320 12631 2372 12640
rect 2320 12597 2329 12631
rect 2329 12597 2363 12631
rect 2363 12597 2372 12631
rect 4712 12631 4764 12640
rect 2320 12588 2372 12597
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 5264 12588 5316 12640
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 15936 12792 15988 12844
rect 16212 12792 16264 12844
rect 17776 12792 17828 12844
rect 6644 12724 6696 12776
rect 9220 12724 9272 12776
rect 5816 12588 5868 12640
rect 7472 12656 7524 12708
rect 10968 12724 11020 12776
rect 10324 12656 10376 12708
rect 8392 12588 8444 12640
rect 9128 12588 9180 12640
rect 10232 12588 10284 12640
rect 10416 12588 10468 12640
rect 12348 12724 12400 12776
rect 12532 12724 12584 12776
rect 14648 12724 14700 12776
rect 14740 12724 14792 12776
rect 11428 12656 11480 12708
rect 14280 12656 14332 12708
rect 16856 12656 16908 12708
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 2320 12384 2372 12436
rect 2964 12427 3016 12436
rect 2964 12393 2973 12427
rect 2973 12393 3007 12427
rect 3007 12393 3016 12427
rect 2964 12384 3016 12393
rect 4712 12384 4764 12436
rect 5264 12384 5316 12436
rect 5632 12384 5684 12436
rect 6460 12384 6512 12436
rect 4160 12316 4212 12368
rect 5356 12316 5408 12368
rect 5908 12316 5960 12368
rect 6092 12316 6144 12368
rect 9036 12384 9088 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 2504 12248 2556 12300
rect 5540 12248 5592 12300
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3608 12223 3660 12232
rect 3608 12189 3617 12223
rect 3617 12189 3651 12223
rect 3651 12189 3660 12223
rect 3608 12180 3660 12189
rect 3700 12180 3752 12232
rect 3424 12044 3476 12096
rect 6184 12044 6236 12096
rect 7656 12316 7708 12368
rect 9772 12316 9824 12368
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 7288 12180 7340 12232
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 8392 12180 8444 12232
rect 9036 12223 9088 12232
rect 9036 12189 9045 12223
rect 9045 12189 9079 12223
rect 9079 12189 9088 12223
rect 9036 12180 9088 12189
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 10600 12384 10652 12436
rect 10784 12316 10836 12368
rect 11980 12316 12032 12368
rect 14464 12384 14516 12436
rect 14648 12427 14700 12436
rect 14648 12393 14657 12427
rect 14657 12393 14691 12427
rect 14691 12393 14700 12427
rect 14648 12384 14700 12393
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 14740 12316 14792 12368
rect 15752 12316 15804 12368
rect 16304 12316 16356 12368
rect 9220 12180 9272 12189
rect 12164 12248 12216 12300
rect 14096 12248 14148 12300
rect 14280 12248 14332 12300
rect 14556 12248 14608 12300
rect 12716 12223 12768 12232
rect 7380 12044 7432 12096
rect 8024 12044 8076 12096
rect 9312 12044 9364 12096
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 10416 12044 10468 12096
rect 11704 12044 11756 12096
rect 13176 12180 13228 12232
rect 15844 12248 15896 12300
rect 16488 12248 16540 12300
rect 16948 12248 17000 12300
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 15292 12112 15344 12164
rect 13912 12044 13964 12096
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 2780 11840 2832 11892
rect 6460 11840 6512 11892
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 9496 11840 9548 11892
rect 11612 11840 11664 11892
rect 12716 11840 12768 11892
rect 3148 11772 3200 11824
rect 4712 11772 4764 11824
rect 7472 11772 7524 11824
rect 13728 11840 13780 11892
rect 14096 11883 14148 11892
rect 14096 11849 14105 11883
rect 14105 11849 14139 11883
rect 14139 11849 14148 11883
rect 14096 11840 14148 11849
rect 14464 11840 14516 11892
rect 2596 11704 2648 11756
rect 9220 11704 9272 11756
rect 13360 11772 13412 11824
rect 15200 11772 15252 11824
rect 13452 11704 13504 11756
rect 13544 11747 13596 11756
rect 13544 11713 13553 11747
rect 13553 11713 13587 11747
rect 13587 11713 13596 11747
rect 13544 11704 13596 11713
rect 13820 11704 13872 11756
rect 3700 11679 3752 11688
rect 3700 11645 3709 11679
rect 3709 11645 3743 11679
rect 3743 11645 3752 11679
rect 3700 11636 3752 11645
rect 3792 11636 3844 11688
rect 4344 11636 4396 11688
rect 6276 11636 6328 11688
rect 7196 11636 7248 11688
rect 3424 11568 3476 11620
rect 4712 11568 4764 11620
rect 8116 11636 8168 11688
rect 10232 11636 10284 11688
rect 10324 11636 10376 11688
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 14464 11679 14516 11688
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 15108 11636 15160 11688
rect 15292 11636 15344 11688
rect 15936 11636 15988 11688
rect 7748 11568 7800 11620
rect 9312 11568 9364 11620
rect 10968 11568 11020 11620
rect 16672 11568 16724 11620
rect 2780 11500 2832 11552
rect 3516 11500 3568 11552
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 5908 11500 5960 11552
rect 6644 11500 6696 11552
rect 7564 11500 7616 11552
rect 8944 11543 8996 11552
rect 8944 11509 8953 11543
rect 8953 11509 8987 11543
rect 8987 11509 8996 11543
rect 8944 11500 8996 11509
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 10600 11500 10652 11552
rect 11060 11500 11112 11552
rect 11612 11500 11664 11552
rect 13176 11500 13228 11552
rect 13268 11500 13320 11552
rect 13728 11500 13780 11552
rect 16948 11500 17000 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2964 11296 3016 11348
rect 3424 11296 3476 11348
rect 3884 11296 3936 11348
rect 5632 11296 5684 11348
rect 7748 11296 7800 11348
rect 7840 11296 7892 11348
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 3700 11228 3752 11280
rect 2320 11203 2372 11212
rect 2320 11169 2354 11203
rect 2354 11169 2372 11203
rect 2320 11160 2372 11169
rect 5080 11160 5132 11212
rect 3792 11092 3844 11144
rect 7472 11228 7524 11280
rect 8300 11228 8352 11280
rect 9772 11296 9824 11348
rect 13360 11296 13412 11348
rect 13452 11296 13504 11348
rect 14464 11339 14516 11348
rect 14464 11305 14473 11339
rect 14473 11305 14507 11339
rect 14507 11305 14516 11339
rect 14464 11296 14516 11305
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 16764 11296 16816 11348
rect 11152 11228 11204 11280
rect 13820 11228 13872 11280
rect 16212 11228 16264 11280
rect 8024 11203 8076 11212
rect 5724 11092 5776 11144
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 2688 10956 2740 11008
rect 6368 11067 6420 11076
rect 6368 11033 6377 11067
rect 6377 11033 6411 11067
rect 6411 11033 6420 11067
rect 6368 11024 6420 11033
rect 7748 11024 7800 11076
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 7932 11092 7984 11144
rect 8668 11160 8720 11212
rect 10140 11160 10192 11212
rect 10232 11160 10284 11212
rect 8024 11024 8076 11076
rect 9772 11092 9824 11144
rect 10968 11092 11020 11144
rect 8944 11024 8996 11076
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 10232 11024 10284 11076
rect 10416 11024 10468 11076
rect 13912 11160 13964 11212
rect 14556 11160 14608 11212
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 15292 11135 15344 11144
rect 12808 11092 12860 11101
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 16580 11160 16632 11212
rect 17316 11092 17368 11144
rect 17776 11092 17828 11144
rect 3700 10956 3752 11008
rect 8484 10956 8536 11008
rect 8668 10956 8720 11008
rect 12348 10956 12400 11008
rect 12624 10956 12676 11008
rect 16212 10956 16264 11008
rect 16948 10956 17000 11008
rect 17776 10956 17828 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 3700 10795 3752 10804
rect 3700 10761 3709 10795
rect 3709 10761 3743 10795
rect 3743 10761 3752 10795
rect 3700 10752 3752 10761
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2872 10684 2924 10736
rect 6828 10752 6880 10804
rect 7012 10752 7064 10804
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 3240 10616 3292 10668
rect 4988 10616 5040 10668
rect 1768 10548 1820 10600
rect 3332 10548 3384 10600
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4712 10548 4764 10600
rect 4896 10548 4948 10600
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5356 10616 5408 10668
rect 6644 10616 6696 10668
rect 9772 10752 9824 10804
rect 10784 10752 10836 10804
rect 11060 10752 11112 10804
rect 7840 10548 7892 10600
rect 8024 10548 8076 10600
rect 8300 10548 8352 10600
rect 1584 10412 1636 10464
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 3792 10412 3844 10464
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 5540 10412 5592 10464
rect 6092 10455 6144 10464
rect 6092 10421 6101 10455
rect 6101 10421 6135 10455
rect 6135 10421 6144 10455
rect 6092 10412 6144 10421
rect 6736 10480 6788 10532
rect 7564 10480 7616 10532
rect 9772 10548 9824 10600
rect 10232 10548 10284 10600
rect 12348 10752 12400 10804
rect 16396 10752 16448 10804
rect 17316 10752 17368 10804
rect 12532 10684 12584 10736
rect 8944 10480 8996 10532
rect 12624 10480 12676 10532
rect 9220 10412 9272 10464
rect 10968 10412 11020 10464
rect 12440 10412 12492 10464
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 15108 10548 15160 10600
rect 15292 10548 15344 10600
rect 15476 10548 15528 10600
rect 13452 10480 13504 10532
rect 17592 10548 17644 10600
rect 13728 10412 13780 10464
rect 14648 10455 14700 10464
rect 14648 10421 14657 10455
rect 14657 10421 14691 10455
rect 14691 10421 14700 10455
rect 14648 10412 14700 10421
rect 15292 10412 15344 10464
rect 16212 10412 16264 10464
rect 16580 10412 16632 10464
rect 16764 10412 16816 10464
rect 17316 10412 17368 10464
rect 17592 10412 17644 10464
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 2504 10208 2556 10260
rect 3608 10208 3660 10260
rect 5448 10208 5500 10260
rect 11244 10208 11296 10260
rect 2688 10140 2740 10192
rect 6644 10140 6696 10192
rect 7012 10140 7064 10192
rect 7472 10140 7524 10192
rect 9496 10140 9548 10192
rect 12532 10140 12584 10192
rect 17040 10208 17092 10260
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3792 10072 3844 10124
rect 7196 10072 7248 10124
rect 7656 10072 7708 10124
rect 8208 10072 8260 10124
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9036 10072 9088 10124
rect 9404 10072 9456 10124
rect 9772 10072 9824 10124
rect 10968 10072 11020 10124
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5356 10004 5408 10056
rect 5448 9936 5500 9988
rect 6736 9936 6788 9988
rect 11980 10004 12032 10056
rect 12716 10004 12768 10056
rect 13636 10140 13688 10192
rect 16396 10140 16448 10192
rect 13728 10072 13780 10124
rect 13636 10004 13688 10056
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 13176 9936 13228 9988
rect 14096 9936 14148 9988
rect 17316 10072 17368 10124
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 17040 10004 17092 10056
rect 17776 10047 17828 10056
rect 16948 9936 17000 9988
rect 17776 10013 17785 10047
rect 17785 10013 17819 10047
rect 17819 10013 17828 10047
rect 17776 10004 17828 10013
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 4988 9868 5040 9920
rect 7472 9868 7524 9920
rect 8300 9868 8352 9920
rect 8668 9868 8720 9920
rect 12348 9868 12400 9920
rect 13268 9868 13320 9920
rect 13728 9868 13780 9920
rect 15476 9911 15528 9920
rect 15476 9877 15485 9911
rect 15485 9877 15519 9911
rect 15519 9877 15528 9911
rect 15476 9868 15528 9877
rect 16764 9868 16816 9920
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 1400 9664 1452 9716
rect 3792 9664 3844 9716
rect 5080 9664 5132 9716
rect 7564 9664 7616 9716
rect 8668 9664 8720 9716
rect 9220 9664 9272 9716
rect 3516 9596 3568 9648
rect 5172 9596 5224 9648
rect 5724 9639 5776 9648
rect 5724 9605 5733 9639
rect 5733 9605 5767 9639
rect 5767 9605 5776 9639
rect 5724 9596 5776 9605
rect 6184 9596 6236 9648
rect 8944 9596 8996 9648
rect 9588 9596 9640 9648
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 4344 9528 4396 9580
rect 4804 9528 4856 9580
rect 11244 9664 11296 9716
rect 13636 9664 13688 9716
rect 14004 9664 14056 9716
rect 14280 9664 14332 9716
rect 14464 9664 14516 9716
rect 16212 9664 16264 9716
rect 16948 9664 17000 9716
rect 17960 9664 18012 9716
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6736 9528 6788 9580
rect 7196 9528 7248 9580
rect 8208 9528 8260 9580
rect 8484 9528 8536 9580
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11152 9528 11204 9580
rect 1952 9392 2004 9444
rect 4528 9460 4580 9512
rect 4620 9460 4672 9512
rect 5172 9460 5224 9512
rect 8116 9460 8168 9512
rect 8576 9460 8628 9512
rect 9220 9460 9272 9512
rect 2504 9392 2556 9444
rect 2688 9392 2740 9444
rect 5724 9392 5776 9444
rect 7564 9392 7616 9444
rect 9312 9392 9364 9444
rect 9772 9392 9824 9444
rect 12348 9460 12400 9512
rect 13544 9596 13596 9648
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 15844 9596 15896 9648
rect 17408 9596 17460 9648
rect 17776 9596 17828 9648
rect 15476 9528 15528 9580
rect 16028 9528 16080 9580
rect 13820 9460 13872 9512
rect 14648 9460 14700 9512
rect 15108 9460 15160 9512
rect 15384 9460 15436 9512
rect 12716 9435 12768 9444
rect 12716 9401 12750 9435
rect 12750 9401 12768 9435
rect 12716 9392 12768 9401
rect 17408 9392 17460 9444
rect 3516 9324 3568 9376
rect 4068 9324 4120 9376
rect 4344 9324 4396 9376
rect 4804 9324 4856 9376
rect 5632 9324 5684 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 6460 9324 6512 9376
rect 6736 9324 6788 9376
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 10324 9324 10376 9376
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 12532 9324 12584 9376
rect 12624 9324 12676 9376
rect 14464 9324 14516 9376
rect 14648 9324 14700 9376
rect 17040 9324 17092 9376
rect 17960 9324 18012 9376
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 4436 9120 4488 9172
rect 7288 9120 7340 9172
rect 8208 9120 8260 9172
rect 10508 9120 10560 9172
rect 11704 9120 11756 9172
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 12532 9120 12584 9172
rect 13268 9120 13320 9172
rect 14004 9120 14056 9172
rect 16488 9120 16540 9172
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 2780 8848 2832 8900
rect 3332 9027 3384 9036
rect 3332 8993 3341 9027
rect 3341 8993 3375 9027
rect 3375 8993 3384 9027
rect 4068 9052 4120 9104
rect 4252 9052 4304 9104
rect 6276 9052 6328 9104
rect 6736 9052 6788 9104
rect 3332 8984 3384 8993
rect 5540 8984 5592 9036
rect 6552 8984 6604 9036
rect 10416 8984 10468 9036
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3332 8848 3384 8900
rect 2412 8780 2464 8832
rect 3792 8916 3844 8968
rect 6736 8916 6788 8968
rect 4712 8780 4764 8832
rect 5724 8780 5776 8832
rect 7104 8780 7156 8832
rect 7564 8780 7616 8832
rect 8024 8780 8076 8832
rect 8116 8780 8168 8832
rect 10968 8916 11020 8968
rect 10968 8780 11020 8832
rect 14096 8984 14148 9036
rect 14556 9027 14608 9036
rect 14556 8993 14565 9027
rect 14565 8993 14599 9027
rect 14599 8993 14608 9027
rect 14556 8984 14608 8993
rect 16672 9052 16724 9104
rect 16304 9027 16356 9036
rect 16304 8993 16327 9027
rect 16327 8993 16356 9027
rect 16304 8984 16356 8993
rect 17776 8984 17828 9036
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 14464 8916 14516 8968
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 16028 8959 16080 8968
rect 14740 8916 14792 8925
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 12992 8848 13044 8900
rect 14556 8780 14608 8832
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 16212 8780 16264 8832
rect 17408 8823 17460 8832
rect 17408 8789 17417 8823
rect 17417 8789 17451 8823
rect 17451 8789 17460 8823
rect 17408 8780 17460 8789
rect 17868 8780 17920 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 3424 8576 3476 8628
rect 3792 8576 3844 8628
rect 2596 8508 2648 8560
rect 5264 8576 5316 8628
rect 6184 8576 6236 8628
rect 7656 8576 7708 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 6276 8508 6328 8560
rect 2872 8440 2924 8492
rect 3424 8440 3476 8492
rect 3608 8440 3660 8492
rect 4252 8440 4304 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 4620 8372 4672 8424
rect 11520 8508 11572 8560
rect 8208 8440 8260 8492
rect 14188 8508 14240 8560
rect 16212 8508 16264 8560
rect 2504 8304 2556 8356
rect 6644 8372 6696 8424
rect 5264 8347 5316 8356
rect 2872 8236 2924 8288
rect 4068 8236 4120 8288
rect 5264 8313 5298 8347
rect 5298 8313 5316 8347
rect 5264 8304 5316 8313
rect 6920 8304 6972 8356
rect 7380 8304 7432 8356
rect 7840 8372 7892 8424
rect 8116 8304 8168 8356
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12532 8440 12584 8492
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 18236 8551 18288 8560
rect 18236 8517 18245 8551
rect 18245 8517 18279 8551
rect 18279 8517 18288 8551
rect 18236 8508 18288 8517
rect 14648 8440 14700 8449
rect 12072 8304 12124 8356
rect 4528 8279 4580 8288
rect 4528 8245 4537 8279
rect 4537 8245 4571 8279
rect 4571 8245 4580 8279
rect 4528 8236 4580 8245
rect 7472 8236 7524 8288
rect 8392 8236 8444 8288
rect 11152 8236 11204 8288
rect 15016 8372 15068 8424
rect 12440 8304 12492 8356
rect 13728 8304 13780 8356
rect 15200 8372 15252 8424
rect 16488 8372 16540 8424
rect 16304 8304 16356 8356
rect 13452 8236 13504 8288
rect 13544 8236 13596 8288
rect 14740 8236 14792 8288
rect 14832 8236 14884 8288
rect 15292 8236 15344 8288
rect 17040 8304 17092 8356
rect 17132 8279 17184 8288
rect 17132 8245 17141 8279
rect 17141 8245 17175 8279
rect 17175 8245 17184 8279
rect 17132 8236 17184 8245
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 3148 8032 3200 8084
rect 10232 8032 10284 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 2412 8007 2464 8016
rect 2412 7973 2421 8007
rect 2421 7973 2455 8007
rect 2455 7973 2464 8007
rect 2412 7964 2464 7973
rect 3608 7964 3660 8016
rect 1492 7896 1544 7948
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 8576 7964 8628 8016
rect 8668 7964 8720 8016
rect 11796 8032 11848 8084
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 13636 8032 13688 8084
rect 15200 8032 15252 8084
rect 11888 7964 11940 8016
rect 14648 7964 14700 8016
rect 4804 7896 4856 7948
rect 6736 7896 6788 7948
rect 8392 7939 8444 7948
rect 8392 7905 8426 7939
rect 8426 7905 8444 7939
rect 8392 7896 8444 7905
rect 8760 7896 8812 7948
rect 9496 7896 9548 7948
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 13544 7896 13596 7948
rect 16856 8032 16908 8084
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 18328 8032 18380 8084
rect 16672 8007 16724 8016
rect 16672 7973 16681 8007
rect 16681 7973 16715 8007
rect 16715 7973 16724 8007
rect 16672 7964 16724 7973
rect 17776 7964 17828 8016
rect 2872 7828 2924 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7288 7828 7340 7880
rect 7472 7828 7524 7880
rect 9312 7828 9364 7880
rect 2872 7692 2924 7744
rect 3608 7692 3660 7744
rect 8024 7760 8076 7812
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 5080 7735 5132 7744
rect 4896 7692 4948 7701
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 5080 7692 5132 7701
rect 5540 7692 5592 7744
rect 7932 7692 7984 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 9588 7692 9640 7744
rect 10508 7828 10560 7880
rect 15660 7828 15712 7880
rect 17408 7896 17460 7948
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 17132 7760 17184 7812
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 16856 7692 16908 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 4712 7488 4764 7540
rect 5264 7488 5316 7540
rect 9312 7488 9364 7540
rect 9404 7488 9456 7540
rect 11888 7531 11940 7540
rect 1400 7352 1452 7404
rect 4896 7420 4948 7472
rect 6184 7420 6236 7472
rect 8668 7420 8720 7472
rect 2964 7284 3016 7336
rect 4160 7327 4212 7336
rect 4160 7293 4169 7327
rect 4169 7293 4203 7327
rect 4203 7293 4212 7327
rect 4160 7284 4212 7293
rect 6552 7352 6604 7404
rect 7564 7352 7616 7404
rect 8208 7352 8260 7404
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 12256 7420 12308 7472
rect 12716 7488 12768 7540
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 18236 7531 18288 7540
rect 13176 7420 13228 7472
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 15292 7352 15344 7404
rect 16212 7352 16264 7404
rect 16488 7352 16540 7404
rect 4620 7284 4672 7336
rect 4068 7216 4120 7268
rect 7380 7284 7432 7336
rect 8760 7284 8812 7336
rect 12532 7284 12584 7336
rect 5356 7216 5408 7268
rect 8300 7216 8352 7268
rect 13176 7284 13228 7336
rect 13636 7284 13688 7336
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 15660 7284 15712 7336
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 15844 7284 15896 7293
rect 16396 7284 16448 7336
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 3056 7191 3108 7200
rect 3056 7157 3065 7191
rect 3065 7157 3099 7191
rect 3099 7157 3108 7191
rect 3056 7148 3108 7157
rect 3332 7148 3384 7200
rect 6184 7148 6236 7200
rect 6736 7148 6788 7200
rect 8024 7148 8076 7200
rect 9772 7148 9824 7200
rect 11980 7148 12032 7200
rect 13820 7148 13872 7200
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 14740 7148 14792 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 15844 7148 15896 7200
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 4344 6944 4396 6996
rect 4988 6944 5040 6996
rect 5264 6944 5316 6996
rect 6644 6944 6696 6996
rect 8300 6944 8352 6996
rect 9588 6944 9640 6996
rect 3148 6876 3200 6928
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 3056 6808 3108 6860
rect 1400 6740 1452 6792
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 5356 6808 5408 6860
rect 8852 6876 8904 6928
rect 10600 6944 10652 6996
rect 12348 6944 12400 6996
rect 12716 6987 12768 6996
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 13268 6944 13320 6996
rect 14464 6944 14516 6996
rect 15200 6944 15252 6996
rect 16764 6987 16816 6996
rect 16764 6953 16773 6987
rect 16773 6953 16807 6987
rect 16807 6953 16816 6987
rect 16764 6944 16816 6953
rect 18144 6944 18196 6996
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 5816 6740 5868 6792
rect 6000 6740 6052 6792
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 7472 6808 7524 6860
rect 8208 6808 8260 6860
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10508 6876 10560 6928
rect 10968 6876 11020 6928
rect 11980 6876 12032 6928
rect 15568 6876 15620 6928
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 11520 6740 11572 6792
rect 12256 6740 12308 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 14740 6808 14792 6860
rect 16580 6876 16632 6928
rect 13084 6740 13136 6792
rect 13728 6740 13780 6792
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 14464 6740 14516 6792
rect 15108 6740 15160 6792
rect 2964 6604 3016 6656
rect 3792 6604 3844 6656
rect 5172 6604 5224 6656
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 13084 6604 13136 6656
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 16948 6808 17000 6860
rect 17592 6740 17644 6792
rect 17868 6740 17920 6792
rect 17500 6715 17552 6724
rect 17500 6681 17509 6715
rect 17509 6681 17543 6715
rect 17543 6681 17552 6715
rect 17500 6672 17552 6681
rect 15660 6604 15712 6656
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2320 6400 2372 6452
rect 3148 6400 3200 6452
rect 4436 6400 4488 6452
rect 5080 6400 5132 6452
rect 5264 6400 5316 6452
rect 6736 6400 6788 6452
rect 6828 6400 6880 6452
rect 8208 6443 8260 6452
rect 4252 6332 4304 6384
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 8668 6332 8720 6384
rect 2596 6264 2648 6316
rect 2872 6307 2924 6316
rect 2872 6273 2881 6307
rect 2881 6273 2915 6307
rect 2915 6273 2924 6307
rect 2872 6264 2924 6273
rect 3148 6264 3200 6316
rect 3424 6264 3476 6316
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 5172 6264 5224 6316
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 5632 6196 5684 6248
rect 9404 6400 9456 6452
rect 12072 6400 12124 6452
rect 12808 6400 12860 6452
rect 14004 6400 14056 6452
rect 17592 6443 17644 6452
rect 17592 6409 17601 6443
rect 17601 6409 17635 6443
rect 17635 6409 17644 6443
rect 17592 6400 17644 6409
rect 18236 6443 18288 6452
rect 18236 6409 18245 6443
rect 18245 6409 18279 6443
rect 18279 6409 18288 6443
rect 18236 6400 18288 6409
rect 13360 6332 13412 6384
rect 12440 6264 12492 6316
rect 14004 6264 14056 6316
rect 15108 6264 15160 6316
rect 5356 6128 5408 6180
rect 1492 6060 1544 6112
rect 1768 6103 1820 6112
rect 1768 6069 1777 6103
rect 1777 6069 1811 6103
rect 1811 6069 1820 6103
rect 1768 6060 1820 6069
rect 2044 6060 2096 6112
rect 5816 6060 5868 6112
rect 6092 6060 6144 6112
rect 6552 6060 6604 6112
rect 10508 6196 10560 6248
rect 12348 6196 12400 6248
rect 13636 6196 13688 6248
rect 6920 6128 6972 6180
rect 7288 6128 7340 6180
rect 7932 6128 7984 6180
rect 8300 6128 8352 6180
rect 9772 6128 9824 6180
rect 11796 6128 11848 6180
rect 12072 6128 12124 6180
rect 13820 6128 13872 6180
rect 16580 6196 16632 6248
rect 14464 6128 14516 6180
rect 8208 6060 8260 6112
rect 8944 6060 8996 6112
rect 11244 6060 11296 6112
rect 12164 6060 12216 6112
rect 13176 6060 13228 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 13728 6060 13780 6112
rect 15200 6060 15252 6112
rect 17040 6128 17092 6180
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 1768 5856 1820 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 5264 5899 5316 5908
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 7288 5856 7340 5908
rect 7472 5856 7524 5908
rect 11888 5856 11940 5908
rect 12256 5856 12308 5908
rect 13452 5856 13504 5908
rect 14004 5899 14056 5908
rect 1400 5720 1452 5772
rect 3700 5720 3752 5772
rect 5264 5720 5316 5772
rect 4344 5652 4396 5704
rect 4528 5584 4580 5636
rect 2596 5516 2648 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 4896 5516 4948 5568
rect 5264 5516 5316 5568
rect 6552 5720 6604 5772
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 7288 5720 7340 5772
rect 9588 5720 9640 5772
rect 10508 5788 10560 5840
rect 14004 5865 14013 5899
rect 14013 5865 14047 5899
rect 14047 5865 14056 5899
rect 14004 5856 14056 5865
rect 14464 5856 14516 5908
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 11244 5720 11296 5772
rect 13728 5720 13780 5772
rect 16672 5720 16724 5772
rect 7380 5652 7432 5704
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 12440 5652 12492 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 16212 5652 16264 5704
rect 16304 5652 16356 5704
rect 7656 5584 7708 5636
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 8208 5516 8260 5568
rect 11704 5584 11756 5636
rect 12164 5584 12216 5636
rect 17500 5627 17552 5636
rect 17500 5593 17509 5627
rect 17509 5593 17543 5627
rect 17543 5593 17552 5627
rect 17500 5584 17552 5593
rect 11888 5516 11940 5568
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 3700 5312 3752 5364
rect 4252 5312 4304 5364
rect 5172 5312 5224 5364
rect 6276 5312 6328 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 2596 5176 2648 5228
rect 4436 5176 4488 5228
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 6736 5176 6788 5228
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 10232 5312 10284 5364
rect 7472 5244 7524 5296
rect 11428 5244 11480 5296
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 3148 5040 3200 5092
rect 2780 5015 2832 5024
rect 2780 4981 2789 5015
rect 2789 4981 2823 5015
rect 2823 4981 2832 5015
rect 6460 5108 6512 5160
rect 4252 5083 4304 5092
rect 4252 5049 4261 5083
rect 4261 5049 4295 5083
rect 4295 5049 4304 5083
rect 4252 5040 4304 5049
rect 7564 5108 7616 5160
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 2780 4972 2832 4981
rect 4528 4972 4580 5024
rect 6920 5040 6972 5092
rect 5264 5015 5316 5024
rect 5264 4981 5273 5015
rect 5273 4981 5307 5015
rect 5307 4981 5316 5015
rect 5264 4972 5316 4981
rect 5448 4972 5500 5024
rect 6276 4972 6328 5024
rect 6552 4972 6604 5024
rect 8300 4972 8352 5024
rect 8760 5176 8812 5228
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 9588 5176 9640 5228
rect 13728 5312 13780 5364
rect 15476 5244 15528 5296
rect 10784 5108 10836 5160
rect 12440 5151 12492 5160
rect 9404 5040 9456 5092
rect 10232 4972 10284 5024
rect 10324 5015 10376 5024
rect 10324 4981 10333 5015
rect 10333 4981 10367 5015
rect 10367 4981 10376 5015
rect 10876 5015 10928 5024
rect 10324 4972 10376 4981
rect 10876 4981 10885 5015
rect 10885 4981 10919 5015
rect 10919 4981 10928 5015
rect 10876 4972 10928 4981
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 16212 5176 16264 5228
rect 12532 5040 12584 5092
rect 13636 5108 13688 5160
rect 14464 5108 14516 5160
rect 17408 5151 17460 5160
rect 17408 5117 17417 5151
rect 17417 5117 17451 5151
rect 17451 5117 17460 5151
rect 17408 5108 17460 5117
rect 13268 5040 13320 5092
rect 15292 4972 15344 5024
rect 16580 5040 16632 5092
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 17592 4972 17644 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 6276 4768 6328 4820
rect 9036 4768 9088 4820
rect 10600 4768 10652 4820
rect 10876 4768 10928 4820
rect 4252 4700 4304 4752
rect 4436 4700 4488 4752
rect 7472 4700 7524 4752
rect 8300 4700 8352 4752
rect 2780 4632 2832 4684
rect 3240 4632 3292 4684
rect 4344 4675 4396 4684
rect 4344 4641 4378 4675
rect 4378 4641 4396 4675
rect 10508 4700 10560 4752
rect 12072 4768 12124 4820
rect 14280 4768 14332 4820
rect 15016 4768 15068 4820
rect 15660 4811 15712 4820
rect 4344 4632 4396 4641
rect 1400 4564 1452 4616
rect 1952 4564 2004 4616
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 6184 4564 6236 4616
rect 5080 4496 5132 4548
rect 10876 4632 10928 4684
rect 11980 4632 12032 4684
rect 13452 4700 13504 4752
rect 13820 4700 13872 4752
rect 14556 4700 14608 4752
rect 15660 4777 15669 4811
rect 15669 4777 15703 4811
rect 15703 4777 15712 4811
rect 15660 4768 15712 4777
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 16580 4700 16632 4752
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 3608 4428 3660 4480
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 5724 4471 5776 4480
rect 5724 4437 5733 4471
rect 5733 4437 5767 4471
rect 5767 4437 5776 4471
rect 5724 4428 5776 4437
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 9312 4496 9364 4548
rect 9588 4496 9640 4548
rect 11704 4564 11756 4616
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 10784 4496 10836 4548
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 14464 4564 14516 4616
rect 16212 4564 16264 4616
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 12164 4428 12216 4480
rect 12440 4428 12492 4480
rect 12624 4471 12676 4480
rect 12624 4437 12633 4471
rect 12633 4437 12667 4471
rect 12667 4437 12676 4471
rect 12624 4428 12676 4437
rect 13544 4428 13596 4480
rect 14004 4428 14056 4480
rect 17868 4428 17920 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 4344 4224 4396 4276
rect 4528 4224 4580 4276
rect 10416 4224 10468 4276
rect 16212 4224 16264 4276
rect 4252 4156 4304 4208
rect 10324 4156 10376 4208
rect 1952 4088 2004 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 6460 4088 6512 4140
rect 8024 4088 8076 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 9404 4088 9456 4140
rect 12624 4088 12676 4140
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 1216 3952 1268 4004
rect 2872 3995 2924 4004
rect 2872 3961 2906 3995
rect 2906 3961 2924 3995
rect 2872 3952 2924 3961
rect 3516 3952 3568 4004
rect 5724 4020 5776 4072
rect 5908 4063 5960 4072
rect 5908 4029 5917 4063
rect 5917 4029 5951 4063
rect 5951 4029 5960 4063
rect 5908 4020 5960 4029
rect 6368 4020 6420 4072
rect 7932 4020 7984 4072
rect 5632 3952 5684 4004
rect 5816 3952 5868 4004
rect 6644 3952 6696 4004
rect 4620 3884 4672 3936
rect 6736 3884 6788 3936
rect 8024 3884 8076 3936
rect 8668 3884 8720 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 12164 4020 12216 4072
rect 12440 4020 12492 4072
rect 10600 3952 10652 4004
rect 12716 4020 12768 4072
rect 13636 4156 13688 4208
rect 16672 4088 16724 4140
rect 17224 4088 17276 4140
rect 13544 4020 13596 4072
rect 13912 3995 13964 4004
rect 13912 3961 13946 3995
rect 13946 3961 13964 3995
rect 13912 3952 13964 3961
rect 14004 3952 14056 4004
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 12532 3884 12584 3936
rect 14648 3884 14700 3936
rect 17592 3927 17644 3936
rect 17592 3893 17601 3927
rect 17601 3893 17635 3927
rect 17635 3893 17644 3927
rect 17592 3884 17644 3893
rect 17868 3884 17920 3936
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 7840 3680 7892 3732
rect 8576 3723 8628 3732
rect 8576 3689 8585 3723
rect 8585 3689 8619 3723
rect 8619 3689 8628 3723
rect 8576 3680 8628 3689
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 9588 3680 9640 3732
rect 9864 3680 9916 3732
rect 10508 3680 10560 3732
rect 10784 3680 10836 3732
rect 10968 3680 11020 3732
rect 14096 3680 14148 3732
rect 17776 3680 17828 3732
rect 5356 3612 5408 3664
rect 5448 3612 5500 3664
rect 8944 3655 8996 3664
rect 8944 3621 8953 3655
rect 8953 3621 8987 3655
rect 8987 3621 8996 3655
rect 8944 3612 8996 3621
rect 15200 3612 15252 3664
rect 2504 3544 2556 3596
rect 2964 3544 3016 3596
rect 2228 3476 2280 3528
rect 4344 3476 4396 3528
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 2872 3408 2924 3460
rect 3608 3408 3660 3460
rect 3792 3340 3844 3392
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 7656 3544 7708 3596
rect 8484 3476 8536 3528
rect 8944 3476 8996 3528
rect 9312 3476 9364 3528
rect 9496 3476 9548 3528
rect 11980 3544 12032 3596
rect 12072 3544 12124 3596
rect 14004 3544 14056 3596
rect 14832 3544 14884 3596
rect 15660 3544 15712 3596
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 12164 3519 12216 3528
rect 11244 3476 11296 3485
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 7288 3340 7340 3392
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 13912 3408 13964 3460
rect 14740 3408 14792 3460
rect 18052 3408 18104 3460
rect 11152 3340 11204 3392
rect 13636 3340 13688 3392
rect 13820 3383 13872 3392
rect 13820 3349 13829 3383
rect 13829 3349 13863 3383
rect 13863 3349 13872 3383
rect 13820 3340 13872 3349
rect 17408 3383 17460 3392
rect 17408 3349 17417 3383
rect 17417 3349 17451 3383
rect 17451 3349 17460 3383
rect 17408 3340 17460 3349
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 3056 3136 3108 3188
rect 4712 3136 4764 3188
rect 5356 3136 5408 3188
rect 7472 3136 7524 3188
rect 9220 3136 9272 3188
rect 388 3068 440 3120
rect 11152 3136 11204 3188
rect 12624 3136 12676 3188
rect 13636 3136 13688 3188
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 3792 3000 3844 3052
rect 5448 3000 5500 3052
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 8116 3000 8168 3052
rect 8300 3000 8352 3052
rect 9772 3000 9824 3052
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 2780 2864 2832 2916
rect 1492 2796 1544 2848
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 4252 2932 4304 2984
rect 3792 2864 3844 2916
rect 5724 2864 5776 2916
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9588 2932 9640 2984
rect 12072 3068 12124 3120
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 11612 2975 11664 2984
rect 11612 2941 11621 2975
rect 11621 2941 11655 2975
rect 11655 2941 11664 2975
rect 11612 2932 11664 2941
rect 12072 2932 12124 2984
rect 14924 3000 14976 3052
rect 14372 2932 14424 2984
rect 15384 2932 15436 2984
rect 6276 2796 6328 2848
rect 10232 2864 10284 2916
rect 8944 2796 8996 2848
rect 10692 2864 10744 2916
rect 12164 2864 12216 2916
rect 12808 2907 12860 2916
rect 12808 2873 12817 2907
rect 12817 2873 12851 2907
rect 12851 2873 12860 2907
rect 12808 2864 12860 2873
rect 14832 2864 14884 2916
rect 10508 2796 10560 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 13912 2796 13964 2848
rect 16672 2932 16724 2984
rect 16856 2975 16908 2984
rect 16856 2941 16865 2975
rect 16865 2941 16899 2975
rect 16899 2941 16908 2975
rect 16856 2932 16908 2941
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 17776 2796 17828 2848
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 4436 2592 4488 2644
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 4988 2592 5040 2601
rect 5080 2592 5132 2644
rect 8944 2592 8996 2644
rect 11796 2635 11848 2644
rect 11796 2601 11805 2635
rect 11805 2601 11839 2635
rect 11839 2601 11848 2635
rect 11796 2592 11848 2601
rect 4528 2524 4580 2576
rect 4896 2567 4948 2576
rect 4896 2533 4905 2567
rect 4905 2533 4939 2567
rect 4939 2533 4948 2567
rect 4896 2524 4948 2533
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 3332 2499 3384 2508
rect 3332 2465 3341 2499
rect 3341 2465 3375 2499
rect 3375 2465 3384 2499
rect 3332 2456 3384 2465
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 7564 2524 7616 2576
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 11244 2524 11296 2576
rect 11704 2567 11756 2576
rect 11704 2533 11713 2567
rect 11713 2533 11747 2567
rect 11747 2533 11756 2567
rect 16304 2592 16356 2644
rect 11704 2524 11756 2533
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 10692 2499 10744 2508
rect 10692 2465 10701 2499
rect 10701 2465 10735 2499
rect 10735 2465 10744 2499
rect 10692 2456 10744 2465
rect 10876 2456 10928 2508
rect 12256 2456 12308 2508
rect 14188 2456 14240 2508
rect 14648 2499 14700 2508
rect 14648 2465 14657 2499
rect 14657 2465 14691 2499
rect 14691 2465 14700 2499
rect 14648 2456 14700 2465
rect 15016 2456 15068 2508
rect 17684 2499 17736 2508
rect 17684 2465 17693 2499
rect 17693 2465 17727 2499
rect 17727 2465 17736 2499
rect 17684 2456 17736 2465
rect 2136 2388 2188 2440
rect 3608 2431 3660 2440
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 4896 2320 4948 2372
rect 7564 2388 7616 2440
rect 10600 2388 10652 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 13084 2388 13136 2440
rect 8484 2320 8536 2372
rect 8576 2320 8628 2372
rect 6092 2252 6144 2304
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 9772 2252 9824 2304
rect 11244 2320 11296 2372
rect 12348 2252 12400 2304
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 17868 2295 17920 2304
rect 17868 2261 17877 2295
rect 17877 2261 17911 2295
rect 17911 2261 17920 2295
rect 17868 2252 17920 2261
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 3332 2048 3384 2100
rect 9772 2048 9824 2100
rect 10692 2048 10744 2100
rect 13360 2048 13412 2100
rect 8668 1980 8720 2032
rect 13820 1980 13872 2032
rect 3240 1844 3292 1896
rect 5172 1844 5224 1896
rect 10232 1436 10284 1488
rect 19432 1436 19484 1488
<< metal2 >>
rect 1122 16520 1178 17000
rect 3330 16520 3386 17000
rect 5538 16520 5594 17000
rect 7746 16520 7802 17000
rect 9494 16688 9550 16697
rect 9494 16623 9550 16632
rect 1136 13433 1164 16520
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 2134 15056 2190 15065
rect 2134 14991 2190 15000
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1400 13728 1452 13734
rect 1400 13670 1452 13676
rect 1122 13424 1178 13433
rect 1122 13359 1178 13368
rect 1412 10674 1440 13670
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1490 11248 1546 11257
rect 1490 11183 1492 11192
rect 1544 11183 1546 11192
rect 1492 11154 1544 11160
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9722 1440 9998
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 7410 1440 8366
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 7857 1532 7890
rect 1490 7848 1546 7857
rect 1490 7783 1546 7792
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6798 1440 7346
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 5778 1440 6734
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5234 1440 5714
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 4622 1440 5170
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1216 4004 1268 4010
rect 1216 3946 1268 3952
rect 388 3120 440 3126
rect 388 3062 440 3068
rect 400 480 428 3062
rect 1228 480 1256 3946
rect 1504 2854 1532 6054
rect 1596 4078 1624 10406
rect 1688 9518 1716 13330
rect 1780 10606 1808 14214
rect 2056 14074 2084 14418
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 2148 9625 2176 14991
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2240 13530 2268 14350
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2516 13326 2544 13874
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2504 13320 2556 13326
rect 2226 13288 2282 13297
rect 2504 13262 2556 13268
rect 2226 13223 2282 13232
rect 2240 13190 2268 13223
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12782 2268 13126
rect 2516 12866 2544 13262
rect 2608 12889 2636 13330
rect 2424 12850 2544 12866
rect 2412 12844 2544 12850
rect 2464 12838 2544 12844
rect 2594 12880 2650 12889
rect 2594 12815 2650 12824
rect 2412 12786 2464 12792
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2332 12442 2360 12582
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2424 12322 2452 12786
rect 2332 12294 2452 12322
rect 2504 12300 2556 12306
rect 2332 11218 2360 12294
rect 2504 12242 2556 12248
rect 2516 11642 2544 12242
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11762 2636 12174
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2516 11614 2636 11642
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2608 10985 2636 11614
rect 2700 11014 2728 14350
rect 2792 13530 2820 15807
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 11898 2820 13262
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2688 11008 2740 11014
rect 2594 10976 2650 10985
rect 2688 10950 2740 10956
rect 2594 10911 2650 10920
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2516 10266 2544 10610
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2134 9616 2190 9625
rect 2134 9551 2190 9560
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 2516 9450 2544 10202
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 2504 9444 2556 9450
rect 2608 9432 2636 10911
rect 2700 10198 2728 10950
rect 2688 10192 2740 10198
rect 2792 10169 2820 11494
rect 2884 10742 2912 14214
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 12442 3004 13806
rect 3068 12986 3096 14418
rect 3344 14346 3372 16520
rect 3698 16280 3754 16289
rect 3698 16215 3754 16224
rect 3712 15230 3740 16215
rect 4066 15464 4122 15473
rect 4066 15399 4068 15408
rect 4120 15399 4122 15408
rect 5080 15428 5132 15434
rect 4068 15370 4120 15376
rect 5080 15370 5132 15376
rect 3700 15224 3752 15230
rect 3700 15166 3752 15172
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3238 14240 3294 14249
rect 3238 14175 3294 14184
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 3160 11830 3188 13330
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3146 11384 3202 11393
rect 2964 11348 3016 11354
rect 3146 11319 3202 11328
rect 2964 11290 3016 11296
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2688 10134 2740 10140
rect 2778 10160 2834 10169
rect 2834 10118 2912 10146
rect 2778 10095 2834 10104
rect 2688 9444 2740 9450
rect 2608 9404 2688 9432
rect 2504 9386 2556 9392
rect 2688 9386 2740 9392
rect 1964 9178 1992 9386
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2596 8968 2648 8974
rect 2226 8936 2282 8945
rect 2596 8910 2648 8916
rect 2226 8871 2282 8880
rect 1674 8528 1730 8537
rect 1674 8463 1730 8472
rect 1688 6866 1716 8463
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1780 5914 1808 6054
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1952 4616 2004 4622
rect 1952 4558 2004 4564
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 4321 1716 4422
rect 1674 4312 1730 4321
rect 1674 4247 1730 4256
rect 1964 4146 1992 4558
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1582 3904 1638 3913
rect 1582 3839 1638 3848
rect 1596 3738 1624 3839
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1688 2650 1716 3431
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 2056 2514 2084 6054
rect 2240 3534 2268 8871
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2424 8022 2452 8774
rect 2608 8566 2636 8910
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2332 6458 2360 6734
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2516 5681 2544 8298
rect 2792 6361 2820 8842
rect 2884 8498 2912 10118
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2976 8401 3004 11290
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2962 8392 3018 8401
rect 2962 8327 3018 8336
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 7886 2912 8230
rect 2872 7880 2924 7886
rect 2924 7828 3004 7834
rect 2872 7822 3004 7828
rect 2884 7806 3004 7822
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2778 6352 2834 6361
rect 2596 6316 2648 6322
rect 2884 6322 2912 7686
rect 2976 7342 3004 7806
rect 3068 7585 3096 10406
rect 3160 8090 3188 11319
rect 3252 10674 3280 14175
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3344 10606 3372 14010
rect 3436 13530 3464 14350
rect 3712 13841 3740 14486
rect 3804 14074 3832 14826
rect 4342 14648 4398 14657
rect 4342 14583 4398 14592
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3698 13832 3754 13841
rect 3698 13767 3754 13776
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3712 13025 3740 13194
rect 3698 13016 3754 13025
rect 3804 12986 3832 13874
rect 4264 13802 4292 14214
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3698 12951 3754 12960
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12238 3648 12650
rect 3712 12238 3740 12718
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11626 3464 12038
rect 3606 11792 3662 11801
rect 3606 11727 3662 11736
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3516 11552 3568 11558
rect 3436 11500 3516 11506
rect 3436 11494 3568 11500
rect 3436 11478 3556 11494
rect 3436 11354 3464 11478
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3054 7576 3110 7585
rect 3054 7511 3110 7520
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 6866 3096 7142
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2778 6287 2834 6296
rect 2872 6316 2924 6322
rect 2596 6258 2648 6264
rect 2872 6258 2924 6264
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2516 3602 2544 5607
rect 2608 5574 2636 6258
rect 2780 6248 2832 6254
rect 2778 6216 2780 6225
rect 2832 6216 2834 6225
rect 2778 6151 2834 6160
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2608 5234 2636 5510
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4690 2820 4966
rect 2976 4729 3004 6598
rect 3068 6304 3096 6802
rect 3160 6458 3188 6870
rect 3252 6769 3280 9862
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3344 9081 3372 9687
rect 3436 9353 3464 11290
rect 3620 10690 3648 11727
rect 3712 11694 3740 12174
rect 3804 11694 3832 12922
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4172 12209 4200 12310
rect 4158 12200 4214 12209
rect 4158 12135 4214 12144
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3882 11792 3938 11801
rect 4356 11778 4384 14583
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4724 14074 4752 14418
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4724 13258 4752 13738
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4632 12918 4660 13126
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4724 12730 4752 13194
rect 3882 11727 3938 11736
rect 4264 11750 4384 11778
rect 4632 12702 4752 12730
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3712 11286 3740 11630
rect 3896 11354 3924 11727
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3712 11132 3740 11222
rect 3792 11144 3844 11150
rect 3712 11104 3792 11132
rect 3792 11086 3844 11092
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3712 10810 3740 10950
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3620 10662 3740 10690
rect 3608 10600 3660 10606
rect 3514 10568 3570 10577
rect 3608 10542 3660 10548
rect 3514 10503 3570 10512
rect 3528 9654 3556 10503
rect 3620 10266 3648 10542
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3516 9376 3568 9382
rect 3422 9344 3478 9353
rect 3516 9318 3568 9324
rect 3422 9279 3478 9288
rect 3330 9072 3386 9081
rect 3330 9007 3332 9016
rect 3384 9007 3386 9016
rect 3332 8978 3384 8984
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3332 8900 3384 8906
rect 3332 8842 3384 8848
rect 3344 7206 3372 8842
rect 3436 8634 3464 8910
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3436 8401 3464 8434
rect 3422 8392 3478 8401
rect 3422 8327 3478 8336
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3238 6760 3294 6769
rect 3238 6695 3294 6704
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3436 6322 3464 8327
rect 3148 6316 3200 6322
rect 3068 6276 3148 6304
rect 3148 6258 3200 6264
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2962 4720 3018 4729
rect 2780 4684 2832 4690
rect 2962 4655 3018 4664
rect 2780 4626 2832 4632
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2884 3466 2912 3946
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2148 480 2176 2382
rect 386 0 442 480
rect 1214 0 1270 480
rect 2134 0 2190 480
rect 2792 241 2820 2858
rect 2976 2650 3004 3538
rect 3068 3194 3096 5102
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3056 2848 3108 2854
rect 3054 2816 3056 2825
rect 3108 2816 3110 2825
rect 3054 2751 3110 2760
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3160 1442 3188 5034
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3252 3058 3280 4626
rect 3436 3097 3464 5510
rect 3528 5273 3556 9318
rect 3606 8936 3662 8945
rect 3606 8871 3662 8880
rect 3620 8498 3648 8871
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3620 8265 3648 8434
rect 3606 8256 3662 8265
rect 3606 8191 3662 8200
rect 3606 8120 3662 8129
rect 3606 8055 3662 8064
rect 3620 8022 3648 8055
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3514 5264 3570 5273
rect 3620 5250 3648 7686
rect 3712 5778 3740 10662
rect 3804 10470 3832 11086
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 4068 10600 4120 10606
rect 4066 10568 4068 10577
rect 4120 10568 4122 10577
rect 4066 10503 4122 10512
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 10130 3832 10406
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3804 9722 3832 10066
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 3792 9716 3844 9722
rect 4264 9704 4292 11750
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 3792 9658 3844 9664
rect 4172 9676 4292 9704
rect 3804 8974 3832 9658
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 9110 4108 9318
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3792 8968 3844 8974
rect 4172 8945 4200 9676
rect 4356 9586 4384 11630
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 3792 8910 3844 8916
rect 4158 8936 4214 8945
rect 3804 8634 3832 8910
rect 4158 8871 4214 8880
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 4264 8498 4292 9046
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7993 4108 8230
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 4158 7440 4214 7449
rect 4158 7375 4214 7384
rect 4172 7342 4200 7375
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 6798 4108 7210
rect 4356 7177 4384 9318
rect 4448 9178 4476 9862
rect 4632 9518 4660 12702
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12442 4752 12582
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4710 12200 4766 12209
rect 4710 12135 4766 12144
rect 4724 11830 4752 12135
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4724 10810 4752 11562
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4540 9081 4568 9454
rect 4526 9072 4582 9081
rect 4526 9007 4582 9016
rect 4434 8936 4490 8945
rect 4724 8922 4752 10542
rect 4816 9586 4844 13806
rect 5092 13376 5120 15370
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5184 13530 5212 14350
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5172 13388 5224 13394
rect 5092 13348 5172 13376
rect 5172 13330 5224 13336
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4908 10606 4936 13262
rect 5184 13025 5212 13330
rect 5170 13016 5226 13025
rect 5170 12951 5226 12960
rect 5276 12646 5304 14350
rect 5552 14090 5580 16520
rect 5908 15224 5960 15230
rect 5908 15166 5960 15172
rect 5356 14068 5408 14074
rect 5552 14062 5856 14090
rect 5356 14010 5408 14016
rect 5368 12782 5396 14010
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5264 12640 5316 12646
rect 5460 12628 5488 12786
rect 5264 12582 5316 12588
rect 5368 12600 5488 12628
rect 5276 12442 5304 12582
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5368 12374 5396 12600
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5552 12306 5580 13942
rect 5828 13802 5856 14062
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 12442 5672 13670
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5736 12850 5764 13194
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5828 12322 5856 12582
rect 5920 12374 5948 15166
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 6090 13832 6146 13841
rect 6090 13767 6146 13776
rect 6104 13734 6132 13767
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6196 13530 6224 13670
rect 6380 13546 6408 13670
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6288 13518 6408 13546
rect 6288 13462 6316 13518
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5644 12294 5856 12322
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11218 5120 11494
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9761 4936 9998
rect 5000 9926 5028 10610
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4894 9752 4950 9761
rect 5092 9722 5120 10406
rect 5170 10160 5226 10169
rect 5170 10095 5226 10104
rect 4894 9687 4950 9696
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5184 9654 5212 10095
rect 5172 9648 5224 9654
rect 4986 9616 5042 9625
rect 4804 9580 4856 9586
rect 5172 9590 5224 9596
rect 4986 9551 5042 9560
rect 4804 9522 4856 9528
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4434 8871 4490 8880
rect 4540 8894 4752 8922
rect 4448 7954 4476 8871
rect 4540 8537 4568 8894
rect 4712 8832 4764 8838
rect 4632 8792 4712 8820
rect 4526 8528 4582 8537
rect 4526 8463 4582 8472
rect 4632 8430 4660 8792
rect 4712 8774 4764 8780
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4342 7168 4398 7177
rect 4342 7103 4398 7112
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 5953 3832 6598
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 3790 5944 3846 5953
rect 3790 5879 3846 5888
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3698 5536 3754 5545
rect 3698 5471 3754 5480
rect 3712 5370 3740 5471
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4264 5370 4292 6326
rect 4356 5710 4384 6938
rect 4448 6458 4476 7890
rect 4540 7449 4568 8230
rect 4632 7886 4660 8366
rect 4816 8129 4844 9318
rect 4802 8120 4858 8129
rect 4802 8055 4858 8064
rect 4804 7948 4856 7954
rect 4724 7908 4804 7936
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4526 7440 4582 7449
rect 4526 7375 4582 7384
rect 4632 7342 4660 7822
rect 4724 7546 4752 7908
rect 4804 7890 4856 7896
rect 5000 7834 5028 9551
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 4816 7806 5028 7834
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4526 7032 4582 7041
rect 4526 6967 4582 6976
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4448 5624 4476 6258
rect 4540 6225 4568 6967
rect 4526 6216 4582 6225
rect 4526 6151 4582 6160
rect 4618 5944 4674 5953
rect 4618 5879 4620 5888
rect 4672 5879 4674 5888
rect 4620 5850 4672 5856
rect 4528 5636 4580 5642
rect 4448 5596 4528 5624
rect 4528 5578 4580 5584
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4434 5264 4490 5273
rect 3620 5222 3740 5250
rect 3514 5199 3570 5208
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3422 3088 3478 3097
rect 3240 3052 3292 3058
rect 3422 3023 3478 3032
rect 3240 2994 3292 3000
rect 3422 2952 3478 2961
rect 3422 2887 3478 2896
rect 3436 2650 3464 2887
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3344 2106 3372 2450
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 3240 1896 3292 1902
rect 3238 1864 3240 1873
rect 3292 1864 3294 1873
rect 3238 1799 3294 1808
rect 3068 1414 3188 1442
rect 3068 480 3096 1414
rect 3528 1057 3556 3946
rect 3620 3466 3648 4422
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3620 2446 3648 3402
rect 3712 2553 3740 5222
rect 4540 5234 4568 5578
rect 4434 5199 4436 5208
rect 4488 5199 4490 5208
rect 4528 5228 4580 5234
rect 4436 5170 4488 5176
rect 4528 5170 4580 5176
rect 4816 5137 4844 7806
rect 4896 7744 4948 7750
rect 5080 7744 5132 7750
rect 4948 7692 5028 7698
rect 4896 7686 5028 7692
rect 5080 7686 5132 7692
rect 4908 7670 5028 7686
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4908 5574 4936 7414
rect 5000 7002 5028 7670
rect 5092 7041 5120 7686
rect 5078 7032 5134 7041
rect 4988 6996 5040 7002
rect 5078 6967 5134 6976
rect 4988 6938 5040 6944
rect 5184 6746 5212 9454
rect 5276 8634 5304 10610
rect 5368 10062 5396 10610
rect 5460 10266 5488 11591
rect 5644 11354 5672 12294
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5368 9586 5396 9998
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5276 8362 5304 8570
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5276 7546 5304 8298
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5368 7274 5396 9522
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5000 6718 5212 6746
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4250 5128 4306 5137
rect 4250 5063 4252 5072
rect 4304 5063 4306 5072
rect 4802 5128 4858 5137
rect 4802 5063 4858 5072
rect 4252 5034 4304 5040
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4894 4992 4950 5001
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 4264 4214 4292 4694
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4356 4282 4384 4626
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4356 3534 4384 4218
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 3804 3058 3832 3334
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 4264 2990 4292 3334
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3698 2544 3754 2553
rect 3698 2479 3754 2488
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3514 1048 3570 1057
rect 3514 983 3570 992
rect 3804 898 3832 2858
rect 4448 2650 4476 4694
rect 4540 4282 4568 4966
rect 4894 4927 4950 4936
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4540 2582 4568 4218
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 3738 4660 3878
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 3194 4752 3470
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4908 2582 4936 4927
rect 5000 2650 5028 6718
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5092 4554 5120 6394
rect 5184 6322 5212 6598
rect 5276 6458 5304 6938
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5368 6322 5396 6802
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5368 6066 5396 6122
rect 5276 6038 5396 6066
rect 5276 5914 5304 6038
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5262 5808 5318 5817
rect 5262 5743 5264 5752
rect 5316 5743 5318 5752
rect 5264 5714 5316 5720
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 4548 5132 4554
rect 5080 4490 5132 4496
rect 5078 2680 5134 2689
rect 4988 2644 5040 2650
rect 5078 2615 5080 2624
rect 4988 2586 5040 2592
rect 5132 2615 5134 2624
rect 5080 2586 5132 2592
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 3804 870 4016 898
rect 3988 480 4016 870
rect 4908 480 4936 2314
rect 5184 1902 5212 5306
rect 5276 5030 5304 5510
rect 5460 5030 5488 9930
rect 5552 9042 5580 10406
rect 5644 10033 5672 11290
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5630 10024 5686 10033
rect 5630 9959 5686 9968
rect 5736 9654 5764 11086
rect 5814 10840 5870 10849
rect 5814 10775 5870 10784
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5630 9480 5686 9489
rect 5630 9415 5686 9424
rect 5724 9444 5776 9450
rect 5644 9382 5672 9415
rect 5724 9386 5776 9392
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5630 9208 5686 9217
rect 5630 9143 5686 9152
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 4146 5488 4422
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3670 5488 4082
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5368 3194 5396 3606
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5460 3058 5488 3606
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5552 2514 5580 7686
rect 5644 6254 5672 9143
rect 5736 8838 5764 9386
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5828 7857 5856 10775
rect 5814 7848 5870 7857
rect 5814 7783 5870 7792
rect 5828 6798 5856 7783
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 4570 5856 6054
rect 5644 4542 5856 4570
rect 5644 4010 5672 4542
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 4078 5764 4422
rect 5920 4078 5948 11494
rect 6012 10169 6040 13262
rect 6092 12368 6144 12374
rect 6092 12310 6144 12316
rect 6104 10470 6132 12310
rect 6380 12288 6408 13398
rect 6472 13190 6500 13874
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13462 6776 13738
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 7484 13530 7512 13874
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6472 12442 6500 12854
rect 6656 12782 6684 13262
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6380 12260 6592 12288
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 5998 10160 6054 10169
rect 5998 10095 6054 10104
rect 6196 9654 6224 12038
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6196 9466 6224 9590
rect 6104 9438 6224 9466
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6012 5001 6040 6734
rect 6104 6118 6132 9438
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 8634 6224 9318
rect 6288 9110 6316 11630
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6288 8566 6316 9046
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6196 7206 6224 7414
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5998 4992 6054 5001
rect 5998 4927 6054 4936
rect 6196 4826 6224 7142
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6288 5273 6316 5306
rect 6274 5264 6330 5273
rect 6274 5199 6330 5208
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4826 6316 4966
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5644 2904 5672 3946
rect 5724 2916 5776 2922
rect 5644 2876 5724 2904
rect 5724 2858 5776 2864
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 5828 480 5856 3946
rect 6196 3058 6224 4558
rect 6274 4176 6330 4185
rect 6274 4111 6330 4120
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6104 2310 6132 2994
rect 6288 2854 6316 4111
rect 6380 4078 6408 11018
rect 6472 9382 6500 11834
rect 6564 10849 6592 12260
rect 6656 11558 6684 12718
rect 7484 12714 7512 13466
rect 7760 13462 7788 16520
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 14074 8156 14214
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 6734 12608 6790 12617
rect 6734 12543 6790 12552
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6550 10840 6606 10849
rect 6550 10775 6606 10784
rect 6656 10674 6684 11494
rect 6748 11121 6776 12543
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7024 11801 7052 12174
rect 7010 11792 7066 11801
rect 7010 11727 7066 11736
rect 7196 11688 7248 11694
rect 7194 11656 7196 11665
rect 7248 11656 7250 11665
rect 7194 11591 7250 11600
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 7012 11144 7064 11150
rect 6734 11112 6790 11121
rect 7012 11086 7064 11092
rect 6734 11047 6790 11056
rect 6826 10976 6882 10985
rect 6826 10911 6882 10920
rect 6840 10810 6868 10911
rect 7024 10810 7052 11086
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6644 10668 6696 10674
rect 6564 10628 6644 10656
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 5953 6500 9318
rect 6564 9042 6592 10628
rect 6644 10610 6696 10616
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6656 8430 6684 10134
rect 6748 9994 6776 10474
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6748 9586 6776 9930
rect 7024 9625 7052 10134
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7010 9616 7066 9625
rect 6736 9580 6788 9586
rect 7208 9586 7236 10066
rect 7010 9551 7066 9560
rect 7196 9580 7248 9586
rect 6736 9522 6788 9528
rect 7196 9522 7248 9528
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 9110 6776 9318
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 7300 9178 7328 12174
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6550 8256 6606 8265
rect 6550 8191 6606 8200
rect 6564 7410 6592 8191
rect 6748 7954 6776 8910
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6918 8392 6974 8401
rect 6918 8327 6920 8336
rect 6972 8327 6974 8336
rect 6920 8298 6972 8304
rect 7116 8276 7144 8774
rect 7392 8362 7420 12038
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7484 11665 7512 11766
rect 7470 11656 7526 11665
rect 7470 11591 7526 11600
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7484 10198 7512 11222
rect 7576 10538 7604 11494
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7668 10248 7696 12310
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7760 11354 7788 11562
rect 7852 11354 7880 13670
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8128 12889 8156 13398
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8220 12918 8248 13126
rect 8208 12912 8260 12918
rect 8114 12880 8170 12889
rect 8208 12854 8260 12860
rect 8114 12815 8170 12824
rect 8128 12730 8156 12815
rect 8128 12702 8248 12730
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8036 11218 8064 12038
rect 8128 11694 8156 12174
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8114 11248 8170 11257
rect 8024 11212 8076 11218
rect 8114 11183 8170 11192
rect 8024 11154 8076 11160
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7576 10220 7696 10248
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7484 8294 7512 9862
rect 7576 9722 7604 10220
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7576 9450 7604 9658
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7472 8288 7524 8294
rect 7116 8248 7328 8276
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7300 7970 7328 8248
rect 7472 8230 7524 8236
rect 6736 7948 6788 7954
rect 7300 7942 7420 7970
rect 6736 7890 6788 7896
rect 6644 7880 6696 7886
rect 7288 7880 7340 7886
rect 6644 7822 6696 7828
rect 6734 7848 6790 7857
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6656 7002 6684 7822
rect 7288 7822 7340 7828
rect 6734 7783 6790 7792
rect 6748 7206 6776 7783
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6748 6882 6776 7142
rect 6886 7100 7182 7120
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6656 6854 6776 6882
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6458 5944 6514 5953
rect 6458 5879 6514 5888
rect 6472 5166 6500 5879
rect 6564 5778 6592 6054
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6656 5681 6684 6854
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6458 6868 6734
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6748 6338 6776 6394
rect 6748 6310 6960 6338
rect 6932 6186 6960 6310
rect 7300 6186 7328 7822
rect 7392 7449 7420 7942
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7378 7440 7434 7449
rect 7378 7375 7434 7384
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 6798 7420 7278
rect 7484 6866 7512 7822
rect 7576 7410 7604 8774
rect 7668 8634 7696 10066
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7300 5914 7328 6122
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7286 5808 7342 5817
rect 7196 5772 7248 5778
rect 7286 5743 7288 5752
rect 7196 5714 7248 5720
rect 7340 5743 7342 5752
rect 7288 5714 7340 5720
rect 7208 5681 7236 5714
rect 7392 5710 7420 6734
rect 7484 5914 7512 6802
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7380 5704 7432 5710
rect 6642 5672 6698 5681
rect 6642 5607 6698 5616
rect 7194 5672 7250 5681
rect 7250 5630 7328 5658
rect 7380 5646 7432 5652
rect 7194 5607 7250 5616
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6472 4146 6500 5102
rect 6748 5080 6776 5170
rect 6920 5092 6972 5098
rect 6748 5052 6920 5080
rect 6920 5034 6972 5040
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6276 2848 6328 2854
rect 6564 2825 6592 4966
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6276 2790 6328 2796
rect 6550 2816 6606 2825
rect 6550 2751 6606 2760
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 6656 1034 6684 3946
rect 6748 3942 6776 4422
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 7300 3398 7328 5630
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 6656 1006 6776 1034
rect 6748 480 6776 1006
rect 7392 649 7420 5510
rect 7576 5386 7604 7346
rect 7668 5642 7696 8570
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7576 5358 7696 5386
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7484 4758 7512 5238
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7484 3194 7512 4694
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7576 2582 7604 5102
rect 7668 3602 7696 5358
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7760 2514 7788 11018
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7852 9976 7880 10542
rect 7944 10452 7972 11086
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 8036 10606 8064 11018
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 7944 10424 8064 10452
rect 7852 9948 7972 9976
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7852 8430 7880 9687
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7838 8256 7894 8265
rect 7838 8191 7894 8200
rect 7852 5794 7880 8191
rect 7944 7750 7972 9948
rect 8036 8838 8064 10424
rect 8128 9518 8156 11183
rect 8220 10130 8248 12702
rect 8312 11286 8340 13126
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12238 8432 12582
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8390 11520 8446 11529
rect 8390 11455 8446 11464
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8312 9926 8340 10542
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8220 9178 8248 9522
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 8650 8156 8774
rect 8036 8622 8156 8650
rect 8036 8401 8064 8622
rect 8220 8498 8248 9114
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8404 8401 8432 11455
rect 8496 11014 8524 13670
rect 8680 11218 8708 13806
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8574 11112 8630 11121
rect 8574 11047 8630 11056
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8496 9081 8524 9522
rect 8588 9518 8616 11047
rect 8668 11008 8720 11014
rect 8666 10976 8668 10985
rect 8720 10976 8722 10985
rect 8666 10911 8722 10920
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8680 9722 8708 9862
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8482 9072 8538 9081
rect 8482 9007 8538 9016
rect 8022 8392 8078 8401
rect 8390 8392 8446 8401
rect 8022 8327 8078 8336
rect 8116 8356 8168 8362
rect 8390 8327 8446 8336
rect 8116 8298 8168 8304
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7930 7440 7986 7449
rect 7930 7375 7986 7384
rect 7944 6186 7972 7375
rect 8036 7206 8064 7754
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7852 5766 7972 5794
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7852 4622 7880 5646
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7852 3738 7880 4558
rect 7944 4078 7972 5766
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8036 3942 8064 4082
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8128 3058 8156 8298
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7954 8432 8230
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 6866 8248 7346
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 7002 8340 7210
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8220 6458 8248 6802
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5574 8248 6054
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8206 5400 8262 5409
rect 8206 5335 8262 5344
rect 8220 5166 8248 5335
rect 8312 5273 8340 6122
rect 8298 5264 8354 5273
rect 8298 5199 8300 5208
rect 8352 5199 8354 5208
rect 8300 5170 8352 5176
rect 8208 5160 8260 5166
rect 8312 5139 8340 5170
rect 8208 5102 8260 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4758 8340 4966
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8312 4146 8340 4694
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8312 3398 8340 4082
rect 8496 3534 8524 9007
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8588 3738 8616 7958
rect 8680 7478 8708 7958
rect 8772 7954 8800 13874
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8864 9761 8892 13806
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13530 9168 13670
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9048 12442 9076 13262
rect 9140 12646 9168 13262
rect 9232 12782 9260 13874
rect 9416 13870 9444 14758
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9324 13530 9352 13738
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9508 13326 9536 16623
rect 9954 16520 10010 17000
rect 12162 16520 12218 17000
rect 14370 16520 14426 17000
rect 16578 16520 16634 17000
rect 17958 16688 18014 16697
rect 17958 16623 18014 16632
rect 9968 14414 9996 16520
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9496 13320 9548 13326
rect 9416 13280 9496 13308
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9232 12238 9260 12718
rect 9036 12232 9088 12238
rect 9034 12200 9036 12209
rect 9220 12232 9272 12238
rect 9088 12200 9090 12209
rect 9220 12174 9272 12180
rect 9034 12135 9090 12144
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 11082 8984 11494
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8956 10538 8984 11018
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 9048 10130 9076 12135
rect 9232 11762 9260 12174
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9324 11898 9352 12038
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8850 9752 8906 9761
rect 8850 9687 8906 9696
rect 8956 9654 8984 10066
rect 9232 9722 9260 10406
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8772 7342 8800 7890
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8680 3942 8708 6326
rect 8864 5370 8892 6870
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8772 5137 8800 5170
rect 8758 5128 8814 5137
rect 8758 5063 8814 5072
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8956 3670 8984 6054
rect 9232 5166 9260 9454
rect 9324 9450 9352 11562
rect 9416 10724 9444 13280
rect 9496 13262 9548 13268
rect 9494 13016 9550 13025
rect 9494 12951 9550 12960
rect 9508 12918 9536 12951
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9508 11257 9536 11834
rect 9494 11248 9550 11257
rect 9494 11183 9550 11192
rect 9416 10696 9536 10724
rect 9508 10198 9536 10696
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9324 7546 9352 7822
rect 9416 7546 9444 10066
rect 9600 9654 9628 13806
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9692 12442 9720 13738
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 10152 13462 10180 13631
rect 10336 13462 10364 14486
rect 10888 14278 10916 14826
rect 11794 14512 11850 14521
rect 11794 14447 11850 14456
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10140 13456 10192 13462
rect 10140 13398 10192 13404
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9784 12374 9812 13126
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 10244 12832 10272 13126
rect 9876 12804 10272 12832
rect 10336 12832 10364 13398
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12986 10456 13262
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10336 12804 10456 12832
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9876 12152 9904 12804
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9692 12124 9904 12152
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9508 7750 9536 7890
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9416 6458 9444 7482
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9402 5264 9458 5273
rect 9402 5199 9458 5208
rect 9220 5160 9272 5166
rect 9218 5128 9220 5137
rect 9272 5128 9274 5137
rect 9416 5098 9444 5199
rect 9218 5063 9274 5072
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9048 3738 9076 4762
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9324 4146 9352 4490
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8312 3058 8340 3334
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8956 2990 8984 3470
rect 9232 3194 9260 3878
rect 9324 3534 9352 4082
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8956 2650 8984 2790
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7378 640 7434 649
rect 7378 575 7434 584
rect 7576 480 7604 2382
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8496 480 8524 2314
rect 8588 1465 8616 2314
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 2038 8708 2246
rect 8668 2032 8720 2038
rect 8668 1974 8720 1980
rect 8574 1456 8630 1465
rect 8574 1391 8630 1400
rect 9416 480 9444 4082
rect 9508 3534 9536 7686
rect 9600 7002 9628 7686
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 5234 9628 5714
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4554 9628 5170
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9692 3890 9720 12124
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10138 11792 10194 11801
rect 10138 11727 10194 11736
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11354 9812 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 10152 11218 10180 11727
rect 10244 11694 10272 12582
rect 10336 11694 10364 12650
rect 10428 12646 10456 12804
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10230 11248 10286 11257
rect 10140 11212 10192 11218
rect 10230 11183 10232 11192
rect 10140 11154 10192 11160
rect 10284 11183 10286 11192
rect 10232 11154 10284 11160
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 10138 11112 10194 11121
rect 9784 10810 9812 11086
rect 10138 11047 10140 11056
rect 10192 11047 10194 11056
rect 10232 11076 10284 11082
rect 10140 11018 10192 11024
rect 10232 11018 10284 11024
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 10244 10606 10272 11018
rect 10336 10985 10364 11494
rect 10428 11082 10456 12038
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10322 10976 10378 10985
rect 10322 10911 10378 10920
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 9784 10130 9812 10542
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 10322 9616 10378 9625
rect 10322 9551 10378 9560
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9784 7993 9812 9386
rect 10336 9382 10364 9551
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 9876 9081 9904 9318
rect 9862 9072 9918 9081
rect 9862 9007 9918 9016
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 9770 7984 9826 7993
rect 9770 7919 9826 7928
rect 10046 7984 10102 7993
rect 10046 7919 10048 7928
rect 10100 7919 10102 7928
rect 10048 7890 10100 7896
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6186 9812 7142
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6769 10088 6802
rect 10046 6760 10102 6769
rect 10046 6695 10102 6704
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9784 4162 9812 6122
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 10244 5370 10272 8026
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10336 5030 10364 9318
rect 10414 9208 10470 9217
rect 10520 9178 10548 13670
rect 10704 13462 10732 14010
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10612 12442 10640 13262
rect 10796 13138 10824 14214
rect 11150 13968 11206 13977
rect 11150 13903 11206 13912
rect 11520 13932 11572 13938
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10704 13110 10824 13138
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 9489 10640 11494
rect 10598 9480 10654 9489
rect 10598 9415 10654 9424
rect 10414 9143 10470 9152
rect 10508 9172 10560 9178
rect 10428 9042 10456 9143
rect 10508 9114 10560 9120
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7410 10548 7822
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10520 6934 10548 7346
rect 10612 7002 10640 9415
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10520 6254 10548 6870
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5846 10548 6190
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 9852 4380 10148 4400
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 9784 4134 9996 4162
rect 9692 3862 9904 3890
rect 9876 3738 9904 3862
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9600 2990 9628 3674
rect 9968 3618 9996 4134
rect 10244 4049 10272 4966
rect 10336 4214 10364 4966
rect 10520 4758 10548 5782
rect 10598 5672 10654 5681
rect 10598 5607 10654 5616
rect 10612 4826 10640 5607
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10508 4752 10560 4758
rect 10414 4720 10470 4729
rect 10508 4694 10560 4700
rect 10414 4655 10470 4664
rect 10428 4282 10456 4655
rect 10598 4448 10654 4457
rect 10598 4383 10654 4392
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10230 4040 10286 4049
rect 10612 4010 10640 4383
rect 10230 3975 10286 3984
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 9784 3590 9996 3618
rect 9784 3058 9812 3590
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9784 2310 9812 2450
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 2106 9812 2246
rect 9852 2204 10148 2224
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 10244 1494 10272 2858
rect 10520 2854 10548 3674
rect 10612 3097 10640 3946
rect 10598 3088 10654 3097
rect 10598 3023 10654 3032
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10612 2446 10640 3023
rect 10704 2922 10732 13110
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10796 12374 10824 12786
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 10810 10824 12310
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10888 8090 10916 13330
rect 11164 13258 11192 13903
rect 11520 13874 11572 13880
rect 11532 13326 11560 13874
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11520 13320 11572 13326
rect 11256 13280 11520 13308
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 11744 11008 12718
rect 10980 11716 11100 11744
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10980 11150 11008 11562
rect 11072 11558 11100 11716
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10130 11008 10406
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9586 11008 10066
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 8974 11008 9522
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10980 7018 11008 8774
rect 11072 8634 11100 10746
rect 11164 9897 11192 11222
rect 11256 10266 11284 13280
rect 11624 13297 11652 13330
rect 11520 13262 11572 13268
rect 11610 13288 11666 13297
rect 11610 13223 11666 13232
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11440 12345 11468 12650
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11426 12336 11482 12345
rect 11348 12294 11426 12322
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11150 9888 11206 9897
rect 11150 9823 11206 9832
rect 11256 9722 11284 10202
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11164 8294 11192 9522
rect 11348 9058 11376 12294
rect 11426 12271 11482 12280
rect 11532 12209 11560 12582
rect 11518 12200 11574 12209
rect 11518 12135 11574 12144
rect 11624 11898 11652 13223
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11716 11694 11744 12038
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11518 11384 11574 11393
rect 11518 11319 11574 11328
rect 11256 9030 11376 9058
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 10980 6990 11100 7018
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10796 4554 10824 5102
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 4826 10916 4966
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10704 2106 10732 2450
rect 10796 2446 10824 3674
rect 10888 3040 10916 4626
rect 10980 3738 11008 6870
rect 11072 4593 11100 6990
rect 11256 6202 11284 9030
rect 11532 8650 11560 11319
rect 11164 6174 11284 6202
rect 11440 8622 11560 8650
rect 11058 4584 11114 4593
rect 11058 4519 11114 4528
rect 11060 4480 11112 4486
rect 11058 4448 11060 4457
rect 11112 4448 11114 4457
rect 11058 4383 11114 4392
rect 11164 4185 11192 6174
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 5778 11284 6054
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11150 4176 11206 4185
rect 11150 4111 11206 4120
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11256 3534 11284 5714
rect 11440 5302 11468 8622
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11532 6798 11560 8502
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 3194 11192 3334
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 3052 11112 3058
rect 10888 3012 11060 3040
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10232 1488 10284 1494
rect 10232 1430 10284 1436
rect 10888 1306 10916 2450
rect 10980 2446 11008 3012
rect 11060 2994 11112 3000
rect 11348 2666 11376 4422
rect 11624 2990 11652 11494
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 9178 11744 9318
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11808 8090 11836 14447
rect 12176 13462 12204 16520
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 14384 14550 14412 16520
rect 15566 15872 15622 15881
rect 15566 15807 15622 15816
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13542 14376 13598 14385
rect 13372 13870 13400 14350
rect 13542 14311 13598 14320
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 12348 13728 12400 13734
rect 12346 13696 12348 13705
rect 12400 13696 12402 13705
rect 12346 13631 12402 13640
rect 12164 13456 12216 13462
rect 12728 13433 12756 13806
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12164 13398 12216 13404
rect 12714 13424 12770 13433
rect 12714 13359 12770 13368
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12532 12776 12584 12782
rect 12584 12736 12664 12764
rect 12532 12718 12584 12724
rect 12084 12430 12296 12458
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11992 10146 12020 12310
rect 12084 11393 12112 12430
rect 12162 12336 12218 12345
rect 12162 12271 12164 12280
rect 12216 12271 12218 12280
rect 12164 12242 12216 12248
rect 12268 12209 12296 12430
rect 12254 12200 12310 12209
rect 12360 12186 12388 12718
rect 12360 12158 12480 12186
rect 12254 12135 12310 12144
rect 12070 11384 12126 11393
rect 12070 11319 12126 11328
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 10810 12388 10950
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12452 10554 12480 12158
rect 12636 11778 12664 12736
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12728 11898 12756 12174
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12636 11750 12756 11778
rect 12622 11656 12678 11665
rect 12622 11591 12678 11600
rect 12728 11642 12756 11750
rect 13188 11665 13216 12174
rect 12806 11656 12862 11665
rect 12728 11614 12806 11642
rect 12636 11014 12664 11591
rect 12728 11132 12756 11614
rect 12806 11591 12862 11600
rect 13174 11656 13230 11665
rect 13174 11591 13230 11600
rect 13280 11558 13308 13466
rect 13372 12900 13400 13806
rect 13452 12912 13504 12918
rect 13372 12872 13452 12900
rect 13452 12854 13504 12860
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13176 11552 13228 11558
rect 13268 11552 13320 11558
rect 13176 11494 13228 11500
rect 13266 11520 13268 11529
rect 13320 11520 13322 11529
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12808 11144 12860 11150
rect 12728 11104 12808 11132
rect 12808 11086 12860 11092
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12820 10826 12848 11086
rect 12636 10798 12848 10826
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12268 10526 12480 10554
rect 11992 10118 12112 10146
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11808 6186 11836 8026
rect 11900 8022 11928 8434
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 11900 7546 11928 7958
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11992 7426 12020 9998
rect 12084 8480 12112 10118
rect 12268 8786 12296 10526
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9761 12388 9862
rect 12346 9752 12402 9761
rect 12346 9687 12402 9696
rect 12348 9512 12400 9518
rect 12452 9500 12480 10406
rect 12544 10198 12572 10678
rect 12636 10538 12664 10798
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12400 9472 12480 9500
rect 12544 9489 12572 10134
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12530 9480 12586 9489
rect 12348 9454 12400 9460
rect 12728 9450 12756 9998
rect 13188 9994 13216 11494
rect 13266 11455 13322 11464
rect 13372 11354 13400 11766
rect 13556 11762 13584 14311
rect 14384 14090 14412 14486
rect 15580 14414 15608 15807
rect 16302 15464 16358 15473
rect 16302 15399 16358 15408
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15120 14278 15148 14350
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 14292 14062 14412 14090
rect 14292 13938 14320 14062
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14278 13832 14334 13841
rect 14278 13767 14334 13776
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14200 13530 14228 13670
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13648 11801 13676 13262
rect 13740 11898 13768 13262
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13634 11792 13690 11801
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13544 11756 13596 11762
rect 13634 11727 13690 11736
rect 13544 11698 13596 11704
rect 13464 11354 13492 11698
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13358 10568 13414 10577
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13280 9926 13308 10542
rect 13464 10538 13492 11290
rect 13358 10503 13414 10512
rect 13452 10532 13504 10538
rect 13372 10130 13400 10503
rect 13452 10474 13504 10480
rect 13556 10418 13584 11698
rect 13740 11558 13768 11834
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13832 11286 13860 11698
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13464 10390 13584 10418
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13268 9920 13320 9926
rect 13174 9888 13230 9897
rect 13268 9862 13320 9868
rect 13174 9823 13230 9832
rect 13188 9489 13216 9823
rect 13174 9480 13230 9489
rect 12530 9415 12586 9424
rect 12716 9444 12768 9450
rect 13174 9415 13230 9424
rect 12716 9386 12768 9392
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12438 9208 12494 9217
rect 12544 9178 12572 9318
rect 12636 9217 12664 9318
rect 12622 9208 12678 9217
rect 12438 9143 12440 9152
rect 12492 9143 12494 9152
rect 12532 9172 12584 9178
rect 12440 9114 12492 9120
rect 12622 9143 12678 9152
rect 12532 9114 12584 9120
rect 12728 8974 12756 9386
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13280 9081 13308 9114
rect 13266 9072 13322 9081
rect 13266 9007 13322 9016
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12176 8758 12296 8786
rect 12176 8548 12204 8758
rect 12176 8520 12296 8548
rect 12084 8452 12204 8480
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11900 7398 12020 7426
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11900 5914 11928 7398
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 6934 12020 7142
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11978 6760 12034 6769
rect 11978 6695 12034 6704
rect 11992 6662 12020 6695
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11716 4706 11744 5578
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11716 4678 11836 4706
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11256 2638 11376 2666
rect 11256 2582 11284 2638
rect 11716 2582 11744 4558
rect 11808 2650 11836 4678
rect 11900 4622 11928 5510
rect 11992 4690 12020 6598
rect 12084 6458 12112 8298
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12084 4826 12112 6122
rect 12176 6118 12204 8452
rect 12268 7478 12296 8520
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 7546 12480 8298
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12544 7342 12572 8434
rect 12728 8090 12756 8910
rect 12992 8900 13044 8906
rect 13044 8860 13216 8888
rect 12992 8842 13044 8848
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12544 7018 12572 7278
rect 12360 7002 12572 7018
rect 12728 7002 12756 7482
rect 13188 7478 13216 8860
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13372 7426 13400 10066
rect 13464 9194 13492 10390
rect 13636 10192 13688 10198
rect 13556 10140 13636 10146
rect 13556 10134 13688 10140
rect 13556 10118 13676 10134
rect 13740 10130 13768 10406
rect 13728 10124 13780 10130
rect 13556 9654 13584 10118
rect 13728 10066 13780 10072
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9722 13676 9998
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13740 9466 13768 9862
rect 13832 9654 13860 11222
rect 13924 11218 13952 12038
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14016 9897 14044 13330
rect 14292 12714 14320 13767
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14108 11898 14136 12242
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14002 9888 14058 9897
rect 14002 9823 14058 9832
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13820 9512 13872 9518
rect 13740 9460 13820 9466
rect 13740 9454 13872 9460
rect 13740 9438 13860 9454
rect 13464 9166 13676 9194
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13648 8242 13676 9166
rect 13740 8362 13768 9438
rect 14016 9330 14044 9658
rect 13832 9302 14044 9330
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13464 7546 13492 8230
rect 13556 7954 13584 8230
rect 13648 8214 13768 8242
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13372 7398 13492 7426
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 12348 6996 12572 7002
rect 12400 6990 12572 6996
rect 12716 6996 12768 7002
rect 12348 6938 12400 6944
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 5642 12204 6054
rect 12268 5914 12296 6734
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6254 12388 6598
rect 12452 6322 12480 6990
rect 12716 6938 12768 6944
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12820 6458 12848 6734
rect 13096 6662 13124 6734
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 13188 6118 13216 7278
rect 13266 7032 13322 7041
rect 13266 6967 13268 6976
rect 13320 6967 13322 6976
rect 13268 6938 13320 6944
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6390 13400 6598
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 13464 5914 13492 7398
rect 13648 7342 13676 8026
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13740 6798 13768 8214
rect 13832 7206 13860 9302
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 13910 8936 13966 8945
rect 13910 8871 13966 8880
rect 13924 7342 13952 8871
rect 14016 8548 14044 9114
rect 14108 9042 14136 9930
rect 14292 9722 14320 12242
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 8650 14136 8978
rect 14108 8622 14320 8650
rect 14188 8560 14240 8566
rect 14016 8520 14136 8548
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12452 5166 12480 5646
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 12254 4584 12310 4593
rect 12254 4519 12310 4528
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12176 4078 12204 4422
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11978 3632 12034 3641
rect 12084 3602 12112 3878
rect 11978 3567 11980 3576
rect 12032 3567 12034 3576
rect 12072 3596 12124 3602
rect 11980 3538 12032 3544
rect 12072 3538 12124 3544
rect 12176 3534 12204 4014
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12084 2990 12112 3062
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 10336 1278 10916 1306
rect 10336 480 10364 1278
rect 11256 480 11284 2314
rect 12176 480 12204 2858
rect 12268 2514 12296 4519
rect 12452 4486 12480 5102
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 12544 4978 12572 5034
rect 12544 4950 12756 4978
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12438 4176 12494 4185
rect 12636 4146 12664 4422
rect 12438 4111 12494 4120
rect 12624 4140 12676 4146
rect 12452 4078 12480 4111
rect 12624 4082 12676 4088
rect 12728 4078 12756 4950
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 13280 4622 13308 5034
rect 13452 4752 13504 4758
rect 13450 4720 13452 4729
rect 13504 4720 13506 4729
rect 13450 4655 13506 4664
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13556 4486 13584 6054
rect 13648 5166 13676 6190
rect 13740 6118 13768 6734
rect 13832 6186 13860 7142
rect 14016 6798 14044 7346
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14016 6458 14044 6734
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 14016 5914 14044 6258
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13740 5370 13768 5714
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13544 4480 13596 4486
rect 13372 4428 13544 4434
rect 13372 4422 13596 4428
rect 13372 4406 13584 4422
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12532 3936 12584 3942
rect 12584 3884 12664 3890
rect 12532 3878 12664 3884
rect 12544 3862 12664 3878
rect 12636 3194 12664 3862
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 13082 3088 13138 3097
rect 13082 3023 13084 3032
rect 13136 3023 13138 3032
rect 13084 2994 13136 3000
rect 12360 2944 12480 2972
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12360 2310 12388 2944
rect 12452 2802 12480 2944
rect 12808 2916 12860 2922
rect 12636 2876 12808 2904
rect 12636 2802 12664 2876
rect 12808 2858 12860 2864
rect 12452 2774 12664 2802
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 13096 480 13124 2382
rect 13372 2106 13400 4406
rect 13648 4298 13676 5102
rect 13556 4270 13676 4298
rect 13556 4078 13584 4270
rect 13636 4208 13688 4214
rect 13740 4196 13768 5306
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13688 4168 13768 4196
rect 13636 4150 13688 4156
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13832 3398 13860 4694
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 4010 14044 4422
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 14004 4004 14056 4010
rect 14004 3946 14056 3952
rect 13924 3466 13952 3946
rect 14108 3738 14136 8520
rect 14188 8502 14240 8508
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13648 3194 13676 3334
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 14016 3058 14044 3538
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 13832 2038 13860 2790
rect 13820 2032 13872 2038
rect 13820 1974 13872 1980
rect 13924 480 13952 2790
rect 14200 2514 14228 8502
rect 14292 4826 14320 8622
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14384 2990 14412 13942
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14554 13424 14610 13433
rect 14464 13388 14516 13394
rect 14554 13359 14610 13368
rect 14464 13330 14516 13336
rect 14476 12850 14504 13330
rect 14568 13258 14596 13359
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14752 13002 14780 13874
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14660 12974 14780 13002
rect 14844 12986 14872 13262
rect 14832 12980 14884 12986
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14476 11898 14504 12378
rect 14568 12306 14596 12922
rect 14660 12782 14688 12974
rect 14832 12922 14884 12928
rect 14648 12776 14700 12782
rect 14740 12776 14792 12782
rect 14648 12718 14700 12724
rect 14738 12744 14740 12753
rect 14792 12744 14794 12753
rect 14660 12442 14688 12718
rect 14738 12679 14794 12688
rect 14844 12594 14872 12922
rect 15106 12880 15162 12889
rect 15106 12815 15162 12824
rect 14752 12566 14872 12594
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14752 12374 14780 12566
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14830 12336 14886 12345
rect 14556 12300 14608 12306
rect 14830 12271 14886 12280
rect 14556 12242 14608 12248
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 11354 14504 11630
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14568 10062 14596 11154
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14476 9382 14504 9658
rect 14660 9518 14688 10406
rect 14648 9512 14700 9518
rect 14554 9480 14610 9489
rect 14700 9460 14780 9466
rect 14648 9454 14780 9460
rect 14660 9438 14780 9454
rect 14554 9415 14610 9424
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14568 9042 14596 9415
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14476 8378 14504 8910
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8498 14596 8774
rect 14660 8498 14688 9318
rect 14752 8974 14780 9438
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14476 8350 14596 8378
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 7002 14504 7142
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14568 6882 14596 8350
rect 14660 8022 14688 8434
rect 14844 8294 14872 12271
rect 15120 11694 15148 12815
rect 15212 11830 15240 14214
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15474 13832 15530 13841
rect 15396 13530 15424 13806
rect 15474 13767 15530 13776
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15304 12442 15332 13194
rect 15382 12744 15438 12753
rect 15382 12679 15438 12688
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15396 12186 15424 12679
rect 15304 12170 15424 12186
rect 15292 12164 15424 12170
rect 15344 12158 15424 12164
rect 15292 12106 15344 12112
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15304 11694 15332 12106
rect 15488 12073 15516 13767
rect 15580 13025 15608 14350
rect 15782 14172 16078 14192
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 16040 13462 16068 13738
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15752 13388 15804 13394
rect 15672 13348 15752 13376
rect 15566 13016 15622 13025
rect 15566 12951 15622 12960
rect 15672 12288 15700 13348
rect 15752 13330 15804 13336
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15842 12880 15898 12889
rect 15842 12815 15898 12824
rect 15936 12844 15988 12850
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15580 12260 15700 12288
rect 15474 12064 15530 12073
rect 15474 11999 15530 12008
rect 15580 11914 15608 12260
rect 15764 12186 15792 12310
rect 15856 12306 15884 12815
rect 15936 12786 15988 12792
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15948 12238 15976 12786
rect 15396 11886 15608 11914
rect 15672 12158 15792 12186
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15108 11688 15160 11694
rect 15292 11688 15344 11694
rect 15108 11630 15160 11636
rect 15198 11656 15254 11665
rect 15292 11630 15344 11636
rect 15198 11591 15254 11600
rect 15212 11234 15240 11591
rect 15120 11206 15240 11234
rect 15120 10606 15148 11206
rect 15304 11150 15332 11630
rect 15292 11144 15344 11150
rect 15198 11112 15254 11121
rect 15292 11086 15344 11092
rect 15198 11047 15254 11056
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14922 9072 14978 9081
rect 14922 9007 14978 9016
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14648 8016 14700 8022
rect 14752 7993 14780 8230
rect 14648 7958 14700 7964
rect 14738 7984 14794 7993
rect 14738 7919 14794 7928
rect 14752 7206 14780 7919
rect 14936 7290 14964 9007
rect 15120 8945 15148 9454
rect 15106 8936 15162 8945
rect 15106 8871 15162 8880
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14844 7262 14964 7290
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14568 6866 14780 6882
rect 14568 6860 14792 6866
rect 14568 6854 14740 6860
rect 14740 6802 14792 6808
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14476 6186 14504 6734
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14476 5914 14504 6122
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14476 4622 14504 5102
rect 14556 4752 14608 4758
rect 14554 4720 14556 4729
rect 14608 4720 14610 4729
rect 14554 4655 14610 4664
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14660 2514 14688 3878
rect 14752 3641 14780 6802
rect 14738 3632 14794 3641
rect 14844 3602 14872 7262
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14738 3567 14794 3576
rect 14832 3596 14884 3602
rect 14752 3466 14780 3567
rect 14832 3538 14884 3544
rect 14740 3460 14792 3466
rect 14740 3402 14792 3408
rect 14936 3058 14964 7142
rect 15028 6304 15056 8366
rect 15120 7528 15148 8774
rect 15212 8514 15240 11047
rect 15304 10606 15332 11086
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 9761 15332 10406
rect 15290 9752 15346 9761
rect 15290 9687 15346 9696
rect 15304 9330 15332 9687
rect 15396 9518 15424 11886
rect 15566 11248 15622 11257
rect 15566 11183 15622 11192
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15488 9926 15516 10542
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15488 9586 15516 9862
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15304 9302 15516 9330
rect 15212 8486 15424 8514
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15212 8090 15240 8366
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15120 7500 15240 7528
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15120 6798 15148 7346
rect 15212 7002 15240 7500
rect 15304 7410 15332 8230
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15108 6316 15160 6322
rect 15028 6276 15108 6304
rect 15108 6258 15160 6264
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 14844 480 14872 2858
rect 15028 2514 15056 4762
rect 15212 3670 15240 6054
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15304 5030 15332 5510
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 15396 2990 15424 8486
rect 15488 5302 15516 9302
rect 15580 6934 15608 11183
rect 15672 9625 15700 12158
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 11257 15976 11630
rect 15934 11248 15990 11257
rect 15934 11183 15990 11192
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 15844 9648 15896 9654
rect 15658 9616 15714 9625
rect 15844 9590 15896 9596
rect 15658 9551 15714 9560
rect 15658 9480 15714 9489
rect 15658 9415 15714 9424
rect 15672 7886 15700 9415
rect 15856 8945 15884 9590
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16040 8974 16068 9522
rect 16028 8968 16080 8974
rect 15842 8936 15898 8945
rect 16028 8910 16080 8916
rect 15842 8871 15898 8880
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15672 7342 15700 7822
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15856 7206 15884 7278
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15672 4826 15700 6598
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 15752 5704 15804 5710
rect 15750 5672 15752 5681
rect 15804 5672 15806 5681
rect 15750 5607 15806 5616
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15750 4992 15806 5001
rect 15750 4927 15806 4936
rect 15764 4826 15792 4927
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15672 3602 15700 4762
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 16132 1034 16160 14350
rect 16316 13394 16344 15399
rect 16394 15056 16450 15065
rect 16394 14991 16450 15000
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16224 12850 16252 13262
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 12986 16344 13194
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16302 12472 16358 12481
rect 16302 12407 16358 12416
rect 16316 12374 16344 12407
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16408 12220 16436 14991
rect 16592 13938 16620 16520
rect 17866 16280 17922 16289
rect 17866 16215 17922 16224
rect 17880 14822 17908 16215
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16684 13977 16712 14010
rect 16670 13968 16726 13977
rect 16580 13932 16632 13938
rect 16670 13903 16726 13912
rect 17224 13932 17276 13938
rect 16580 13874 16632 13880
rect 17224 13874 17276 13880
rect 17130 13424 17186 13433
rect 16580 13388 16632 13394
rect 17130 13359 17186 13368
rect 16580 13330 16632 13336
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16500 12424 16528 13126
rect 16592 12986 16620 13330
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16500 12396 16620 12424
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16316 12192 16436 12220
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16224 11121 16252 11222
rect 16210 11112 16266 11121
rect 16210 11047 16266 11056
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16224 10849 16252 10950
rect 16210 10840 16266 10849
rect 16210 10775 16266 10784
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 9897 16252 10406
rect 16210 9888 16266 9897
rect 16210 9823 16266 9832
rect 16224 9722 16252 9823
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16316 9217 16344 12192
rect 16500 10826 16528 12242
rect 16592 11218 16620 12396
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16684 11354 16712 11562
rect 16776 11354 16804 13262
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16408 10810 16620 10826
rect 16396 10804 16620 10810
rect 16448 10798 16620 10804
rect 16396 10746 16448 10752
rect 16394 10704 16450 10713
rect 16394 10639 16450 10648
rect 16408 10441 16436 10639
rect 16592 10554 16620 10798
rect 16500 10526 16620 10554
rect 16394 10432 16450 10441
rect 16394 10367 16450 10376
rect 16408 10198 16436 10367
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16500 9738 16528 10526
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16408 9710 16528 9738
rect 16302 9208 16358 9217
rect 16302 9143 16358 9152
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8566 16252 8774
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16316 8362 16344 8978
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 7410 16252 7686
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16408 7342 16436 9710
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16500 8673 16528 9114
rect 16486 8664 16542 8673
rect 16486 8599 16542 8608
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16500 7410 16528 8366
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16592 6934 16620 10406
rect 16776 10062 16804 10406
rect 16764 10056 16816 10062
rect 16764 9998 16816 10004
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16684 8022 16712 9046
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16670 7032 16726 7041
rect 16776 7002 16804 9862
rect 16868 8090 16896 12650
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16960 11558 16988 12242
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11014 16988 11494
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 17052 10266 17080 12582
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16946 10160 17002 10169
rect 16946 10095 17002 10104
rect 16960 9994 16988 10095
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7342 16896 7686
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16670 6967 16726 6976
rect 16764 6996 16816 7002
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16224 5234 16252 5646
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16224 4622 16252 5170
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16224 4282 16252 4558
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16316 2650 16344 5646
rect 16592 5098 16620 6190
rect 16684 5778 16712 6967
rect 16764 6938 16816 6944
rect 16960 6866 16988 9658
rect 17052 9382 17080 9998
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17144 8378 17172 13359
rect 17052 8362 17172 8378
rect 17040 8356 17172 8362
rect 17092 8350 17172 8356
rect 17040 8298 17092 8304
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17052 6186 17080 8298
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 7818 17172 8230
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16960 5273 16988 5510
rect 16946 5264 17002 5273
rect 16946 5199 17002 5208
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16500 4865 16528 4966
rect 16486 4856 16542 4865
rect 16486 4791 16542 4800
rect 16592 4758 16620 5034
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 17236 4146 17264 13874
rect 17328 11150 17356 14350
rect 17406 11520 17462 11529
rect 17406 11455 17462 11464
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10810 17356 11086
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17328 10470 17356 10746
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 8090 17356 10066
rect 17420 9654 17448 11455
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17420 8838 17448 9386
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17420 5166 17448 7890
rect 17512 6730 17540 14418
rect 17604 13530 17632 14418
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17590 13424 17646 13433
rect 17590 13359 17592 13368
rect 17644 13359 17646 13368
rect 17592 13330 17644 13336
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17604 10606 17632 13194
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17604 6798 17632 10406
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17590 6488 17646 6497
rect 17590 6423 17592 6432
rect 17644 6423 17646 6432
rect 17592 6394 17644 6400
rect 17498 5672 17554 5681
rect 17498 5607 17500 5616
rect 17552 5607 17554 5616
rect 17500 5578 17552 5584
rect 17408 5160 17460 5166
rect 17408 5102 17460 5108
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4457 17632 4966
rect 17590 4448 17646 4457
rect 17590 4383 17646 4392
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 16684 2990 16712 4082
rect 16854 4040 16910 4049
rect 16854 3975 16910 3984
rect 16868 2990 16896 3975
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17604 3641 17632 3878
rect 17590 3632 17646 3641
rect 17590 3567 17646 3576
rect 17696 3516 17724 13806
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17788 13297 17816 13398
rect 17774 13288 17830 13297
rect 17774 13223 17830 13232
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12102 17816 12786
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 11150 17816 12038
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10062 17816 10950
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17788 9042 17816 9590
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17880 8922 17908 14758
rect 17972 13161 18000 16623
rect 18786 16520 18842 17000
rect 18800 14550 18828 16520
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18064 13870 18092 14282
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17958 13152 18014 13161
rect 17958 13087 18014 13096
rect 17972 9722 18000 13087
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17788 8894 17908 8922
rect 17788 8022 17816 8894
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17880 7886 17908 8774
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17788 3738 17816 7822
rect 17972 7698 18000 9318
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17880 7670 18000 7698
rect 17880 6798 17908 7670
rect 18064 7449 18092 8774
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 18156 7002 18184 9998
rect 18326 9072 18382 9081
rect 18326 9007 18382 9016
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18248 8265 18276 8502
rect 18234 8256 18290 8265
rect 18234 8191 18290 8200
rect 18340 8090 18368 9007
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18234 7848 18290 7857
rect 18234 7783 18290 7792
rect 18248 7546 18276 7783
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18234 7032 18290 7041
rect 18144 6996 18196 7002
rect 18234 6967 18290 6976
rect 18144 6938 18196 6944
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 18248 6458 18276 6967
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18050 6080 18106 6089
rect 18050 6015 18106 6024
rect 18064 5914 18092 6015
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 17880 4690 17908 5063
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4865 18276 4966
rect 18234 4856 18290 4865
rect 18234 4791 18290 4800
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 4049 17908 4422
rect 17866 4040 17922 4049
rect 17866 3975 17922 3984
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17604 3488 17724 3516
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 3097 17448 3334
rect 17406 3088 17462 3097
rect 17406 3023 17462 3032
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 15764 1006 16160 1034
rect 15764 480 15792 1006
rect 16684 480 16712 2926
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 17052 2281 17080 2790
rect 17316 2304 17368 2310
rect 17038 2272 17094 2281
rect 17316 2246 17368 2252
rect 17038 2207 17094 2216
rect 17328 1465 17356 2246
rect 17314 1456 17370 1465
rect 17314 1391 17370 1400
rect 17604 480 17632 3488
rect 17776 2848 17828 2854
rect 17880 2825 17908 3878
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17776 2790 17828 2796
rect 17866 2816 17922 2825
rect 17682 2680 17738 2689
rect 17682 2615 17738 2624
rect 17696 2514 17724 2615
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 17788 1057 17816 2790
rect 17866 2751 17922 2760
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17880 1873 17908 2246
rect 17866 1864 17922 1873
rect 17866 1799 17922 1808
rect 17774 1048 17830 1057
rect 17774 983 17830 992
rect 17972 649 18000 3334
rect 18064 2990 18092 3402
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17958 640 18014 649
rect 17958 575 18014 584
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3054 0 3110 480
rect 3974 0 4030 480
rect 4894 0 4950 480
rect 5814 0 5870 480
rect 6734 0 6790 480
rect 7562 0 7618 480
rect 8482 0 8538 480
rect 9402 0 9458 480
rect 10322 0 10378 480
rect 11242 0 11298 480
rect 12162 0 12218 480
rect 13082 0 13138 480
rect 13910 0 13966 480
rect 14830 0 14886 480
rect 15750 0 15806 480
rect 16670 0 16726 480
rect 17590 0 17646 480
rect 18248 241 18276 2790
rect 18524 480 18552 13942
rect 19432 1488 19484 1494
rect 19432 1430 19484 1436
rect 19444 480 19472 1430
rect 18234 232 18290 241
rect 18234 167 18290 176
rect 18510 0 18566 480
rect 19430 0 19486 480
<< via2 >>
rect 9494 16632 9550 16688
rect 2778 15816 2834 15872
rect 2134 15000 2190 15056
rect 1122 13368 1178 13424
rect 1490 11212 1546 11248
rect 1490 11192 1492 11212
rect 1492 11192 1544 11212
rect 1544 11192 1546 11212
rect 1490 7792 1546 7848
rect 2226 13232 2282 13288
rect 2594 12824 2650 12880
rect 2594 10920 2650 10976
rect 2134 9560 2190 9616
rect 3698 16224 3754 16280
rect 4066 15428 4122 15464
rect 4066 15408 4068 15428
rect 4068 15408 4120 15428
rect 4120 15408 4122 15428
rect 3238 14184 3294 14240
rect 3146 11328 3202 11384
rect 2778 10104 2834 10160
rect 2226 8880 2282 8936
rect 1674 8472 1730 8528
rect 1674 4256 1730 4312
rect 1582 3848 1638 3904
rect 1674 3440 1730 3496
rect 2962 8336 3018 8392
rect 2778 6296 2834 6352
rect 4342 14592 4398 14648
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 3698 13776 3754 13832
rect 3698 12960 3754 13016
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3606 11736 3662 11792
rect 3054 7520 3110 7576
rect 2502 5616 2558 5672
rect 2778 6196 2780 6216
rect 2780 6196 2832 6216
rect 2832 6196 2834 6216
rect 2778 6160 2834 6196
rect 3330 9696 3386 9752
rect 4158 12144 4214 12200
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3882 11736 3938 11792
rect 3514 10512 3570 10568
rect 3422 9288 3478 9344
rect 3330 9036 3386 9072
rect 3330 9016 3332 9036
rect 3332 9016 3384 9036
rect 3384 9016 3386 9036
rect 3422 8336 3478 8392
rect 3238 6704 3294 6760
rect 2962 4664 3018 4720
rect 3054 2796 3056 2816
rect 3056 2796 3108 2816
rect 3108 2796 3110 2816
rect 3054 2760 3110 2796
rect 3606 8880 3662 8936
rect 3606 8200 3662 8256
rect 3606 8064 3662 8120
rect 3514 5208 3570 5264
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 4066 10548 4068 10568
rect 4068 10548 4120 10568
rect 4120 10548 4122 10568
rect 4066 10512 4122 10548
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 4158 8880 4214 8936
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 4066 7928 4122 7984
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 4158 7384 4214 7440
rect 4710 12144 4766 12200
rect 4526 9016 4582 9072
rect 4434 8880 4490 8936
rect 5170 12960 5226 13016
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 6090 13776 6146 13832
rect 5446 11600 5502 11656
rect 4894 9696 4950 9752
rect 5170 10104 5226 10160
rect 4986 9560 5042 9616
rect 4526 8472 4582 8528
rect 4342 7112 4398 7168
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3790 5888 3846 5944
rect 3698 5480 3754 5536
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 4802 8064 4858 8120
rect 4526 7384 4582 7440
rect 4526 6976 4582 7032
rect 4526 6160 4582 6216
rect 4618 5908 4674 5944
rect 4618 5888 4620 5908
rect 4620 5888 4672 5908
rect 4672 5888 4674 5908
rect 3422 3032 3478 3088
rect 3422 2896 3478 2952
rect 3238 1844 3240 1864
rect 3240 1844 3292 1864
rect 3292 1844 3294 1864
rect 3238 1808 3294 1844
rect 4434 5228 4490 5264
rect 4434 5208 4436 5228
rect 4436 5208 4488 5228
rect 4488 5208 4490 5228
rect 5078 6976 5134 7032
rect 4250 5092 4306 5128
rect 4250 5072 4252 5092
rect 4252 5072 4304 5092
rect 4304 5072 4306 5092
rect 4802 5072 4858 5128
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3698 2488 3754 2544
rect 3514 992 3570 1048
rect 4894 4936 4950 4992
rect 5262 5772 5318 5808
rect 5262 5752 5264 5772
rect 5264 5752 5316 5772
rect 5316 5752 5318 5772
rect 5078 2644 5134 2680
rect 5078 2624 5080 2644
rect 5080 2624 5132 2644
rect 5132 2624 5134 2644
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 5630 9968 5686 10024
rect 5814 10784 5870 10840
rect 5630 9424 5686 9480
rect 5630 9152 5686 9208
rect 5814 7792 5870 7848
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 5998 10104 6054 10160
rect 5998 4936 6054 4992
rect 6274 5208 6330 5264
rect 6274 4120 6330 4176
rect 6734 12552 6790 12608
rect 6550 10784 6606 10840
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 7010 11736 7066 11792
rect 7194 11636 7196 11656
rect 7196 11636 7248 11656
rect 7248 11636 7250 11656
rect 7194 11600 7250 11636
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6734 11056 6790 11112
rect 6826 10920 6882 10976
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 7010 9560 7066 9616
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 6550 8200 6606 8256
rect 6918 8356 6974 8392
rect 6918 8336 6920 8356
rect 6920 8336 6972 8356
rect 6972 8336 6974 8356
rect 7470 11600 7526 11656
rect 8114 12824 8170 12880
rect 8114 11192 8170 11248
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6734 7792 6790 7848
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6458 5888 6514 5944
rect 7378 7384 7434 7440
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 7286 5772 7342 5808
rect 7286 5752 7288 5772
rect 7288 5752 7340 5772
rect 7340 5752 7342 5772
rect 6642 5616 6698 5672
rect 7194 5616 7250 5672
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6550 2760 6606 2816
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 7838 9696 7894 9752
rect 7838 8200 7894 8256
rect 8390 11464 8446 11520
rect 8574 11056 8630 11112
rect 8666 10956 8668 10976
rect 8668 10956 8720 10976
rect 8720 10956 8722 10976
rect 8666 10920 8722 10956
rect 8482 9016 8538 9072
rect 8022 8336 8078 8392
rect 8390 8336 8446 8392
rect 7930 7384 7986 7440
rect 8206 5344 8262 5400
rect 8298 5228 8354 5264
rect 8298 5208 8300 5228
rect 8300 5208 8352 5228
rect 8352 5208 8354 5228
rect 17958 16632 18014 16688
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9034 12180 9036 12200
rect 9036 12180 9088 12200
rect 9088 12180 9090 12200
rect 9034 12144 9090 12180
rect 8850 9696 8906 9752
rect 8758 5072 8814 5128
rect 9494 12960 9550 13016
rect 9494 11192 9550 11248
rect 10138 13640 10194 13696
rect 11794 14456 11850 14512
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9402 5208 9458 5264
rect 9218 5108 9220 5128
rect 9220 5108 9272 5128
rect 9272 5108 9274 5128
rect 9218 5072 9274 5108
rect 7378 584 7434 640
rect 8574 1400 8630 1456
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10138 11736 10194 11792
rect 10230 11212 10286 11248
rect 10230 11192 10232 11212
rect 10232 11192 10284 11212
rect 10284 11192 10286 11212
rect 10138 11076 10194 11112
rect 10138 11056 10140 11076
rect 10140 11056 10192 11076
rect 10192 11056 10194 11076
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10322 10920 10378 10976
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10322 9560 10378 9616
rect 9862 9016 9918 9072
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9770 7928 9826 7984
rect 10046 7948 10102 7984
rect 10046 7928 10048 7948
rect 10048 7928 10100 7948
rect 10100 7928 10102 7948
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10046 6704 10102 6760
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10414 9152 10470 9208
rect 11150 13912 11206 13968
rect 10598 9424 10654 9480
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10598 5616 10654 5672
rect 10414 4664 10470 4720
rect 10598 4392 10654 4448
rect 10230 3984 10286 4040
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 10598 3032 10654 3088
rect 11610 13232 11666 13288
rect 11150 9832 11206 9888
rect 11426 12280 11482 12336
rect 11518 12144 11574 12200
rect 11518 11328 11574 11384
rect 11058 4528 11114 4584
rect 11058 4428 11060 4448
rect 11060 4428 11112 4448
rect 11112 4428 11114 4448
rect 11058 4392 11114 4428
rect 11150 4120 11206 4176
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 15566 15816 15622 15872
rect 13542 14320 13598 14376
rect 12346 13676 12348 13696
rect 12348 13676 12400 13696
rect 12400 13676 12402 13696
rect 12346 13640 12402 13676
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 12714 13368 12770 13424
rect 12162 12300 12218 12336
rect 12162 12280 12164 12300
rect 12164 12280 12216 12300
rect 12216 12280 12218 12300
rect 12254 12144 12310 12200
rect 12070 11328 12126 11384
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12622 11600 12678 11656
rect 12806 11600 12862 11656
rect 13174 11600 13230 11656
rect 13266 11500 13268 11520
rect 13268 11500 13320 11520
rect 13320 11500 13322 11520
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12346 9696 12402 9752
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12530 9424 12586 9480
rect 13266 11464 13322 11500
rect 16302 15408 16358 15464
rect 14278 13776 14334 13832
rect 13634 11736 13690 11792
rect 13358 10512 13414 10568
rect 13174 9832 13230 9888
rect 13174 9424 13230 9480
rect 12438 9172 12494 9208
rect 12438 9152 12440 9172
rect 12440 9152 12492 9172
rect 12492 9152 12494 9172
rect 12622 9152 12678 9208
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 13266 9016 13322 9072
rect 11978 6704 12034 6760
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 14002 9832 14058 9888
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 13266 6996 13322 7032
rect 13266 6976 13268 6996
rect 13268 6976 13320 6996
rect 13320 6976 13322 6996
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 13910 8880 13966 8936
rect 12254 4528 12310 4584
rect 11978 3596 12034 3632
rect 11978 3576 11980 3596
rect 11980 3576 12032 3596
rect 12032 3576 12034 3596
rect 12438 4120 12494 4176
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13450 4700 13452 4720
rect 13452 4700 13504 4720
rect 13504 4700 13506 4720
rect 13450 4664 13506 4700
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 13082 3052 13138 3088
rect 13082 3032 13084 3052
rect 13084 3032 13136 3052
rect 13136 3032 13138 3052
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 14554 13368 14610 13424
rect 14738 12724 14740 12744
rect 14740 12724 14792 12744
rect 14792 12724 14794 12744
rect 14738 12688 14794 12724
rect 15106 12824 15162 12880
rect 14830 12280 14886 12336
rect 14554 9424 14610 9480
rect 15474 13776 15530 13832
rect 15382 12688 15438 12744
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15566 12960 15622 13016
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15842 12824 15898 12880
rect 15474 12008 15530 12064
rect 15198 11600 15254 11656
rect 15198 11056 15254 11112
rect 14922 9016 14978 9072
rect 14738 7928 14794 7984
rect 15106 8880 15162 8936
rect 14554 4700 14556 4720
rect 14556 4700 14608 4720
rect 14608 4700 14610 4720
rect 14554 4664 14610 4700
rect 14738 3576 14794 3632
rect 15290 9696 15346 9752
rect 15566 11192 15622 11248
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 15934 11192 15990 11248
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 15658 9560 15714 9616
rect 15658 9424 15714 9480
rect 15842 8880 15898 8936
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 15750 5652 15752 5672
rect 15752 5652 15804 5672
rect 15804 5652 15806 5672
rect 15750 5616 15806 5652
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15750 4936 15806 4992
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 16394 15000 16450 15056
rect 16302 12416 16358 12472
rect 17866 16224 17922 16280
rect 16670 13912 16726 13968
rect 17130 13368 17186 13424
rect 16210 11056 16266 11112
rect 16210 10784 16266 10840
rect 16210 9832 16266 9888
rect 16394 10648 16450 10704
rect 16394 10376 16450 10432
rect 16302 9152 16358 9208
rect 16486 8608 16542 8664
rect 16670 6976 16726 7032
rect 16946 10104 17002 10160
rect 16946 5208 17002 5264
rect 16486 4800 16542 4856
rect 17406 11464 17462 11520
rect 17590 13388 17646 13424
rect 17590 13368 17592 13388
rect 17592 13368 17644 13388
rect 17644 13368 17646 13388
rect 17590 6452 17646 6488
rect 17590 6432 17592 6452
rect 17592 6432 17644 6452
rect 17644 6432 17646 6452
rect 17498 5636 17554 5672
rect 17498 5616 17500 5636
rect 17500 5616 17552 5636
rect 17552 5616 17554 5636
rect 17590 4392 17646 4448
rect 16854 3984 16910 4040
rect 17590 3576 17646 3632
rect 17774 13232 17830 13288
rect 17958 13096 18014 13152
rect 18050 7384 18106 7440
rect 18326 9016 18382 9072
rect 18234 8200 18290 8256
rect 18234 7792 18290 7848
rect 18234 6976 18290 7032
rect 18050 6024 18106 6080
rect 17866 5072 17922 5128
rect 18234 4800 18290 4856
rect 17866 3984 17922 4040
rect 17406 3032 17462 3088
rect 17038 2216 17094 2272
rect 17314 1400 17370 1456
rect 17682 2624 17738 2680
rect 17866 2760 17922 2816
rect 17866 1808 17922 1864
rect 17774 992 17830 1048
rect 17958 584 18014 640
rect 2778 176 2834 232
rect 18234 176 18290 232
<< metal3 >>
rect 0 16690 480 16720
rect 9489 16690 9555 16693
rect 0 16688 9555 16690
rect 0 16632 9494 16688
rect 9550 16632 9555 16688
rect 0 16630 9555 16632
rect 0 16600 480 16630
rect 9489 16627 9555 16630
rect 17953 16690 18019 16693
rect 19520 16690 20000 16720
rect 17953 16688 20000 16690
rect 17953 16632 17958 16688
rect 18014 16632 20000 16688
rect 17953 16630 20000 16632
rect 17953 16627 18019 16630
rect 19520 16600 20000 16630
rect 0 16282 480 16312
rect 3693 16282 3759 16285
rect 0 16280 3759 16282
rect 0 16224 3698 16280
rect 3754 16224 3759 16280
rect 0 16222 3759 16224
rect 0 16192 480 16222
rect 3693 16219 3759 16222
rect 17861 16282 17927 16285
rect 19520 16282 20000 16312
rect 17861 16280 20000 16282
rect 17861 16224 17866 16280
rect 17922 16224 20000 16280
rect 17861 16222 20000 16224
rect 17861 16219 17927 16222
rect 19520 16192 20000 16222
rect 0 15874 480 15904
rect 2773 15874 2839 15877
rect 0 15872 2839 15874
rect 0 15816 2778 15872
rect 2834 15816 2839 15872
rect 0 15814 2839 15816
rect 0 15784 480 15814
rect 2773 15811 2839 15814
rect 15561 15874 15627 15877
rect 19520 15874 20000 15904
rect 15561 15872 20000 15874
rect 15561 15816 15566 15872
rect 15622 15816 20000 15872
rect 15561 15814 20000 15816
rect 15561 15811 15627 15814
rect 19520 15784 20000 15814
rect 0 15466 480 15496
rect 4061 15466 4127 15469
rect 0 15464 4127 15466
rect 0 15408 4066 15464
rect 4122 15408 4127 15464
rect 0 15406 4127 15408
rect 0 15376 480 15406
rect 4061 15403 4127 15406
rect 16297 15466 16363 15469
rect 19520 15466 20000 15496
rect 16297 15464 20000 15466
rect 16297 15408 16302 15464
rect 16358 15408 20000 15464
rect 16297 15406 20000 15408
rect 16297 15403 16363 15406
rect 19520 15376 20000 15406
rect 0 15058 480 15088
rect 2129 15058 2195 15061
rect 0 15056 2195 15058
rect 0 15000 2134 15056
rect 2190 15000 2195 15056
rect 0 14998 2195 15000
rect 0 14968 480 14998
rect 2129 14995 2195 14998
rect 16389 15058 16455 15061
rect 19520 15058 20000 15088
rect 16389 15056 20000 15058
rect 16389 15000 16394 15056
rect 16450 15000 20000 15056
rect 16389 14998 20000 15000
rect 16389 14995 16455 14998
rect 19520 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 480 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 4337 14650 4403 14653
rect 19520 14650 20000 14680
rect 0 14648 4403 14650
rect 0 14592 4342 14648
rect 4398 14592 4403 14648
rect 0 14590 4403 14592
rect 0 14560 480 14590
rect 4337 14587 4403 14590
rect 15886 14590 20000 14650
rect 11789 14514 11855 14517
rect 15886 14514 15946 14590
rect 19520 14560 20000 14590
rect 11789 14512 15946 14514
rect 11789 14456 11794 14512
rect 11850 14456 15946 14512
rect 11789 14454 15946 14456
rect 11789 14451 11855 14454
rect 13537 14378 13603 14381
rect 13537 14376 16268 14378
rect 13537 14320 13542 14376
rect 13598 14320 16268 14376
rect 13537 14318 16268 14320
rect 13537 14315 13603 14318
rect 0 14242 480 14272
rect 3233 14242 3299 14245
rect 0 14240 3299 14242
rect 0 14184 3238 14240
rect 3294 14184 3299 14240
rect 0 14182 3299 14184
rect 16208 14242 16268 14318
rect 19520 14242 20000 14272
rect 16208 14182 20000 14242
rect 0 14152 480 14182
rect 3233 14179 3299 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19520 14152 20000 14182
rect 15770 14111 16090 14112
rect 11145 13970 11211 13973
rect 16665 13970 16731 13973
rect 11145 13968 16731 13970
rect 11145 13912 11150 13968
rect 11206 13912 16670 13968
rect 16726 13912 16731 13968
rect 11145 13910 16731 13912
rect 11145 13907 11211 13910
rect 16665 13907 16731 13910
rect 0 13834 480 13864
rect 3693 13834 3759 13837
rect 0 13832 3759 13834
rect 0 13776 3698 13832
rect 3754 13776 3759 13832
rect 0 13774 3759 13776
rect 0 13744 480 13774
rect 3693 13771 3759 13774
rect 6085 13834 6151 13837
rect 14273 13834 14339 13837
rect 6085 13832 14339 13834
rect 6085 13776 6090 13832
rect 6146 13776 14278 13832
rect 14334 13776 14339 13832
rect 6085 13774 14339 13776
rect 6085 13771 6151 13774
rect 14273 13771 14339 13774
rect 15469 13834 15535 13837
rect 19520 13834 20000 13864
rect 15469 13832 20000 13834
rect 15469 13776 15474 13832
rect 15530 13776 20000 13832
rect 15469 13774 20000 13776
rect 15469 13771 15535 13774
rect 19520 13744 20000 13774
rect 10133 13698 10199 13701
rect 12341 13698 12407 13701
rect 10133 13696 12407 13698
rect 10133 13640 10138 13696
rect 10194 13640 12346 13696
rect 12402 13640 12407 13696
rect 10133 13638 12407 13640
rect 10133 13635 10199 13638
rect 12341 13635 12407 13638
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 0 13426 480 13456
rect 1117 13426 1183 13429
rect 12709 13426 12775 13429
rect 0 13366 1042 13426
rect 0 13336 480 13366
rect 982 13290 1042 13366
rect 1117 13424 12775 13426
rect 1117 13368 1122 13424
rect 1178 13368 12714 13424
rect 12770 13368 12775 13424
rect 1117 13366 12775 13368
rect 1117 13363 1183 13366
rect 12709 13363 12775 13366
rect 14549 13426 14615 13429
rect 17125 13426 17191 13429
rect 17585 13426 17651 13429
rect 14549 13424 17651 13426
rect 14549 13368 14554 13424
rect 14610 13368 17130 13424
rect 17186 13368 17590 13424
rect 17646 13368 17651 13424
rect 14549 13366 17651 13368
rect 14549 13363 14615 13366
rect 17125 13363 17191 13366
rect 17585 13363 17651 13366
rect 2221 13290 2287 13293
rect 982 13288 2287 13290
rect 982 13232 2226 13288
rect 2282 13232 2287 13288
rect 982 13230 2287 13232
rect 2221 13227 2287 13230
rect 11605 13290 11671 13293
rect 17769 13290 17835 13293
rect 19520 13290 20000 13320
rect 11605 13288 16268 13290
rect 11605 13232 11610 13288
rect 11666 13232 16268 13288
rect 11605 13230 16268 13232
rect 11605 13227 11671 13230
rect 16208 13154 16268 13230
rect 17769 13288 20000 13290
rect 17769 13232 17774 13288
rect 17830 13232 20000 13288
rect 17769 13230 20000 13232
rect 17769 13227 17835 13230
rect 19520 13200 20000 13230
rect 17953 13154 18019 13157
rect 16208 13152 18019 13154
rect 16208 13096 17958 13152
rect 18014 13096 18019 13152
rect 16208 13094 18019 13096
rect 17953 13091 18019 13094
rect 3909 13088 4229 13089
rect 0 13018 480 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 13023 16090 13024
rect 3693 13018 3759 13021
rect 0 13016 3759 13018
rect 0 12960 3698 13016
rect 3754 12960 3759 13016
rect 0 12958 3759 12960
rect 0 12928 480 12958
rect 3693 12955 3759 12958
rect 5165 13018 5231 13021
rect 9489 13018 9555 13021
rect 15561 13018 15627 13021
rect 5165 13016 9555 13018
rect 5165 12960 5170 13016
rect 5226 12960 9494 13016
rect 9550 12960 9555 13016
rect 5165 12958 9555 12960
rect 5165 12955 5231 12958
rect 9489 12955 9555 12958
rect 15150 13016 15627 13018
rect 15150 12960 15566 13016
rect 15622 12960 15627 13016
rect 15150 12958 15627 12960
rect 15150 12885 15210 12958
rect 15561 12955 15627 12958
rect 2589 12882 2655 12885
rect 8109 12882 8175 12885
rect 2589 12880 8175 12882
rect 2589 12824 2594 12880
rect 2650 12824 8114 12880
rect 8170 12824 8175 12880
rect 2589 12822 8175 12824
rect 2589 12819 2655 12822
rect 8109 12819 8175 12822
rect 15101 12880 15210 12885
rect 15101 12824 15106 12880
rect 15162 12824 15210 12880
rect 15101 12822 15210 12824
rect 15837 12882 15903 12885
rect 19520 12882 20000 12912
rect 15837 12880 20000 12882
rect 15837 12824 15842 12880
rect 15898 12824 20000 12880
rect 15837 12822 20000 12824
rect 15101 12819 15167 12822
rect 15837 12819 15903 12822
rect 19520 12792 20000 12822
rect 14733 12746 14799 12749
rect 15377 12746 15443 12749
rect 14733 12744 15443 12746
rect 14733 12688 14738 12744
rect 14794 12688 15382 12744
rect 15438 12688 15443 12744
rect 14733 12686 15443 12688
rect 14733 12683 14799 12686
rect 15377 12683 15443 12686
rect 0 12610 480 12640
rect 6729 12610 6795 12613
rect 0 12608 6795 12610
rect 0 12552 6734 12608
rect 6790 12552 6795 12608
rect 0 12550 6795 12552
rect 0 12520 480 12550
rect 6729 12547 6795 12550
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 16297 12474 16363 12477
rect 19520 12474 20000 12504
rect 16297 12472 20000 12474
rect 16297 12416 16302 12472
rect 16358 12416 20000 12472
rect 16297 12414 20000 12416
rect 16297 12411 16363 12414
rect 19520 12384 20000 12414
rect 11421 12338 11487 12341
rect 2776 12336 11487 12338
rect 2776 12304 11426 12336
rect 2638 12280 11426 12304
rect 11482 12280 11487 12336
rect 2638 12278 11487 12280
rect 2638 12244 2836 12278
rect 11421 12275 11487 12278
rect 12157 12338 12223 12341
rect 14825 12338 14891 12341
rect 12157 12336 14891 12338
rect 12157 12280 12162 12336
rect 12218 12280 14830 12336
rect 14886 12280 14891 12336
rect 12157 12278 14891 12280
rect 12157 12275 12223 12278
rect 14825 12275 14891 12278
rect 0 12202 480 12232
rect 2638 12202 2698 12244
rect 0 12142 2698 12202
rect 4153 12202 4219 12205
rect 4705 12202 4771 12205
rect 4153 12200 4771 12202
rect 4153 12144 4158 12200
rect 4214 12144 4710 12200
rect 4766 12144 4771 12200
rect 4153 12142 4771 12144
rect 0 12112 480 12142
rect 4153 12139 4219 12142
rect 4705 12139 4771 12142
rect 9029 12202 9095 12205
rect 11513 12202 11579 12205
rect 12249 12202 12315 12205
rect 9029 12200 10426 12202
rect 9029 12144 9034 12200
rect 9090 12144 10426 12200
rect 9029 12142 10426 12144
rect 9029 12139 9095 12142
rect 10366 12066 10426 12142
rect 11513 12200 16314 12202
rect 11513 12144 11518 12200
rect 11574 12144 12254 12200
rect 12310 12144 16314 12200
rect 11513 12142 16314 12144
rect 11513 12139 11579 12142
rect 12249 12139 12315 12142
rect 15469 12066 15535 12069
rect 10366 12064 15535 12066
rect 10366 12008 15474 12064
rect 15530 12008 15535 12064
rect 10366 12006 15535 12008
rect 16254 12066 16314 12142
rect 19520 12066 20000 12096
rect 16254 12006 20000 12066
rect 15469 12003 15535 12006
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 19520 11976 20000 12006
rect 15770 11935 16090 11936
rect 0 11794 480 11824
rect 3601 11794 3667 11797
rect 0 11792 3667 11794
rect 0 11736 3606 11792
rect 3662 11736 3667 11792
rect 0 11734 3667 11736
rect 0 11704 480 11734
rect 3601 11731 3667 11734
rect 3877 11794 3943 11797
rect 7005 11794 7071 11797
rect 3877 11792 7071 11794
rect 3877 11736 3882 11792
rect 3938 11736 7010 11792
rect 7066 11736 7071 11792
rect 3877 11734 7071 11736
rect 3877 11731 3943 11734
rect 7005 11731 7071 11734
rect 10133 11794 10199 11797
rect 13629 11794 13695 11797
rect 10133 11792 13695 11794
rect 10133 11736 10138 11792
rect 10194 11736 13634 11792
rect 13690 11736 13695 11792
rect 10133 11734 13695 11736
rect 10133 11731 10199 11734
rect 13629 11731 13695 11734
rect 5441 11658 5507 11661
rect 7189 11658 7255 11661
rect 5441 11656 7255 11658
rect 5441 11600 5446 11656
rect 5502 11600 7194 11656
rect 7250 11600 7255 11656
rect 5441 11598 7255 11600
rect 5441 11595 5507 11598
rect 7189 11595 7255 11598
rect 7465 11658 7531 11661
rect 12617 11658 12683 11661
rect 7465 11656 12683 11658
rect 7465 11600 7470 11656
rect 7526 11600 12622 11656
rect 12678 11600 12683 11656
rect 7465 11598 12683 11600
rect 7465 11595 7531 11598
rect 8342 11525 8402 11598
rect 12617 11595 12683 11598
rect 12801 11658 12867 11661
rect 13169 11658 13235 11661
rect 12801 11656 13235 11658
rect 12801 11600 12806 11656
rect 12862 11600 13174 11656
rect 13230 11600 13235 11656
rect 12801 11598 13235 11600
rect 12801 11595 12867 11598
rect 13169 11595 13235 11598
rect 15193 11658 15259 11661
rect 19520 11658 20000 11688
rect 15193 11656 20000 11658
rect 15193 11600 15198 11656
rect 15254 11600 20000 11656
rect 15193 11598 20000 11600
rect 15193 11595 15259 11598
rect 19520 11568 20000 11598
rect 8342 11520 8451 11525
rect 8342 11464 8390 11520
rect 8446 11464 8451 11520
rect 8342 11462 8451 11464
rect 8385 11459 8451 11462
rect 13261 11522 13327 11525
rect 17401 11522 17467 11525
rect 13261 11520 17467 11522
rect 13261 11464 13266 11520
rect 13322 11464 17406 11520
rect 17462 11464 17467 11520
rect 13261 11462 17467 11464
rect 13261 11459 13327 11462
rect 17401 11459 17467 11462
rect 6874 11456 7194 11457
rect 0 11386 480 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 3141 11386 3207 11389
rect 0 11384 3207 11386
rect 0 11328 3146 11384
rect 3202 11328 3207 11384
rect 0 11326 3207 11328
rect 0 11296 480 11326
rect 3141 11323 3207 11326
rect 11513 11386 11579 11389
rect 12065 11386 12131 11389
rect 11513 11384 12131 11386
rect 11513 11328 11518 11384
rect 11574 11328 12070 11384
rect 12126 11328 12131 11384
rect 11513 11326 12131 11328
rect 11513 11323 11579 11326
rect 12065 11323 12131 11326
rect 1485 11250 1551 11253
rect 8109 11250 8175 11253
rect 9489 11250 9555 11253
rect 1485 11248 9555 11250
rect 1485 11192 1490 11248
rect 1546 11192 8114 11248
rect 8170 11192 9494 11248
rect 9550 11192 9555 11248
rect 1485 11190 9555 11192
rect 1485 11187 1551 11190
rect 8109 11187 8175 11190
rect 9489 11187 9555 11190
rect 10225 11250 10291 11253
rect 15561 11250 15627 11253
rect 10225 11248 15627 11250
rect 10225 11192 10230 11248
rect 10286 11192 15566 11248
rect 15622 11192 15627 11248
rect 10225 11190 15627 11192
rect 10225 11187 10291 11190
rect 15561 11187 15627 11190
rect 15929 11250 15995 11253
rect 19520 11250 20000 11280
rect 15929 11248 20000 11250
rect 15929 11192 15934 11248
rect 15990 11192 20000 11248
rect 15929 11190 20000 11192
rect 15929 11187 15995 11190
rect 19520 11160 20000 11190
rect 6729 11114 6795 11117
rect 8569 11114 8635 11117
rect 6729 11112 8635 11114
rect 6729 11056 6734 11112
rect 6790 11056 8574 11112
rect 8630 11056 8635 11112
rect 6729 11054 8635 11056
rect 6729 11051 6795 11054
rect 8569 11051 8635 11054
rect 10133 11114 10199 11117
rect 15193 11114 15259 11117
rect 16205 11114 16271 11117
rect 10133 11112 15259 11114
rect 10133 11056 10138 11112
rect 10194 11056 15198 11112
rect 15254 11056 15259 11112
rect 10133 11054 15259 11056
rect 10133 11051 10199 11054
rect 15193 11051 15259 11054
rect 15564 11112 16271 11114
rect 15564 11056 16210 11112
rect 16266 11056 16271 11112
rect 15564 11054 16271 11056
rect 0 10978 480 11008
rect 2589 10978 2655 10981
rect 0 10976 2655 10978
rect 0 10920 2594 10976
rect 2650 10920 2655 10976
rect 0 10918 2655 10920
rect 0 10888 480 10918
rect 2589 10915 2655 10918
rect 6821 10978 6887 10981
rect 8661 10978 8727 10981
rect 6821 10976 8727 10978
rect 6821 10920 6826 10976
rect 6882 10920 8666 10976
rect 8722 10920 8727 10976
rect 6821 10918 8727 10920
rect 6821 10915 6887 10918
rect 8661 10915 8727 10918
rect 10317 10978 10383 10981
rect 15564 10978 15624 11054
rect 16205 11051 16271 11054
rect 10317 10976 15624 10978
rect 10317 10920 10322 10976
rect 10378 10920 15624 10976
rect 10317 10918 15624 10920
rect 10317 10915 10383 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 5809 10842 5875 10845
rect 6545 10842 6611 10845
rect 16205 10842 16271 10845
rect 19520 10842 20000 10872
rect 5809 10840 6746 10842
rect 5809 10784 5814 10840
rect 5870 10784 6550 10840
rect 6606 10784 6746 10840
rect 5809 10782 6746 10784
rect 5809 10779 5875 10782
rect 6545 10779 6611 10782
rect 6686 10706 6746 10782
rect 16205 10840 20000 10842
rect 16205 10784 16210 10840
rect 16266 10784 20000 10840
rect 16205 10782 20000 10784
rect 16205 10779 16271 10782
rect 19520 10752 20000 10782
rect 16389 10706 16455 10709
rect 6686 10704 16455 10706
rect 6686 10648 16394 10704
rect 16450 10648 16455 10704
rect 6686 10646 16455 10648
rect 16389 10643 16455 10646
rect 0 10570 480 10600
rect 3509 10570 3575 10573
rect 0 10568 3575 10570
rect 0 10512 3514 10568
rect 3570 10512 3575 10568
rect 0 10510 3575 10512
rect 0 10480 480 10510
rect 3509 10507 3575 10510
rect 4061 10570 4127 10573
rect 13353 10570 13419 10573
rect 4061 10568 13419 10570
rect 4061 10512 4066 10568
rect 4122 10512 13358 10568
rect 13414 10512 13419 10568
rect 4061 10510 13419 10512
rect 4061 10507 4127 10510
rect 13353 10507 13419 10510
rect 16389 10434 16455 10437
rect 19520 10434 20000 10464
rect 16389 10432 20000 10434
rect 16389 10376 16394 10432
rect 16450 10376 20000 10432
rect 16389 10374 20000 10376
rect 16389 10371 16455 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19520 10344 20000 10374
rect 12805 10303 13125 10304
rect 0 10162 480 10192
rect 2773 10162 2839 10165
rect 0 10160 2839 10162
rect 0 10104 2778 10160
rect 2834 10104 2839 10160
rect 0 10102 2839 10104
rect 0 10072 480 10102
rect 2773 10099 2839 10102
rect 5165 10162 5231 10165
rect 5993 10162 6059 10165
rect 16941 10162 17007 10165
rect 17718 10162 17724 10164
rect 5165 10160 17724 10162
rect 5165 10104 5170 10160
rect 5226 10104 5998 10160
rect 6054 10104 16946 10160
rect 17002 10104 17724 10160
rect 5165 10102 17724 10104
rect 5165 10099 5231 10102
rect 5993 10099 6059 10102
rect 16941 10099 17007 10102
rect 17718 10100 17724 10102
rect 17788 10100 17794 10164
rect 5625 10026 5691 10029
rect 3328 10024 5691 10026
rect 3328 9968 5630 10024
rect 5686 9968 5691 10024
rect 3328 9966 5691 9968
rect 0 9754 480 9784
rect 3328 9757 3388 9966
rect 5625 9963 5691 9966
rect 11145 9890 11211 9893
rect 13169 9890 13235 9893
rect 13997 9890 14063 9893
rect 11145 9888 14063 9890
rect 11145 9832 11150 9888
rect 11206 9832 13174 9888
rect 13230 9832 14002 9888
rect 14058 9832 14063 9888
rect 11145 9830 14063 9832
rect 11145 9827 11211 9830
rect 13169 9827 13235 9830
rect 13997 9827 14063 9830
rect 16205 9890 16271 9893
rect 19520 9890 20000 9920
rect 16205 9888 20000 9890
rect 16205 9832 16210 9888
rect 16266 9832 20000 9888
rect 16205 9830 20000 9832
rect 16205 9827 16271 9830
rect 3909 9824 4229 9825
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 19520 9800 20000 9830
rect 15770 9759 16090 9760
rect 3325 9754 3391 9757
rect 0 9752 3391 9754
rect 0 9696 3330 9752
rect 3386 9696 3391 9752
rect 0 9694 3391 9696
rect 0 9664 480 9694
rect 3325 9691 3391 9694
rect 4889 9754 4955 9757
rect 7833 9754 7899 9757
rect 8845 9754 8911 9757
rect 4889 9752 8911 9754
rect 4889 9696 4894 9752
rect 4950 9696 7838 9752
rect 7894 9696 8850 9752
rect 8906 9696 8911 9752
rect 4889 9694 8911 9696
rect 4889 9691 4955 9694
rect 7833 9691 7899 9694
rect 8845 9691 8911 9694
rect 12341 9754 12407 9757
rect 15285 9754 15351 9757
rect 12341 9752 15351 9754
rect 12341 9696 12346 9752
rect 12402 9696 15290 9752
rect 15346 9696 15351 9752
rect 12341 9694 15351 9696
rect 12341 9691 12407 9694
rect 15285 9691 15351 9694
rect 2129 9618 2195 9621
rect 4981 9618 5047 9621
rect 2129 9616 5047 9618
rect 2129 9560 2134 9616
rect 2190 9560 4986 9616
rect 5042 9560 5047 9616
rect 2129 9558 5047 9560
rect 2129 9555 2195 9558
rect 4981 9555 5047 9558
rect 6678 9556 6684 9620
rect 6748 9618 6754 9620
rect 7005 9618 7071 9621
rect 6748 9616 7071 9618
rect 6748 9560 7010 9616
rect 7066 9560 7071 9616
rect 6748 9558 7071 9560
rect 6748 9556 6754 9558
rect 7005 9555 7071 9558
rect 10317 9618 10383 9621
rect 15653 9618 15719 9621
rect 10317 9616 15719 9618
rect 10317 9560 10322 9616
rect 10378 9560 15658 9616
rect 15714 9560 15719 9616
rect 10317 9558 15719 9560
rect 10317 9555 10383 9558
rect 15653 9555 15719 9558
rect 5625 9482 5691 9485
rect 10593 9482 10659 9485
rect 12525 9484 12591 9485
rect 12525 9482 12572 9484
rect 5625 9480 10659 9482
rect 5625 9424 5630 9480
rect 5686 9424 10598 9480
rect 10654 9424 10659 9480
rect 5625 9422 10659 9424
rect 12480 9480 12572 9482
rect 12480 9424 12530 9480
rect 12480 9422 12572 9424
rect 5625 9419 5691 9422
rect 10593 9419 10659 9422
rect 12525 9420 12572 9422
rect 12636 9420 12642 9484
rect 13169 9482 13235 9485
rect 14549 9482 14615 9485
rect 13169 9480 14615 9482
rect 13169 9424 13174 9480
rect 13230 9424 14554 9480
rect 14610 9424 14615 9480
rect 13169 9422 14615 9424
rect 12525 9419 12591 9420
rect 13169 9419 13235 9422
rect 14549 9419 14615 9422
rect 15653 9482 15719 9485
rect 19520 9482 20000 9512
rect 15653 9480 20000 9482
rect 15653 9424 15658 9480
rect 15714 9424 20000 9480
rect 15653 9422 20000 9424
rect 15653 9419 15719 9422
rect 19520 9392 20000 9422
rect 0 9346 480 9376
rect 3417 9346 3483 9349
rect 0 9344 3483 9346
rect 0 9288 3422 9344
rect 3478 9288 3483 9344
rect 0 9286 3483 9288
rect 0 9256 480 9286
rect 3417 9283 3483 9286
rect 3420 9210 3480 9283
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 9215 13125 9216
rect 5625 9210 5691 9213
rect 10409 9210 10475 9213
rect 12433 9210 12499 9213
rect 12617 9210 12683 9213
rect 16297 9212 16363 9213
rect 3420 9208 6746 9210
rect 3420 9152 5630 9208
rect 5686 9152 6746 9208
rect 3420 9150 6746 9152
rect 5625 9147 5691 9150
rect 3325 9076 3391 9077
rect 3325 9074 3372 9076
rect 3280 9072 3372 9074
rect 3280 9016 3330 9072
rect 3280 9014 3372 9016
rect 3325 9012 3372 9014
rect 3436 9012 3442 9076
rect 4521 9074 4587 9077
rect 6686 9074 6746 9150
rect 10409 9208 12683 9210
rect 10409 9152 10414 9208
rect 10470 9152 12438 9208
rect 12494 9152 12622 9208
rect 12678 9152 12683 9208
rect 10409 9150 12683 9152
rect 10409 9147 10475 9150
rect 12433 9147 12499 9150
rect 12617 9147 12683 9150
rect 16246 9148 16252 9212
rect 16316 9210 16363 9212
rect 16316 9208 16408 9210
rect 16358 9152 16408 9208
rect 16316 9150 16408 9152
rect 16316 9148 16363 9150
rect 16297 9147 16363 9148
rect 8477 9074 8543 9077
rect 4521 9072 4722 9074
rect 4521 9016 4526 9072
rect 4582 9016 4722 9072
rect 4521 9014 4722 9016
rect 6686 9072 8543 9074
rect 6686 9016 8482 9072
rect 8538 9016 8543 9072
rect 6686 9014 8543 9016
rect 3325 9011 3391 9012
rect 4521 9011 4587 9014
rect 0 8938 480 8968
rect 2221 8938 2287 8941
rect 3601 8938 3667 8941
rect 0 8936 3667 8938
rect 0 8880 2226 8936
rect 2282 8880 3606 8936
rect 3662 8880 3667 8936
rect 0 8878 3667 8880
rect 0 8848 480 8878
rect 2221 8875 2287 8878
rect 3601 8875 3667 8878
rect 4153 8938 4219 8941
rect 4429 8938 4495 8941
rect 4153 8936 4495 8938
rect 4153 8880 4158 8936
rect 4214 8880 4434 8936
rect 4490 8880 4495 8936
rect 4153 8878 4495 8880
rect 4662 8938 4722 9014
rect 8477 9011 8543 9014
rect 9857 9074 9923 9077
rect 13261 9074 13327 9077
rect 14917 9074 14983 9077
rect 18321 9074 18387 9077
rect 19520 9074 20000 9104
rect 9857 9072 20000 9074
rect 9857 9016 9862 9072
rect 9918 9016 13266 9072
rect 13322 9016 14922 9072
rect 14978 9016 18326 9072
rect 18382 9016 20000 9072
rect 9857 9014 20000 9016
rect 9857 9011 9923 9014
rect 13261 9011 13327 9014
rect 14917 9011 14983 9014
rect 18321 9011 18387 9014
rect 19520 8984 20000 9014
rect 13905 8938 13971 8941
rect 15101 8938 15167 8941
rect 4662 8936 15167 8938
rect 4662 8880 13910 8936
rect 13966 8880 15106 8936
rect 15162 8880 15167 8936
rect 4662 8878 15167 8880
rect 4153 8875 4219 8878
rect 4429 8875 4495 8878
rect 13905 8875 13971 8878
rect 15101 8875 15167 8878
rect 15510 8876 15516 8940
rect 15580 8938 15586 8940
rect 15837 8938 15903 8941
rect 15580 8936 15903 8938
rect 15580 8880 15842 8936
rect 15898 8880 15903 8936
rect 15580 8878 15903 8880
rect 15580 8876 15586 8878
rect 15837 8875 15903 8878
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 16481 8666 16547 8669
rect 19520 8666 20000 8696
rect 16481 8664 20000 8666
rect 16481 8608 16486 8664
rect 16542 8608 20000 8664
rect 16481 8606 20000 8608
rect 16481 8603 16547 8606
rect 19520 8576 20000 8606
rect 1669 8530 1735 8533
rect 4521 8530 4587 8533
rect 1669 8528 4587 8530
rect 1669 8472 1674 8528
rect 1730 8472 4526 8528
rect 4582 8472 4587 8528
rect 1669 8470 4587 8472
rect 1669 8467 1735 8470
rect 4521 8467 4587 8470
rect 0 8394 480 8424
rect 2957 8394 3023 8397
rect 0 8392 3023 8394
rect 0 8336 2962 8392
rect 3018 8336 3023 8392
rect 0 8334 3023 8336
rect 0 8304 480 8334
rect 2957 8331 3023 8334
rect 3417 8394 3483 8397
rect 6913 8394 6979 8397
rect 8017 8394 8083 8397
rect 8385 8396 8451 8397
rect 8334 8394 8340 8396
rect 3417 8392 8083 8394
rect 3417 8336 3422 8392
rect 3478 8336 6918 8392
rect 6974 8336 8022 8392
rect 8078 8336 8083 8392
rect 3417 8334 8083 8336
rect 8294 8334 8340 8394
rect 8404 8392 8451 8396
rect 8446 8336 8451 8392
rect 3417 8331 3483 8334
rect 6913 8331 6979 8334
rect 7790 8261 7850 8334
rect 8017 8331 8083 8334
rect 8334 8332 8340 8334
rect 8404 8332 8451 8336
rect 8385 8331 8451 8332
rect 3601 8258 3667 8261
rect 6545 8258 6611 8261
rect 3601 8256 6611 8258
rect 3601 8200 3606 8256
rect 3662 8200 6550 8256
rect 6606 8200 6611 8256
rect 3601 8198 6611 8200
rect 7790 8256 7899 8261
rect 7790 8200 7838 8256
rect 7894 8200 7899 8256
rect 7790 8198 7899 8200
rect 3601 8195 3667 8198
rect 6545 8195 6611 8198
rect 7833 8195 7899 8198
rect 18229 8258 18295 8261
rect 19520 8258 20000 8288
rect 18229 8256 20000 8258
rect 18229 8200 18234 8256
rect 18290 8200 20000 8256
rect 18229 8198 20000 8200
rect 18229 8195 18295 8198
rect 6874 8192 7194 8193
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 19520 8168 20000 8198
rect 12805 8127 13125 8128
rect 3601 8122 3667 8125
rect 4797 8122 4863 8125
rect 3601 8120 4863 8122
rect 3601 8064 3606 8120
rect 3662 8064 4802 8120
rect 4858 8064 4863 8120
rect 3601 8062 4863 8064
rect 3601 8059 3667 8062
rect 4797 8059 4863 8062
rect 0 7986 480 8016
rect 4061 7986 4127 7989
rect 0 7984 4127 7986
rect 0 7928 4066 7984
rect 4122 7928 4127 7984
rect 0 7926 4127 7928
rect 0 7896 480 7926
rect 4061 7923 4127 7926
rect 9765 7986 9831 7989
rect 10041 7986 10107 7989
rect 14733 7986 14799 7989
rect 9765 7984 14799 7986
rect 9765 7928 9770 7984
rect 9826 7928 10046 7984
rect 10102 7928 14738 7984
rect 14794 7928 14799 7984
rect 9765 7926 14799 7928
rect 9765 7923 9831 7926
rect 10041 7923 10107 7926
rect 14733 7923 14799 7926
rect 1485 7850 1551 7853
rect 5809 7850 5875 7853
rect 6729 7852 6795 7853
rect 6678 7850 6684 7852
rect 1485 7848 5875 7850
rect 1485 7792 1490 7848
rect 1546 7792 5814 7848
rect 5870 7792 5875 7848
rect 1485 7790 5875 7792
rect 6638 7790 6684 7850
rect 6748 7848 6795 7852
rect 6790 7792 6795 7848
rect 1485 7787 1551 7790
rect 5809 7787 5875 7790
rect 6678 7788 6684 7790
rect 6748 7788 6795 7792
rect 6729 7787 6795 7788
rect 18229 7850 18295 7853
rect 19520 7850 20000 7880
rect 18229 7848 20000 7850
rect 18229 7792 18234 7848
rect 18290 7792 20000 7848
rect 18229 7790 20000 7792
rect 18229 7787 18295 7790
rect 19520 7760 20000 7790
rect 3909 7648 4229 7649
rect 0 7578 480 7608
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 3049 7578 3115 7581
rect 0 7576 3115 7578
rect 0 7520 3054 7576
rect 3110 7520 3115 7576
rect 0 7518 3115 7520
rect 0 7488 480 7518
rect 3049 7515 3115 7518
rect 4153 7442 4219 7445
rect 4521 7442 4587 7445
rect 4153 7440 4587 7442
rect 4153 7384 4158 7440
rect 4214 7384 4526 7440
rect 4582 7384 4587 7440
rect 4153 7382 4587 7384
rect 4153 7379 4219 7382
rect 4521 7379 4587 7382
rect 7373 7442 7439 7445
rect 7925 7442 7991 7445
rect 7373 7440 7991 7442
rect 7373 7384 7378 7440
rect 7434 7384 7930 7440
rect 7986 7384 7991 7440
rect 7373 7382 7991 7384
rect 7373 7379 7439 7382
rect 7925 7379 7991 7382
rect 18045 7442 18111 7445
rect 19520 7442 20000 7472
rect 18045 7440 20000 7442
rect 18045 7384 18050 7440
rect 18106 7384 20000 7440
rect 18045 7382 20000 7384
rect 18045 7379 18111 7382
rect 19520 7352 20000 7382
rect 0 7170 480 7200
rect 4337 7170 4403 7173
rect 0 7168 4403 7170
rect 0 7112 4342 7168
rect 4398 7112 4403 7168
rect 0 7110 4403 7112
rect 0 7080 480 7110
rect 4337 7107 4403 7110
rect 6874 7104 7194 7105
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 4521 7034 4587 7037
rect 5073 7034 5139 7037
rect 4521 7032 5139 7034
rect 4521 6976 4526 7032
rect 4582 6976 5078 7032
rect 5134 6976 5139 7032
rect 4521 6974 5139 6976
rect 4521 6971 4587 6974
rect 5073 6971 5139 6974
rect 13261 7034 13327 7037
rect 16665 7034 16731 7037
rect 13261 7032 16731 7034
rect 13261 6976 13266 7032
rect 13322 6976 16670 7032
rect 16726 6976 16731 7032
rect 13261 6974 16731 6976
rect 13261 6971 13327 6974
rect 16665 6971 16731 6974
rect 18229 7034 18295 7037
rect 19520 7034 20000 7064
rect 18229 7032 20000 7034
rect 18229 6976 18234 7032
rect 18290 6976 20000 7032
rect 18229 6974 20000 6976
rect 18229 6971 18295 6974
rect 19520 6944 20000 6974
rect 0 6762 480 6792
rect 3233 6762 3299 6765
rect 0 6760 3299 6762
rect 0 6704 3238 6760
rect 3294 6704 3299 6760
rect 0 6702 3299 6704
rect 0 6672 480 6702
rect 3233 6699 3299 6702
rect 10041 6762 10107 6765
rect 11973 6762 12039 6765
rect 10041 6760 12039 6762
rect 10041 6704 10046 6760
rect 10102 6704 11978 6760
rect 12034 6704 12039 6760
rect 10041 6702 12039 6704
rect 10041 6699 10107 6702
rect 11973 6699 12039 6702
rect 3909 6560 4229 6561
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 6495 16090 6496
rect 17585 6490 17651 6493
rect 19520 6490 20000 6520
rect 17585 6488 20000 6490
rect 17585 6432 17590 6488
rect 17646 6432 20000 6488
rect 17585 6430 20000 6432
rect 17585 6427 17651 6430
rect 19520 6400 20000 6430
rect 0 6354 480 6384
rect 2773 6354 2839 6357
rect 0 6352 2839 6354
rect 0 6296 2778 6352
rect 2834 6296 2839 6352
rect 0 6294 2839 6296
rect 0 6264 480 6294
rect 2773 6291 2839 6294
rect 2773 6218 2839 6221
rect 4521 6218 4587 6221
rect 2773 6216 4587 6218
rect 2773 6160 2778 6216
rect 2834 6160 4526 6216
rect 4582 6160 4587 6216
rect 2773 6158 4587 6160
rect 2773 6155 2839 6158
rect 4521 6155 4587 6158
rect 18045 6082 18111 6085
rect 19520 6082 20000 6112
rect 18045 6080 20000 6082
rect 18045 6024 18050 6080
rect 18106 6024 20000 6080
rect 18045 6022 20000 6024
rect 18045 6019 18111 6022
rect 6874 6016 7194 6017
rect 0 5946 480 5976
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 19520 5992 20000 6022
rect 12805 5951 13125 5952
rect 3785 5946 3851 5949
rect 0 5944 3851 5946
rect 0 5888 3790 5944
rect 3846 5888 3851 5944
rect 0 5886 3851 5888
rect 0 5856 480 5886
rect 3785 5883 3851 5886
rect 4613 5946 4679 5949
rect 6453 5946 6519 5949
rect 4613 5944 6519 5946
rect 4613 5888 4618 5944
rect 4674 5888 6458 5944
rect 6514 5888 6519 5944
rect 4613 5886 6519 5888
rect 4613 5883 4679 5886
rect 6453 5883 6519 5886
rect 5257 5810 5323 5813
rect 7281 5810 7347 5813
rect 5257 5808 7347 5810
rect 5257 5752 5262 5808
rect 5318 5752 7286 5808
rect 7342 5752 7347 5808
rect 5257 5750 7347 5752
rect 5257 5747 5323 5750
rect 7281 5747 7347 5750
rect 2497 5674 2563 5677
rect 6637 5674 6703 5677
rect 7189 5674 7255 5677
rect 2497 5672 7255 5674
rect 2497 5616 2502 5672
rect 2558 5616 6642 5672
rect 6698 5616 7194 5672
rect 7250 5616 7255 5672
rect 2497 5614 7255 5616
rect 2497 5611 2563 5614
rect 6637 5611 6703 5614
rect 7189 5611 7255 5614
rect 10593 5674 10659 5677
rect 15745 5674 15811 5677
rect 16246 5674 16252 5676
rect 10593 5672 16252 5674
rect 10593 5616 10598 5672
rect 10654 5616 15750 5672
rect 15806 5616 16252 5672
rect 10593 5614 16252 5616
rect 10593 5611 10659 5614
rect 15745 5611 15811 5614
rect 16246 5612 16252 5614
rect 16316 5612 16322 5676
rect 17493 5674 17559 5677
rect 19520 5674 20000 5704
rect 17493 5672 20000 5674
rect 17493 5616 17498 5672
rect 17554 5616 20000 5672
rect 17493 5614 20000 5616
rect 17493 5611 17559 5614
rect 19520 5584 20000 5614
rect 0 5538 480 5568
rect 3693 5538 3759 5541
rect 0 5536 3759 5538
rect 0 5480 3698 5536
rect 3754 5480 3759 5536
rect 0 5478 3759 5480
rect 0 5448 480 5478
rect 3693 5475 3759 5478
rect 3909 5472 4229 5473
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15770 5407 16090 5408
rect 8201 5402 8267 5405
rect 8334 5402 8340 5404
rect 8201 5400 8340 5402
rect 8201 5344 8206 5400
rect 8262 5344 8340 5400
rect 8201 5342 8340 5344
rect 8201 5339 8267 5342
rect 8334 5340 8340 5342
rect 8404 5340 8410 5404
rect 3509 5266 3575 5269
rect 1534 5264 3575 5266
rect 1534 5208 3514 5264
rect 3570 5208 3575 5264
rect 1534 5206 3575 5208
rect 0 5130 480 5160
rect 1534 5130 1594 5206
rect 3509 5203 3575 5206
rect 4429 5266 4495 5269
rect 6269 5266 6335 5269
rect 4429 5264 6335 5266
rect 4429 5208 4434 5264
rect 4490 5208 6274 5264
rect 6330 5208 6335 5264
rect 4429 5206 6335 5208
rect 4429 5203 4495 5206
rect 6269 5203 6335 5206
rect 8293 5266 8359 5269
rect 9397 5266 9463 5269
rect 8293 5264 9463 5266
rect 8293 5208 8298 5264
rect 8354 5208 9402 5264
rect 9458 5208 9463 5264
rect 8293 5206 9463 5208
rect 8293 5203 8359 5206
rect 9397 5203 9463 5206
rect 16941 5266 17007 5269
rect 19520 5266 20000 5296
rect 16941 5264 20000 5266
rect 16941 5208 16946 5264
rect 17002 5208 20000 5264
rect 16941 5206 20000 5208
rect 16941 5203 17007 5206
rect 19520 5176 20000 5206
rect 0 5070 1594 5130
rect 4245 5130 4311 5133
rect 4797 5130 4863 5133
rect 8753 5130 8819 5133
rect 4245 5128 8819 5130
rect 4245 5072 4250 5128
rect 4306 5072 4802 5128
rect 4858 5072 8758 5128
rect 8814 5072 8819 5128
rect 4245 5070 8819 5072
rect 0 5040 480 5070
rect 4245 5067 4311 5070
rect 4797 5067 4863 5070
rect 8753 5067 8819 5070
rect 9213 5130 9279 5133
rect 17861 5130 17927 5133
rect 9213 5128 17927 5130
rect 9213 5072 9218 5128
rect 9274 5072 17866 5128
rect 17922 5072 17927 5128
rect 9213 5070 17927 5072
rect 9213 5067 9279 5070
rect 17861 5067 17927 5070
rect 4889 4994 4955 4997
rect 5993 4994 6059 4997
rect 4889 4992 6059 4994
rect 4889 4936 4894 4992
rect 4950 4936 5998 4992
rect 6054 4936 6059 4992
rect 4889 4934 6059 4936
rect 4889 4931 4955 4934
rect 5993 4931 6059 4934
rect 15510 4932 15516 4996
rect 15580 4994 15586 4996
rect 15745 4994 15811 4997
rect 15580 4992 15811 4994
rect 15580 4936 15750 4992
rect 15806 4936 15811 4992
rect 15580 4934 15811 4936
rect 15580 4932 15586 4934
rect 15745 4931 15811 4934
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 16481 4858 16547 4861
rect 13310 4856 16547 4858
rect 13310 4800 16486 4856
rect 16542 4800 16547 4856
rect 13310 4798 16547 4800
rect 0 4722 480 4752
rect 2957 4722 3023 4725
rect 0 4720 3023 4722
rect 0 4664 2962 4720
rect 3018 4664 3023 4720
rect 0 4662 3023 4664
rect 0 4632 480 4662
rect 2957 4659 3023 4662
rect 10409 4722 10475 4725
rect 12566 4722 12572 4724
rect 10409 4720 12572 4722
rect 10409 4664 10414 4720
rect 10470 4664 12572 4720
rect 10409 4662 12572 4664
rect 10409 4659 10475 4662
rect 12566 4660 12572 4662
rect 12636 4722 12642 4724
rect 13310 4722 13370 4798
rect 16481 4795 16547 4798
rect 18229 4858 18295 4861
rect 19520 4858 20000 4888
rect 18229 4856 20000 4858
rect 18229 4800 18234 4856
rect 18290 4800 20000 4856
rect 18229 4798 20000 4800
rect 18229 4795 18295 4798
rect 19520 4768 20000 4798
rect 12636 4662 13370 4722
rect 13445 4722 13511 4725
rect 14549 4722 14615 4725
rect 13445 4720 14615 4722
rect 13445 4664 13450 4720
rect 13506 4664 14554 4720
rect 14610 4664 14615 4720
rect 13445 4662 14615 4664
rect 12636 4660 12642 4662
rect 13445 4659 13511 4662
rect 14549 4659 14615 4662
rect 11053 4586 11119 4589
rect 12249 4586 12315 4589
rect 11053 4584 12315 4586
rect 11053 4528 11058 4584
rect 11114 4528 12254 4584
rect 12310 4528 12315 4584
rect 11053 4526 12315 4528
rect 11053 4523 11119 4526
rect 12249 4523 12315 4526
rect 10593 4450 10659 4453
rect 11053 4450 11119 4453
rect 10593 4448 11119 4450
rect 10593 4392 10598 4448
rect 10654 4392 11058 4448
rect 11114 4392 11119 4448
rect 10593 4390 11119 4392
rect 10593 4387 10659 4390
rect 11053 4387 11119 4390
rect 17585 4450 17651 4453
rect 19520 4450 20000 4480
rect 17585 4448 20000 4450
rect 17585 4392 17590 4448
rect 17646 4392 20000 4448
rect 17585 4390 20000 4392
rect 17585 4387 17651 4390
rect 3909 4384 4229 4385
rect 0 4314 480 4344
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 19520 4360 20000 4390
rect 15770 4319 16090 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 480 4254
rect 1669 4251 1735 4254
rect 6269 4178 6335 4181
rect 11145 4178 11211 4181
rect 12433 4178 12499 4181
rect 6269 4176 12499 4178
rect 6269 4120 6274 4176
rect 6330 4120 11150 4176
rect 11206 4120 12438 4176
rect 12494 4120 12499 4176
rect 6269 4118 12499 4120
rect 6269 4115 6335 4118
rect 11145 4115 11211 4118
rect 12433 4115 12499 4118
rect 10225 4042 10291 4045
rect 16849 4042 16915 4045
rect 10225 4040 16915 4042
rect 10225 3984 10230 4040
rect 10286 3984 16854 4040
rect 16910 3984 16915 4040
rect 10225 3982 16915 3984
rect 10225 3979 10291 3982
rect 16849 3979 16915 3982
rect 17861 4042 17927 4045
rect 19520 4042 20000 4072
rect 17861 4040 20000 4042
rect 17861 3984 17866 4040
rect 17922 3984 20000 4040
rect 17861 3982 20000 3984
rect 17861 3979 17927 3982
rect 19520 3952 20000 3982
rect 0 3906 480 3936
rect 1577 3906 1643 3909
rect 0 3904 1643 3906
rect 0 3848 1582 3904
rect 1638 3848 1643 3904
rect 0 3846 1643 3848
rect 0 3816 480 3846
rect 1577 3843 1643 3846
rect 6874 3840 7194 3841
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 11973 3634 12039 3637
rect 14733 3634 14799 3637
rect 11973 3632 14799 3634
rect 11973 3576 11978 3632
rect 12034 3576 14738 3632
rect 14794 3576 14799 3632
rect 11973 3574 14799 3576
rect 11973 3571 12039 3574
rect 14733 3571 14799 3574
rect 17585 3634 17651 3637
rect 19520 3634 20000 3664
rect 17585 3632 20000 3634
rect 17585 3576 17590 3632
rect 17646 3576 20000 3632
rect 17585 3574 20000 3576
rect 17585 3571 17651 3574
rect 19520 3544 20000 3574
rect 0 3498 480 3528
rect 1669 3498 1735 3501
rect 0 3496 1735 3498
rect 0 3440 1674 3496
rect 1730 3440 1735 3496
rect 0 3438 1735 3440
rect 0 3408 480 3438
rect 1669 3435 1735 3438
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 0 3090 480 3120
rect 3417 3090 3483 3093
rect 0 3088 3483 3090
rect 0 3032 3422 3088
rect 3478 3032 3483 3088
rect 0 3030 3483 3032
rect 0 3000 480 3030
rect 3417 3027 3483 3030
rect 10593 3090 10659 3093
rect 13077 3090 13143 3093
rect 10593 3088 13143 3090
rect 10593 3032 10598 3088
rect 10654 3032 13082 3088
rect 13138 3032 13143 3088
rect 10593 3030 13143 3032
rect 10593 3027 10659 3030
rect 13077 3027 13143 3030
rect 17401 3090 17467 3093
rect 19520 3090 20000 3120
rect 17401 3088 20000 3090
rect 17401 3032 17406 3088
rect 17462 3032 20000 3088
rect 17401 3030 20000 3032
rect 17401 3027 17467 3030
rect 19520 3000 20000 3030
rect 3417 2956 3483 2957
rect 3366 2954 3372 2956
rect 3326 2894 3372 2954
rect 3436 2952 3483 2956
rect 3478 2896 3483 2952
rect 3366 2892 3372 2894
rect 3436 2892 3483 2896
rect 3417 2891 3483 2892
rect 3049 2818 3115 2821
rect 6545 2818 6611 2821
rect 3049 2816 6611 2818
rect 3049 2760 3054 2816
rect 3110 2760 6550 2816
rect 6606 2760 6611 2816
rect 3049 2758 6611 2760
rect 3049 2755 3115 2758
rect 6545 2755 6611 2758
rect 17861 2818 17927 2821
rect 17861 2816 17970 2818
rect 17861 2760 17866 2816
rect 17922 2760 17970 2816
rect 17861 2755 17970 2760
rect 6874 2752 7194 2753
rect 0 2682 480 2712
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2687 13125 2688
rect 5073 2682 5139 2685
rect 0 2680 5139 2682
rect 0 2624 5078 2680
rect 5134 2624 5139 2680
rect 0 2622 5139 2624
rect 0 2592 480 2622
rect 5073 2619 5139 2622
rect 17677 2684 17743 2685
rect 17677 2680 17724 2684
rect 17788 2682 17794 2684
rect 17910 2682 17970 2755
rect 19520 2682 20000 2712
rect 17677 2624 17682 2680
rect 17677 2620 17724 2624
rect 17788 2622 17834 2682
rect 17910 2622 20000 2682
rect 17788 2620 17794 2622
rect 17677 2619 17743 2620
rect 19520 2592 20000 2622
rect 3693 2546 3759 2549
rect 3190 2544 3759 2546
rect 3190 2488 3698 2544
rect 3754 2488 3759 2544
rect 3190 2486 3759 2488
rect 0 2274 480 2304
rect 3190 2274 3250 2486
rect 3693 2483 3759 2486
rect 0 2214 3250 2274
rect 17033 2274 17099 2277
rect 19520 2274 20000 2304
rect 17033 2272 20000 2274
rect 17033 2216 17038 2272
rect 17094 2216 20000 2272
rect 17033 2214 20000 2216
rect 0 2184 480 2214
rect 17033 2211 17099 2214
rect 3909 2208 4229 2209
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 19520 2184 20000 2214
rect 15770 2143 16090 2144
rect 0 1866 480 1896
rect 3233 1866 3299 1869
rect 0 1864 3299 1866
rect 0 1808 3238 1864
rect 3294 1808 3299 1864
rect 0 1806 3299 1808
rect 0 1776 480 1806
rect 3233 1803 3299 1806
rect 17861 1866 17927 1869
rect 19520 1866 20000 1896
rect 17861 1864 20000 1866
rect 17861 1808 17866 1864
rect 17922 1808 20000 1864
rect 17861 1806 20000 1808
rect 17861 1803 17927 1806
rect 19520 1776 20000 1806
rect 0 1458 480 1488
rect 8569 1458 8635 1461
rect 0 1456 8635 1458
rect 0 1400 8574 1456
rect 8630 1400 8635 1456
rect 0 1398 8635 1400
rect 0 1368 480 1398
rect 8569 1395 8635 1398
rect 17309 1458 17375 1461
rect 19520 1458 20000 1488
rect 17309 1456 20000 1458
rect 17309 1400 17314 1456
rect 17370 1400 20000 1456
rect 17309 1398 20000 1400
rect 17309 1395 17375 1398
rect 19520 1368 20000 1398
rect 0 1050 480 1080
rect 3509 1050 3575 1053
rect 0 1048 3575 1050
rect 0 992 3514 1048
rect 3570 992 3575 1048
rect 0 990 3575 992
rect 0 960 480 990
rect 3509 987 3575 990
rect 17769 1050 17835 1053
rect 19520 1050 20000 1080
rect 17769 1048 20000 1050
rect 17769 992 17774 1048
rect 17830 992 20000 1048
rect 17769 990 20000 992
rect 17769 987 17835 990
rect 19520 960 20000 990
rect 0 642 480 672
rect 7373 642 7439 645
rect 0 640 7439 642
rect 0 584 7378 640
rect 7434 584 7439 640
rect 0 582 7439 584
rect 0 552 480 582
rect 7373 579 7439 582
rect 17953 642 18019 645
rect 19520 642 20000 672
rect 17953 640 20000 642
rect 17953 584 17958 640
rect 18014 584 20000 640
rect 17953 582 20000 584
rect 17953 579 18019 582
rect 19520 552 20000 582
rect 0 234 480 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 480 174
rect 2773 171 2839 174
rect 18229 234 18295 237
rect 19520 234 20000 264
rect 18229 232 20000 234
rect 18229 176 18234 232
rect 18290 176 20000 232
rect 18229 174 20000 176
rect 18229 171 18295 174
rect 19520 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 17724 10100 17788 10164
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 6684 9556 6748 9620
rect 12572 9480 12636 9484
rect 12572 9424 12586 9480
rect 12586 9424 12636 9480
rect 12572 9420 12636 9424
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 3372 9072 3436 9076
rect 3372 9016 3386 9072
rect 3386 9016 3436 9072
rect 3372 9012 3436 9016
rect 16252 9208 16316 9212
rect 16252 9152 16302 9208
rect 16302 9152 16316 9208
rect 16252 9148 16316 9152
rect 15516 8876 15580 8940
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 8340 8392 8404 8396
rect 8340 8336 8390 8392
rect 8390 8336 8404 8392
rect 8340 8332 8404 8336
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 6684 7848 6748 7852
rect 6684 7792 6734 7848
rect 6734 7792 6748 7848
rect 6684 7788 6748 7792
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 16252 5612 16316 5676
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 8340 5340 8404 5404
rect 15516 4932 15580 4996
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 12572 4660 12636 4724
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 3372 2952 3436 2956
rect 3372 2896 3422 2952
rect 3422 2896 3436 2952
rect 3372 2892 3436 2896
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 17724 2680 17788 2684
rect 17724 2624 17738 2680
rect 17738 2624 17788 2680
rect 17724 2620 17788 2624
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3371 9076 3437 9077
rect 3371 9012 3372 9076
rect 3436 9012 3437 9076
rect 3371 9011 3437 9012
rect 3374 2957 3434 9011
rect 3909 8736 4229 9760
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6683 9620 6749 9621
rect 6683 9556 6684 9620
rect 6748 9556 6749 9620
rect 6683 9555 6749 9556
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 7648 4229 8672
rect 6686 7853 6746 9555
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12571 9484 12637 9485
rect 12571 9420 12572 9484
rect 12636 9420 12637 9484
rect 12571 9419 12637 9420
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 8339 8396 8405 8397
rect 8339 8332 8340 8396
rect 8404 8332 8405 8396
rect 8339 8331 8405 8332
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6683 7852 6749 7853
rect 6683 7788 6684 7852
rect 6748 7788 6749 7852
rect 6683 7787 6749 7788
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3371 2956 3437 2957
rect 3371 2892 3372 2956
rect 3436 2892 3437 2956
rect 3371 2891 3437 2892
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 8342 5405 8402 8331
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 8339 5404 8405 5405
rect 8339 5340 8340 5404
rect 8404 5340 8405 5404
rect 8339 5339 8405 5340
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 4384 10160 5408
rect 12574 4725 12634 9419
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12805 8192 13125 9216
rect 15770 14176 16090 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 15770 13088 16090 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 15770 12000 16090 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 10912 16090 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 9824 16090 10848
rect 17723 10164 17789 10165
rect 17723 10100 17724 10164
rect 17788 10100 17789 10164
rect 17723 10099 17789 10100
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15515 8940 15581 8941
rect 15515 8876 15516 8940
rect 15580 8876 15581 8940
rect 15515 8875 15581 8876
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 4928 13125 5952
rect 15518 4997 15578 8875
rect 15770 8736 16090 9760
rect 16251 9212 16317 9213
rect 16251 9148 16252 9212
rect 16316 9148 16317 9212
rect 16251 9147 16317 9148
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 7648 16090 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 6560 16090 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 15770 5472 16090 6496
rect 16254 5677 16314 9147
rect 16251 5676 16317 5677
rect 16251 5612 16252 5676
rect 16316 5612 16317 5676
rect 16251 5611 16317 5612
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 15515 4996 15581 4997
rect 15515 4932 15516 4996
rect 15580 4932 15581 4996
rect 15515 4931 15581 4932
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12571 4724 12637 4725
rect 12571 4660 12572 4724
rect 12636 4660 12637 4724
rect 12571 4659 12637 4660
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 3840 13125 4864
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15770 4384 16090 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 3296 16090 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 2208 16090 3232
rect 17726 2685 17786 10099
rect 17723 2684 17789 2685
rect 17723 2620 17724 2684
rect 17788 2620 17789 2684
rect 17723 2619 17789 2620
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2128 16090 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8
timestamp 1606821651
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1564 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _49_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1472 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2116 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _32_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4508 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4600 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3864 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1606821651
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1606821651
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1606821651
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_36
timestamp 1606821651
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47
timestamp 1606821651
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46
timestamp 1606821651
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5520 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5612 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1606821651
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1606821651
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1606821651
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 7728 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6992 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7176 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1606821651
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_78
timestamp 1606821651
transform 1 0 8280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1606821651
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 9476 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10304 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606821651
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1606821651
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_89
timestamp 1606821651
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1606821651
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_111
timestamp 1606821651
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109
timestamp 1606821651
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11316 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11592 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1606821651
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13892 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13156 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14444 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1606821651
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1606821651
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1606821651
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606821651
transform 1 0 16100 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15180 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606821651
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1606821651
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_159
timestamp 1606821651
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1606821651
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_168
timestamp 1606821651
transform 1 0 16560 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1606821651
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1606821651
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606821651
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606821651
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1606821651
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1932 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1606821651
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1606821651
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4232 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1606821651
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5244 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 1606821651
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_61
timestamp 1606821651
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6900 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_79
timestamp 1606821651
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10672 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1606821651
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1606821651
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12144 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_113
timestamp 1606821651
transform 1 0 11500 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_119
timestamp 1606821651
transform 1 0 12052 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13800 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_136
timestamp 1606821651
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_147
timestamp 1606821651
transform 1 0 14628 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_166 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 16376 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606821651
transform 1 0 17756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_174
timestamp 1606821651
transform 1 0 17112 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_179
timestamp 1606821651
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1606821651
transform 1 0 18124 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1606821651
transform 1 0 18492 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2576 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1606821651
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606821651
transform 1 0 4232 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_32
timestamp 1606821651
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_38
timestamp 1606821651
transform 1 0 4600 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5888 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1606821651
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1606821651
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_68
timestamp 1606821651
transform 1 0 7360 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1606821651
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 10672 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9752 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1606821651
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_100
timestamp 1606821651
transform 1 0 10304 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1606821651
transform 1 0 12604 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1606821651
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13616 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1606821651
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1606821651
transform 1 0 15088 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_164
timestamp 1606821651
transform 1 0 16192 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1606821651
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_176
timestamp 1606821651
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606821651
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1606821651
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1606821651
transform 1 0 1472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2024 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_8
timestamp 1606821651
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_26
timestamp 1606821651
transform 1 0 3496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1606821651
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 6716 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_48
timestamp 1606821651
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1606821651
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7820 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_70
timestamp 1606821651
transform 1 0 7544 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1606821651
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12604 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 11316 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12328 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_109
timestamp 1606821651
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1606821651
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1606821651
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1606821651
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_163
timestamp 1606821651
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_175
timestamp 1606821651
transform 1 0 17204 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_181
timestamp 1606821651
transform 1 0 17756 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1606821651
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_19
timestamp 1606821651
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 3864 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 4876 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 3036 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606821651
transform 1 0 5888 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_50
timestamp 1606821651
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_56
timestamp 1606821651
transform 1 0 6256 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1606821651
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1606821651
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1606821651
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8832 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1606821651
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_104
timestamp 1606821651
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1606821651
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1606821651
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1606821651
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606821651
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 14352 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1606821651
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_143
timestamp 1606821651
transform 1 0 14260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16008 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_160
timestamp 1606821651
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_171
timestamp 1606821651
transform 1 0 16836 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606821651
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1606821651
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1564 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2392 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_12
timestamp 1606821651
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_28
timestamp 1606821651
transform 1 0 3680 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1606821651
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1606821651
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 3404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3772 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606821651
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_38
timestamp 1606821651
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4140 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4784 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1606821651
transform 1 0 5796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 5520 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 5244 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_42
timestamp 1606821651
transform 1 0 4968 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_49
timestamp 1606821651
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_55
timestamp 1606821651
transform 1 0 6164 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606821651
transform 1 0 8740 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606821651
transform 1 0 7176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7820 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1606821651
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_70
timestamp 1606821651
transform 1 0 7544 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1606821651
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp 1606821651
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9200 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10120 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1606821651
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1606821651
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1606821651
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_104
timestamp 1606821651
transform 1 0 10672 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_114
timestamp 1606821651
transform 1 0 11592 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_122
timestamp 1606821651
transform 1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_110
timestamp 1606821651
transform 1 0 11224 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606821651
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14076 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13064 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1606821651
transform 1 0 14076 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_129
timestamp 1606821651
transform 1 0 12972 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1606821651
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606821651
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_147
timestamp 1606821651
transform 1 0 14628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606821651
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_163
timestamp 1606821651
transform 1 0 16100 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1606821651
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_168
timestamp 1606821651
transform 1 0 16560 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1606821651
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1606821651
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606821651
transform 1 0 16744 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606821651
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_176
timestamp 1606821651
transform 1 0 17296 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_180
timestamp 1606821651
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606821651
transform 1 0 17296 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606821651
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606821651
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_186
timestamp 1606821651
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1606821651
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1606821651
transform 1 0 1656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2300 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_10
timestamp 1606821651
transform 1 0 2024 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1606821651
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1606821651
transform 1 0 5704 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6348 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp 1606821651
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_54
timestamp 1606821651
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7360 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1606821651
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10304 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 9844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1606821651
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_98
timestamp 1606821651
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12328 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 11960 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1606821651
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_121
timestamp 1606821651
transform 1 0 12236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_131
timestamp 1606821651
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_142
timestamp 1606821651
transform 1 0 14168 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1606821651
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1606821651
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1606821651
transform 1 0 17480 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_174
timestamp 1606821651
transform 1 0 17112 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_187
timestamp 1606821651
transform 1 0 18308 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1656 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1606821651
transform 1 0 3312 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 3772 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1606821651
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1606821651
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_38
timestamp 1606821651
transform 1 0 4600 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1606821651
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7176 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_75
timestamp 1606821651
transform 1 0 8004 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_81
timestamp 1606821651
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 10488 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1606821651
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1606821651
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1606821651
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1606821651
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1606821651
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1606821651
transform 1 0 15456 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1606821651
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1606821651
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1606821651
transform 1 0 16468 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_176
timestamp 1606821651
transform 1 0 17296 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606821651
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1606821651
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1606821651
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1606821651
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606821651
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1606821651
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 6164 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_52
timestamp 1606821651
transform 1 0 5888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8096 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 7268 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_64
timestamp 1606821651
transform 1 0 6992 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1606821651
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1606821651
transform 1 0 10856 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1606821651
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606821651
transform 1 0 12972 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 13432 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1606821651
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1606821651
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1606821651
transform 1 0 16284 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1606821651
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 1606821651
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 17296 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_174
timestamp 1606821651
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1606821651
transform 1 0 18124 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1606821651
transform 1 0 18492 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_19
timestamp 1606821651
transform 1 0 2852 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606821651
transform 1 0 4508 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3496 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1606821651
transform 1 0 3404 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1606821651
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_40
timestamp 1606821651
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4968 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_58
timestamp 1606821651
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1606821651
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606821651
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 8464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1606821651
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_83
timestamp 1606821651
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8924 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_105
timestamp 1606821651
transform 1 0 10764 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_132
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1606821651
transform 1 0 13984 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 15088 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1606821651
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16744 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1606821651
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1606821651
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1606821651
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1932 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1606821651
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1606821651
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606821651
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1606821651
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7360 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1606821651
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10120 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1606821651
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1606821651
transform 1 0 10028 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12052 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11040 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp 1606821651
transform 1 0 10948 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1606821651
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13064 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1606821651
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_139
timestamp 1606821651
transform 1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606821651
transform 1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16008 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606821651
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1606821651
transform 1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606821651
transform 1 0 17848 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_178
timestamp 1606821651
transform 1 0 17480 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1606821651
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1606821651
transform 1 0 1656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2300 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_10
timestamp 1606821651
transform 1 0 2024 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1606821651
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606821651
transform 1 0 3956 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606821651
transform 1 0 3036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4692 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1606821651
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_35
timestamp 1606821651
transform 1 0 4324 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1606821651
transform 1 0 3404 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5428 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1606821651
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1606821651
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1606821651
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1606821651
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1606821651
transform 1 0 8556 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606821651
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1606821651
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1606821651
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1606821651
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1606821651
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1606821651
transform 1 0 8832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9476 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10304 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_87
timestamp 1606821651
transform 1 0 9108 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606821651
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1606821651
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606821651
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1606821651
transform 1 0 11132 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1606821651
transform 1 0 11868 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14076 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13984 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1606821651
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 1606821651
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1606821651
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16284 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 1606821651
transform 1 0 15548 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1606821651
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1606821651
transform 1 0 15732 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606821651
transform 1 0 18124 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1606821651
transform 1 0 17112 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606821651
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1606821651
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1606821651
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1606821651
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606821651
transform 1 0 2852 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1840 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_6
timestamp 1606821651
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_17
timestamp 1606821651
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4692 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 3680 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 3404 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1606821651
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_37
timestamp 1606821651
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1606821651
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606821651
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1606821651
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10120 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1606821651
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 11776 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1606821651
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1606821651
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 12696 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_129
timestamp 1606821651
transform 1 0 12972 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16100 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15088 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1606821651
transform 1 0 14720 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1606821651
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1606821651
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_184
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606821651
transform 1 0 1472 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2024 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_8
timestamp 1606821651
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_26
timestamp 1606821651
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1606821651
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1606821651
transform 1 0 6348 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1606821651
transform 1 0 5520 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_56
timestamp 1606821651
transform 1 0 6256 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_66
timestamp 1606821651
transform 1 0 7176 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1606821651
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1606821651
transform 1 0 10120 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1606821651
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11132 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_107
timestamp 1606821651
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1606821651
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606821651
transform 1 0 14444 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 12788 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1606821651
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1606821651
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606821651
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606821651
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_181
timestamp 1606821651
transform 1 0 17756 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1606821651
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2668 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 1656 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1606821651
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 3680 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1606821651
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_44
timestamp 1606821651
transform 1 0 5152 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606821651
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 7544 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 7268 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_66
timestamp 1606821651
transform 1 0 7176 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10304 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_86
timestamp 1606821651
transform 1 0 9016 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_98
timestamp 1606821651
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1606821651
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1606821651
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1606821651
transform 1 0 13064 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1606821651
transform 1 0 14076 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1606821651
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1606821651
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15364 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1606821651
transform 1 0 14904 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_154
timestamp 1606821651
transform 1 0 15272 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1606821651
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_184
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1606821651
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606821651
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1606821651
transform 1 0 5704 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1606821651
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_53
timestamp 1606821651
transform 1 0 5980 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1606821651
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1606821651
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1606821651
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10212 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606821651
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_96
timestamp 1606821651
transform 1 0 9936 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_115
timestamp 1606821651
transform 1 0 11684 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1606821651
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16376 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1606821651
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1606821651
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_163
timestamp 1606821651
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_182
timestamp 1606821651
transform 1 0 17848 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1606821651
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1606821651
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2852 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4784 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1606821651
transform 1 0 4324 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606821651
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5704 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1606821651
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606821651
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1606821651
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1606821651
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8464 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1606821651
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1606821651
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_78
timestamp 1606821651
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1606821651
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1606821651
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1606821651
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_107
timestamp 1606821651
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 10948 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11132 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_124
timestamp 1606821651
transform 1 0 12512 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1606821651
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1606821651
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606821651
transform 1 0 14444 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1606821651
transform 1 0 14168 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_139
timestamp 1606821651
transform 1 0 13892 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1606821651
transform 1 0 13064 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1606821651
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 14904 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16284 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1606821651
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1606821651
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606821651
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606821651
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1606821651
transform 1 0 17296 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1606821651
transform 1 0 16560 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1606821651
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1606821651
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1606821651
transform 1 0 18124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1606821651
transform 1 0 18492 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2024 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1606821651
transform 1 0 1932 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_19
timestamp 1606821651
transform 1 0 2852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 4692 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_27
timestamp 1606821651
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_37
timestamp 1606821651
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1606821651
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606821651
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8096 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1606821651
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1606821651
transform 1 0 8004 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_85
timestamp 1606821651
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1606821651
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_107
timestamp 1606821651
transform 1 0 10948 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1606821651
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12972 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1606821651
transform 1 0 14168 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1606821651
transform 1 0 13800 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15456 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15916 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_21_151
timestamp 1606821651
transform 1 0 14996 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_155
timestamp 1606821651
transform 1 0 15364 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_159
timestamp 1606821651
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606821651
transform 1 0 17296 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_174
timestamp 1606821651
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1606821651
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1606821651
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1748 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_16
timestamp 1606821651
transform 1 0 2576 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4692 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1606821651
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_38
timestamp 1606821651
transform 1 0 4600 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_48
timestamp 1606821651
transform 1 0 5520 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1606821651
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1606821651
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1606821651
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1606821651
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1606821651
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1606821651
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1606821651
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1606821651
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1606821651
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1606821651
transform 1 0 15732 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1606821651
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_156
timestamp 1606821651
transform 1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1606821651
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_172
timestamp 1606821651
transform 1 0 16928 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_183
timestamp 1606821651
transform 1 0 17940 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1606821651
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 1122 16520 1178 17000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal2 s 17590 0 17646 480 6 SC_IN_BOT
port 1 nsew default input
rlabel metal2 s 3330 16520 3386 17000 6 SC_IN_TOP
port 2 nsew default input
rlabel metal2 s 18510 0 18566 480 6 SC_OUT_BOT
port 3 nsew default tristate
rlabel metal2 s 5538 16520 5594 17000 6 SC_OUT_TOP
port 4 nsew default tristate
rlabel metal2 s 1214 0 1270 480 6 bottom_grid_pin_0_
port 5 nsew default tristate
rlabel metal2 s 10322 0 10378 480 6 bottom_grid_pin_10_
port 6 nsew default tristate
rlabel metal2 s 11242 0 11298 480 6 bottom_grid_pin_11_
port 7 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 bottom_grid_pin_12_
port 8 nsew default tristate
rlabel metal2 s 13082 0 13138 480 6 bottom_grid_pin_13_
port 9 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 bottom_grid_pin_14_
port 10 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 bottom_grid_pin_15_
port 11 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 bottom_grid_pin_1_
port 12 nsew default tristate
rlabel metal2 s 3054 0 3110 480 6 bottom_grid_pin_2_
port 13 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 bottom_grid_pin_3_
port 14 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_4_
port 15 nsew default tristate
rlabel metal2 s 5814 0 5870 480 6 bottom_grid_pin_5_
port 16 nsew default tristate
rlabel metal2 s 6734 0 6790 480 6 bottom_grid_pin_6_
port 17 nsew default tristate
rlabel metal2 s 7562 0 7618 480 6 bottom_grid_pin_7_
port 18 nsew default tristate
rlabel metal2 s 8482 0 8538 480 6 bottom_grid_pin_8_
port 19 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 bottom_grid_pin_9_
port 20 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 bottom_width_0_height_0__pin_0_
port 21 nsew default input
rlabel metal2 s 16670 0 16726 480 6 bottom_width_0_height_0__pin_1_lower
port 22 nsew default tristate
rlabel metal2 s 386 0 442 480 6 bottom_width_0_height_0__pin_1_upper
port 23 nsew default tristate
rlabel metal2 s 7746 16520 7802 17000 6 ccff_head
port 24 nsew default input
rlabel metal2 s 9954 16520 10010 17000 6 ccff_tail
port 25 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[0]
port 26 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[10]
port 27 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[11]
port 28 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[12]
port 29 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[13]
port 30 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[14]
port 31 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[15]
port 32 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[16]
port 33 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[17]
port 34 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[18]
port 35 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[19]
port 36 nsew default input
rlabel metal3 s 0 9256 480 9376 6 chanx_left_in[1]
port 37 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[2]
port 38 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[3]
port 39 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[4]
port 40 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[5]
port 41 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[6]
port 42 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[7]
port 43 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[8]
port 44 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[9]
port 45 nsew default input
rlabel metal3 s 0 552 480 672 6 chanx_left_out[0]
port 46 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 chanx_left_out[10]
port 47 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[11]
port 48 nsew default tristate
rlabel metal3 s 0 5448 480 5568 6 chanx_left_out[12]
port 49 nsew default tristate
rlabel metal3 s 0 5856 480 5976 6 chanx_left_out[13]
port 50 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[14]
port 51 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_out[15]
port 52 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 chanx_left_out[16]
port 53 nsew default tristate
rlabel metal3 s 0 7488 480 7608 6 chanx_left_out[17]
port 54 nsew default tristate
rlabel metal3 s 0 7896 480 8016 6 chanx_left_out[18]
port 55 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 chanx_left_out[19]
port 56 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[1]
port 57 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 58 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[3]
port 59 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[4]
port 60 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[5]
port 61 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[6]
port 62 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[7]
port 63 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[8]
port 64 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_out[9]
port 65 nsew default tristate
rlabel metal3 s 19520 8576 20000 8696 6 chanx_right_in[0]
port 66 nsew default input
rlabel metal3 s 19520 12792 20000 12912 6 chanx_right_in[10]
port 67 nsew default input
rlabel metal3 s 19520 13200 20000 13320 6 chanx_right_in[11]
port 68 nsew default input
rlabel metal3 s 19520 13744 20000 13864 6 chanx_right_in[12]
port 69 nsew default input
rlabel metal3 s 19520 14152 20000 14272 6 chanx_right_in[13]
port 70 nsew default input
rlabel metal3 s 19520 14560 20000 14680 6 chanx_right_in[14]
port 71 nsew default input
rlabel metal3 s 19520 14968 20000 15088 6 chanx_right_in[15]
port 72 nsew default input
rlabel metal3 s 19520 15376 20000 15496 6 chanx_right_in[16]
port 73 nsew default input
rlabel metal3 s 19520 15784 20000 15904 6 chanx_right_in[17]
port 74 nsew default input
rlabel metal3 s 19520 16192 20000 16312 6 chanx_right_in[18]
port 75 nsew default input
rlabel metal3 s 19520 16600 20000 16720 6 chanx_right_in[19]
port 76 nsew default input
rlabel metal3 s 19520 8984 20000 9104 6 chanx_right_in[1]
port 77 nsew default input
rlabel metal3 s 19520 9392 20000 9512 6 chanx_right_in[2]
port 78 nsew default input
rlabel metal3 s 19520 9800 20000 9920 6 chanx_right_in[3]
port 79 nsew default input
rlabel metal3 s 19520 10344 20000 10464 6 chanx_right_in[4]
port 80 nsew default input
rlabel metal3 s 19520 10752 20000 10872 6 chanx_right_in[5]
port 81 nsew default input
rlabel metal3 s 19520 11160 20000 11280 6 chanx_right_in[6]
port 82 nsew default input
rlabel metal3 s 19520 11568 20000 11688 6 chanx_right_in[7]
port 83 nsew default input
rlabel metal3 s 19520 11976 20000 12096 6 chanx_right_in[8]
port 84 nsew default input
rlabel metal3 s 19520 12384 20000 12504 6 chanx_right_in[9]
port 85 nsew default input
rlabel metal3 s 19520 144 20000 264 6 chanx_right_out[0]
port 86 nsew default tristate
rlabel metal3 s 19520 4360 20000 4480 6 chanx_right_out[10]
port 87 nsew default tristate
rlabel metal3 s 19520 4768 20000 4888 6 chanx_right_out[11]
port 88 nsew default tristate
rlabel metal3 s 19520 5176 20000 5296 6 chanx_right_out[12]
port 89 nsew default tristate
rlabel metal3 s 19520 5584 20000 5704 6 chanx_right_out[13]
port 90 nsew default tristate
rlabel metal3 s 19520 5992 20000 6112 6 chanx_right_out[14]
port 91 nsew default tristate
rlabel metal3 s 19520 6400 20000 6520 6 chanx_right_out[15]
port 92 nsew default tristate
rlabel metal3 s 19520 6944 20000 7064 6 chanx_right_out[16]
port 93 nsew default tristate
rlabel metal3 s 19520 7352 20000 7472 6 chanx_right_out[17]
port 94 nsew default tristate
rlabel metal3 s 19520 7760 20000 7880 6 chanx_right_out[18]
port 95 nsew default tristate
rlabel metal3 s 19520 8168 20000 8288 6 chanx_right_out[19]
port 96 nsew default tristate
rlabel metal3 s 19520 552 20000 672 6 chanx_right_out[1]
port 97 nsew default tristate
rlabel metal3 s 19520 960 20000 1080 6 chanx_right_out[2]
port 98 nsew default tristate
rlabel metal3 s 19520 1368 20000 1488 6 chanx_right_out[3]
port 99 nsew default tristate
rlabel metal3 s 19520 1776 20000 1896 6 chanx_right_out[4]
port 100 nsew default tristate
rlabel metal3 s 19520 2184 20000 2304 6 chanx_right_out[5]
port 101 nsew default tristate
rlabel metal3 s 19520 2592 20000 2712 6 chanx_right_out[6]
port 102 nsew default tristate
rlabel metal3 s 19520 3000 20000 3120 6 chanx_right_out[7]
port 103 nsew default tristate
rlabel metal3 s 19520 3544 20000 3664 6 chanx_right_out[8]
port 104 nsew default tristate
rlabel metal3 s 19520 3952 20000 4072 6 chanx_right_out[9]
port 105 nsew default tristate
rlabel metal2 s 14370 16520 14426 17000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 106 nsew default tristate
rlabel metal2 s 16578 16520 16634 17000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 107 nsew default input
rlabel metal2 s 18786 16520 18842 17000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 108 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 prog_clk_0_S_in
port 109 nsew default input
rlabel metal3 s 0 144 480 264 6 prog_clk_0_W_out
port 110 nsew default tristate
rlabel metal2 s 12162 16520 12218 17000 6 top_grid_pin_0_
port 111 nsew default tristate
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 112 nsew default input
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 113 nsew default input
<< properties >>
string FIXED_BBOX 0 0 20000 17000
<< end >>
