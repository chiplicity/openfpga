* NGSPICE file created from sb_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt sb_1__2_ SC_IN_BOT SC_OUT_BOT bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ left_top_grid_pin_1_ prog_clk_0_S_in right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ right_top_grid_pin_1_
+ VPWR VGND
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_3.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_062_ chanx_right_in[4] VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
X_114_ chanx_right_in[1] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_0_ bottom_left_grid_pin_46_ chanx_right_in[13] mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_028_ VGND VGND VPWR VPWR _028_/HI _028_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _098_/A sky130_fd_sc_hd__buf_4
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[4] mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_061_ _061_/A VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _061_/A sky130_fd_sc_hd__buf_4
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_113_ chanx_right_in[3] VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_3_ _043_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_mem_bottom_track_1.prog_clk clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ chanx_right_in[2] VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_112_ chanx_right_in[7] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[16] mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xprog_clk_0_FTB00 prog_clk_0_S_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
X_111_ chanx_right_in[11] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ chany_bottom_in[9] chany_bottom_in[2] mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_11.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_11.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_110_ _110_/A VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_11.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__buf_4
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ right_bottom_grid_pin_41_ mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_11.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_13.mux_l2_in_0_ mux_bottom_track_13.mux_l1_in_1_/X mux_bottom_track_13.mux_l1_in_0_/X
+ mux_bottom_track_13.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_13.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_11.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l1_in_0_ right_bottom_grid_pin_37_ right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _110_/A sky130_fd_sc_hd__buf_4
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l2_in_1_ _052_/HI chanx_left_in[18] mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_13.mux_l1_in_1_ _046_/HI chanx_left_in[10] mux_bottom_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_13.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_099_ _099_/A VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_9.mux_l2_in_1_ _029_/HI chanx_left_in[15] mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _093_/A sky130_fd_sc_hd__buf_4
XFILLER_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_6_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.mux_l2_in_3_ _033_/HI left_bottom_grid_pin_40_ mux_left_track_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_13.mux_l1_in_0_ bottom_left_grid_pin_44_ chanx_right_in[10] mux_bottom_track_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l2_in_0_ bottom_left_grid_pin_42_ mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_098_ _098_/A VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.mux_l2_in_0_ chanx_left_in[8] mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l1_in_5_ chany_bottom_in[17] chany_bottom_in[10] mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _059_/A sky130_fd_sc_hd__buf_4
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.mux_l2_in_2_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_4.mux_l2_in_3_ _042_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_097_ _097_/A VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_25.mux_l1_in_0_ chanx_right_in[19] chanx_right_in[18] mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_4_ chany_bottom_in[3] right_bottom_grid_pin_41_ mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[8] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _101_/A sky130_fd_sc_hd__buf_4
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_3.mux_l2_in_1_ left_bottom_grid_pin_34_ chany_bottom_in[14] mux_left_track_3.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_096_ chanx_left_in[18] VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_079_ _079_/A VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_3_ _038_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_3_ right_bottom_grid_pin_40_ right_bottom_grid_pin_39_
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_27.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_095_ chanx_left_in[17] VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_078_ _078_/A VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] chany_bottom_in[15] mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_38_ right_bottom_grid_pin_37_
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_mem_bottom_track_1.prog_clk clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[4] mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_094_ chanx_left_in[16] VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_27_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_077_ _077_/A VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_36_ right_bottom_grid_pin_35_
+ mux_right_track_4.mux_l1_in_6_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_6_/S
+ sky130_fd_sc_hd__dfxtp_1
X_093_ _093_/A VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_21.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_21.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l1_in_3_ _055_/HI chanx_left_in[7] mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_076_ chanx_right_in[18] VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _108_/A sky130_fd_sc_hd__buf_4
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_0_ right_bottom_grid_pin_34_ right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_6_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_38_ right_bottom_grid_pin_34_
+ mux_right_track_16.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__buf_4
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_059_ _059_/A VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ chanx_left_in[14] VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l1_in_2_ chanx_left_in[5] bottom_left_grid_pin_48_ mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_075_ chanx_right_in[17] VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__buf_4
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_058_ _058_/A VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_19.mux_l2_in_0_ mux_bottom_track_19.mux_l1_in_1_/X mux_bottom_track_19.mux_l1_in_0_/X
+ mux_bottom_track_19.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_19.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_21.mux_l2_in_0_ mux_bottom_track_21.mux_l1_in_1_/X mux_bottom_track_21.mux_l1_in_0_/X
+ mux_bottom_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_21.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_27.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_27.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_19.mux_l1_in_1_ _049_/HI chanx_left_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_19.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_21.mux_l1_in_1_ _050_/HI chanx_left_in[16] mux_bottom_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _057_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_091_ chanx_left_in[13] VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ chanx_right_in[16] VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_44_
+ mux_bottom_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_057_ _057_/A VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_27.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_9.mux_l2_in_3_ _036_/HI left_bottom_grid_pin_41_ mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ _109_/A VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_3_ _037_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_19.mux_l1_in_0_ bottom_left_grid_pin_47_ chanx_right_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_21.mux_l1_in_0_ bottom_left_grid_pin_48_ chanx_right_in[16] mux_bottom_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_090_ chanx_left_in[12] VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _099_/A sky130_fd_sc_hd__buf_4
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[5] mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_073_ _073_/A VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_056_ SC_IN_BOT VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_3_ _031_/HI left_bottom_grid_pin_38_ mux_left_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ _108_/A VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l2_in_2_ left_bottom_grid_pin_37_ left_top_grid_pin_1_ mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] chany_bottom_in[19] mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__buf_4
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_072_ chanx_right_in[14] VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_2_ left_bottom_grid_pin_34_ chany_bottom_in[17] mux_left_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_107_ _107_/A VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_9.mux_l2_in_1_ chany_bottom_in[16] chany_bottom_in[9] mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_1_ chany_bottom_in[12] mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[5] right_bottom_grid_pin_41_ mux_right_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_13.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_13.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ chanx_right_in[13] VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.mux_l1_in_3_ _040_/HI chanx_left_in[18] mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_1_ chany_bottom_in[10] chany_bottom_in[3] mux_left_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_106_ _106_/A VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_9.mux_l2_in_0_ chany_bottom_in[2] mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_0.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_13.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_070_ chanx_right_in[12] VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[9] chany_bottom_in[14] mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_19.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_19.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_105_ _105_/A VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chanx_right_in[17] chanx_right_in[8] mux_left_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__buf_4
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l1_in_3_ _044_/HI chanx_left_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l1_in_0_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_35_ right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__buf_4
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_19.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_5.mux_l1_in_6_ left_bottom_grid_pin_41_ left_bottom_grid_pin_40_ mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
X_104_ _104_/A VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_2_ chanx_left_in[1] bottom_left_grid_pin_48_ mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_0_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_15.mux_l2_in_0_ mux_bottom_track_15.mux_l1_in_1_/X mux_bottom_track_15.mux_l1_in_0_/X
+ mux_bottom_track_15.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_39_ right_bottom_grid_pin_35_
+ mux_right_track_24.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_15.mux_l1_in_1_ _047_/HI chanx_left_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_15.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_5.mux_l1_in_5_ left_bottom_grid_pin_39_ left_bottom_grid_pin_38_ mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
X_103_ _103_/A VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_44_
+ mux_bottom_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l2_in_3_ _035_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_15.mux_l1_in_0_ bottom_left_grid_pin_45_ chanx_right_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_27.mux_l2_in_0_ _053_/HI mux_bottom_track_27.mux_l1_in_0_/X mux_bottom_track_27.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_27.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
X_102_ _102_/A VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _097_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_5.mux_l1_in_4_ left_bottom_grid_pin_37_ left_bottom_grid_pin_36_ mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_032_ VGND VGND VPWR VPWR _032_/HI _032_/LO sky130_fd_sc_hd__conb_1
X_101_ _101_/A VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_3_ left_bottom_grid_pin_35_ left_bottom_grid_pin_34_ mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_27.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[15] mux_bottom_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_27.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _065_/A sky130_fd_sc_hd__buf_4
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
X_031_ VGND VGND VPWR VPWR _031_/HI _031_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ _100_/A VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l1_in_3_ _032_/HI left_bottom_grid_pin_39_ mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_1_ chany_bottom_in[15] mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_23.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_23.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_030_ VGND VGND VPWR VPWR _030_/HI _030_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.mux_l1_in_2_ left_bottom_grid_pin_35_ chany_bottom_in[18] mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_33.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l1_in_0_ chanx_right_in[14] chanx_right_in[5] mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_21.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_23.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_11.mux_l3_in_0_ mux_bottom_track_11.mux_l2_in_1_/X mux_bottom_track_11.mux_l2_in_0_/X
+ mux_bottom_track_11.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_089_ _089_/A VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_25.mux_l1_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_11.mux_l2_in_1_ _045_/HI chanx_left_in[19] mux_bottom_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_32.mux_l2_in_1_ _041_/HI chanx_left_in[10] mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_088_ chanx_left_in[10] VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l1_in_0_ chanx_right_in[18] chanx_right_in[9] mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_11.mux_l2_in_0_ chanx_left_in[9] mux_bottom_track_11.mux_l1_in_0_/X
+ mux_bottom_track_11.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_7.mux_l1_in_3_ _028_/HI chanx_left_in[11] mux_bottom_track_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _109_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _106_/A sky130_fd_sc_hd__buf_4
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_7.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_7.mux_l2_in_1_ mux_bottom_track_7.mux_l1_in_3_/X mux_bottom_track_7.mux_l1_in_2_/X
+ mux_bottom_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_087_ chanx_left_in[9] VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _089_/A sky130_fd_sc_hd__buf_4
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l1_in_2_ chanx_left_in[6] bottom_left_grid_pin_49_ mux_bottom_track_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_3_ _030_/HI left_bottom_grid_pin_41_ mux_left_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_11.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[9] mux_bottom_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_mem_bottom_track_1.prog_clk clkbuf_3_7_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_23.mux_l2_in_0_ mux_bottom_track_23.mux_l1_in_1_/X mux_bottom_track_23.mux_l1_in_0_/X
+ mux_bottom_track_23.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_23.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_32.mux_l1_in_0_ right_bottom_grid_pin_40_ right_bottom_grid_pin_36_
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_23.mux_l1_in_1_ _051_/HI chanx_left_in[17] mux_bottom_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_23.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_086_ chanx_left_in[8] VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _058_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_069_ _069_/A VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_7.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_7.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_1.mux_l2_in_2_ left_bottom_grid_pin_39_ left_bottom_grid_pin_37_ mux_left_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_3_ _039_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_23.mux_l1_in_0_ bottom_left_grid_pin_49_ chanx_right_in[17] mux_bottom_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_15.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_15.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ _085_/A VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_068_ chanx_right_in[10] VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _100_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_7.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[6] mux_bottom_track_7.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_1_ left_bottom_grid_pin_35_ left_top_grid_pin_1_ mux_left_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] chany_bottom_in[18] mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_13.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_15.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_084_ chanx_left_in[6] VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_067_ chanx_right_in[9] VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l2_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ chanx_left_in[5] VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_066_ chanx_right_in[8] VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail VGND VGND VPWR VPWR mux_left_track_33.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[2] mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ _034_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_082_ chanx_left_in[4] VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_33.mux_l1_in_2_ left_bottom_grid_pin_40_ left_bottom_grid_pin_36_
+ mux_left_track_33.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_065_ _065_/A VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xclkbuf_3_5_0_mem_bottom_track_1.prog_clk clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
XANTENNA_2 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l1_in_3_ _054_/HI chanx_left_in[4] mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_081_ _081_/A VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l1_in_1_ chany_bottom_in[19] chany_bottom_in[12] mux_left_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_0_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__buf_4
X_064_ chanx_right_in[6] VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_116_ chanx_left_in[0] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l1_in_2_ chanx_left_in[3] bottom_left_grid_pin_49_ mux_bottom_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_080_ chanx_left_in[2] VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l1_in_0_ chany_bottom_in[5] chanx_right_in[10] mux_left_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_063_ chanx_right_in[5] VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_2_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ chanx_right_in[0] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_17.mux_l1_in_1_ _048_/HI chanx_left_in[13] mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_029_ VGND VGND VPWR VPWR _029_/HI _029_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

