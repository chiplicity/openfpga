magic
tech EFS8A
magscale 1 2
timestamp 1603804078
<< locali >>
rect 9505 8415 9539 8585
<< viali >>
rect 8125 37281 8159 37315
rect 10977 36873 11011 36907
rect 6996 36669 7030 36703
rect 8033 36669 8067 36703
rect 8585 36669 8619 36703
rect 10793 36669 10827 36703
rect 7067 36533 7101 36567
rect 7389 36533 7423 36567
rect 7849 36533 7883 36567
rect 8309 36533 8343 36567
rect 11345 36533 11379 36567
rect 9873 36329 9907 36363
rect 11437 36329 11471 36363
rect 7297 36261 7331 36295
rect 9689 36193 9723 36227
rect 11253 36193 11287 36227
rect 7205 36125 7239 36159
rect 7757 36057 7791 36091
rect 8769 35989 8803 36023
rect 8125 35785 8159 35819
rect 10425 35785 10459 35819
rect 11483 35785 11517 35819
rect 12633 35785 12667 35819
rect 7757 35717 7791 35751
rect 7205 35649 7239 35683
rect 8677 35581 8711 35615
rect 9229 35581 9263 35615
rect 10241 35581 10275 35615
rect 10793 35581 10827 35615
rect 11412 35581 11446 35615
rect 12449 35581 12483 35615
rect 6285 35513 6319 35547
rect 7297 35513 7331 35547
rect 6653 35445 6687 35479
rect 8493 35445 8527 35479
rect 8769 35445 8803 35479
rect 9781 35445 9815 35479
rect 11805 35445 11839 35479
rect 12173 35445 12207 35479
rect 13001 35445 13035 35479
rect 7849 35241 7883 35275
rect 11713 35241 11747 35275
rect 12909 35241 12943 35275
rect 7021 35173 7055 35207
rect 9965 35173 9999 35207
rect 5892 35105 5926 35139
rect 8620 35105 8654 35139
rect 11529 35105 11563 35139
rect 12725 35105 12759 35139
rect 6929 35037 6963 35071
rect 7573 35037 7607 35071
rect 8723 35037 8757 35071
rect 9873 35037 9907 35071
rect 10517 35037 10551 35071
rect 5963 34969 5997 35003
rect 6653 34969 6687 35003
rect 5273 34901 5307 34935
rect 10885 34901 10919 34935
rect 4307 34697 4341 34731
rect 6285 34697 6319 34731
rect 7757 34697 7791 34731
rect 8493 34697 8527 34731
rect 13645 34697 13679 34731
rect 8217 34561 8251 34595
rect 8677 34561 8711 34595
rect 10517 34561 10551 34595
rect 10885 34561 10919 34595
rect 12587 34561 12621 34595
rect 4204 34493 4238 34527
rect 4629 34493 4663 34527
rect 5089 34493 5123 34527
rect 5181 34493 5215 34527
rect 5641 34493 5675 34527
rect 5917 34493 5951 34527
rect 6837 34493 6871 34527
rect 9597 34493 9631 34527
rect 9873 34493 9907 34527
rect 11529 34493 11563 34527
rect 12484 34493 12518 34527
rect 12909 34493 12943 34527
rect 13277 34493 13311 34527
rect 13461 34493 13495 34527
rect 14013 34493 14047 34527
rect 7158 34425 7192 34459
rect 9039 34425 9073 34459
rect 10609 34425 10643 34459
rect 6561 34357 6595 34391
rect 10333 34357 10367 34391
rect 7389 34153 7423 34187
rect 9413 34153 9447 34187
rect 10609 34153 10643 34187
rect 13553 34153 13587 34187
rect 6187 34085 6221 34119
rect 7021 34085 7055 34119
rect 7757 34085 7791 34119
rect 10051 34085 10085 34119
rect 11529 34085 11563 34119
rect 11621 34085 11655 34119
rect 4848 34017 4882 34051
rect 6745 34017 6779 34051
rect 13369 34017 13403 34051
rect 5825 33949 5859 33983
rect 7665 33949 7699 33983
rect 7941 33949 7975 33983
rect 9689 33949 9723 33983
rect 11989 33949 12023 33983
rect 4951 33881 4985 33915
rect 5273 33813 5307 33847
rect 5641 33813 5675 33847
rect 8677 33813 8711 33847
rect 10885 33813 10919 33847
rect 12541 33813 12575 33847
rect 4813 33609 4847 33643
rect 7849 33609 7883 33643
rect 8309 33609 8343 33643
rect 10057 33609 10091 33643
rect 10425 33609 10459 33643
rect 11713 33609 11747 33643
rect 9689 33541 9723 33575
rect 5917 33473 5951 33507
rect 6561 33473 6595 33507
rect 7573 33473 7607 33507
rect 8769 33473 8803 33507
rect 10517 33473 10551 33507
rect 12817 33473 12851 33507
rect 3893 33405 3927 33439
rect 4077 33405 4111 33439
rect 5273 33405 5307 33439
rect 5641 33405 5675 33439
rect 3525 33337 3559 33371
rect 6929 33337 6963 33371
rect 7021 33337 7055 33371
rect 8677 33337 8711 33371
rect 9090 33337 9124 33371
rect 10838 33337 10872 33371
rect 12541 33337 12575 33371
rect 12633 33337 12667 33371
rect 3893 33269 3927 33303
rect 6193 33269 6227 33303
rect 11437 33269 11471 33303
rect 12173 33269 12207 33303
rect 13553 33269 13587 33303
rect 3709 33065 3743 33099
rect 4859 33065 4893 33099
rect 5641 33065 5675 33099
rect 8861 33065 8895 33099
rect 9873 33065 9907 33099
rect 11529 33065 11563 33099
rect 6095 32997 6129 33031
rect 8033 32997 8067 33031
rect 10333 32997 10367 33031
rect 10885 32997 10919 33031
rect 11805 32997 11839 33031
rect 11897 32997 11931 33031
rect 4756 32929 4790 32963
rect 13344 32929 13378 32963
rect 5733 32861 5767 32895
rect 7941 32861 7975 32895
rect 8309 32861 8343 32895
rect 10241 32861 10275 32895
rect 12081 32861 12115 32895
rect 5181 32725 5215 32759
rect 6653 32725 6687 32759
rect 7021 32725 7055 32759
rect 7389 32725 7423 32759
rect 13415 32725 13449 32759
rect 4997 32521 5031 32555
rect 8309 32521 8343 32555
rect 8585 32521 8619 32555
rect 10977 32521 11011 32555
rect 11713 32521 11747 32555
rect 12173 32521 12207 32555
rect 12587 32521 12621 32555
rect 6561 32385 6595 32419
rect 9505 32385 9539 32419
rect 10057 32385 10091 32419
rect 10701 32385 10735 32419
rect 4236 32317 4270 32351
rect 4629 32317 4663 32351
rect 5181 32317 5215 32351
rect 5641 32317 5675 32351
rect 7389 32317 7423 32351
rect 12484 32317 12518 32351
rect 12909 32317 12943 32351
rect 5917 32249 5951 32283
rect 7711 32249 7745 32283
rect 9873 32249 9907 32283
rect 10149 32249 10183 32283
rect 4307 32181 4341 32215
rect 6285 32181 6319 32215
rect 7205 32181 7239 32215
rect 11345 32181 11379 32215
rect 13369 32181 13403 32215
rect 6285 31977 6319 32011
rect 7849 31977 7883 32011
rect 8217 31977 8251 32011
rect 8723 31977 8757 32011
rect 9781 31977 9815 32011
rect 11391 31977 11425 32011
rect 6009 31909 6043 31943
rect 7021 31909 7055 31943
rect 7573 31909 7607 31943
rect 4112 31841 4146 31875
rect 5457 31841 5491 31875
rect 5733 31841 5767 31875
rect 8652 31841 8686 31875
rect 9965 31841 9999 31875
rect 10149 31841 10183 31875
rect 11320 31841 11354 31875
rect 4215 31773 4249 31807
rect 6918 31773 6952 31807
rect 9137 31637 9171 31671
rect 10701 31637 10735 31671
rect 5733 31433 5767 31467
rect 6561 31433 6595 31467
rect 7021 31433 7055 31467
rect 8125 31365 8159 31399
rect 7573 31297 7607 31331
rect 9597 31297 9631 31331
rect 10793 31297 10827 31331
rect 11437 31297 11471 31331
rect 4537 31229 4571 31263
rect 5181 31229 5215 31263
rect 9045 31229 9079 31263
rect 9505 31229 9539 31263
rect 4169 31161 4203 31195
rect 7665 31161 7699 31195
rect 10425 31161 10459 31195
rect 10885 31161 10919 31195
rect 4905 31093 4939 31127
rect 6101 31093 6135 31127
rect 8677 31093 8711 31127
rect 10057 31093 10091 31127
rect 11805 31093 11839 31127
rect 9045 30889 9079 30923
rect 10609 30889 10643 30923
rect 10885 30889 10919 30923
rect 4813 30821 4847 30855
rect 7849 30821 7883 30855
rect 10051 30821 10085 30855
rect 11621 30821 11655 30855
rect 6285 30753 6319 30787
rect 6469 30753 6503 30787
rect 4721 30685 4755 30719
rect 5365 30685 5399 30719
rect 7757 30685 7791 30719
rect 9689 30685 9723 30719
rect 11529 30685 11563 30719
rect 11989 30685 12023 30719
rect 8309 30617 8343 30651
rect 8677 30617 8711 30651
rect 5733 30549 5767 30583
rect 6561 30549 6595 30583
rect 7113 30549 7147 30583
rect 7573 30549 7607 30583
rect 4721 30345 4755 30379
rect 6377 30345 6411 30379
rect 7757 30345 7791 30379
rect 8033 30345 8067 30379
rect 11529 30345 11563 30379
rect 3893 30277 3927 30311
rect 8815 30277 8849 30311
rect 10609 30277 10643 30311
rect 11805 30277 11839 30311
rect 3985 30209 4019 30243
rect 5365 30209 5399 30243
rect 9689 30209 9723 30243
rect 6837 30141 6871 30175
rect 8712 30141 8746 30175
rect 5089 30073 5123 30107
rect 5181 30073 5215 30107
rect 7158 30073 7192 30107
rect 9137 30073 9171 30107
rect 9505 30073 9539 30107
rect 10010 30073 10044 30107
rect 8401 30005 8435 30039
rect 10885 30005 10919 30039
rect 4629 29801 4663 29835
rect 7573 29801 7607 29835
rect 7849 29801 7883 29835
rect 8401 29801 8435 29835
rect 9505 29801 9539 29835
rect 11253 29801 11287 29835
rect 12403 29801 12437 29835
rect 4905 29733 4939 29767
rect 6974 29733 7008 29767
rect 9873 29733 9907 29767
rect 3040 29665 3074 29699
rect 12332 29665 12366 29699
rect 4813 29597 4847 29631
rect 6653 29597 6687 29631
rect 9781 29597 9815 29631
rect 10425 29597 10459 29631
rect 5365 29529 5399 29563
rect 3111 29461 3145 29495
rect 5733 29461 5767 29495
rect 6377 29461 6411 29495
rect 10793 29461 10827 29495
rect 13001 29257 13035 29291
rect 6561 29189 6595 29223
rect 4997 29121 5031 29155
rect 5365 29121 5399 29155
rect 7389 29121 7423 29155
rect 10425 29121 10459 29155
rect 10885 29121 10919 29155
rect 3944 29053 3978 29087
rect 4353 29053 4387 29087
rect 6285 29053 6319 29087
rect 7021 29053 7055 29087
rect 7297 29053 7331 29087
rect 8585 29053 8619 29087
rect 9505 29053 9539 29087
rect 12449 29053 12483 29087
rect 13277 29053 13311 29087
rect 13496 29053 13530 29087
rect 13921 29053 13955 29087
rect 3065 28985 3099 29019
rect 4031 28985 4065 29019
rect 5089 28985 5123 29019
rect 8125 28985 8159 29019
rect 8906 28985 8940 29019
rect 9873 28985 9907 29019
rect 10241 28985 10275 29019
rect 10517 28985 10551 29019
rect 13599 28985 13633 29019
rect 4721 28917 4755 28951
rect 8401 28917 8435 28951
rect 12633 28917 12667 28951
rect 4629 28713 4663 28747
rect 6193 28713 6227 28747
rect 9965 28713 9999 28747
rect 4721 28645 4755 28679
rect 7297 28645 7331 28679
rect 8769 28645 8803 28679
rect 10333 28645 10367 28679
rect 11897 28645 11931 28679
rect 4813 28577 4847 28611
rect 5733 28577 5767 28611
rect 6561 28577 6595 28611
rect 6745 28577 6779 28611
rect 8033 28577 8067 28611
rect 8585 28577 8619 28611
rect 10885 28577 10919 28611
rect 13312 28577 13346 28611
rect 6837 28509 6871 28543
rect 10241 28509 10275 28543
rect 11805 28509 11839 28543
rect 12357 28441 12391 28475
rect 13415 28441 13449 28475
rect 4537 28169 4571 28203
rect 5917 28169 5951 28203
rect 9781 28169 9815 28203
rect 11161 28169 11195 28203
rect 11437 28169 11471 28203
rect 11805 28169 11839 28203
rect 13645 28169 13679 28203
rect 3341 28033 3375 28067
rect 4905 28033 4939 28067
rect 7941 28033 7975 28067
rect 13277 28033 13311 28067
rect 3709 27965 3743 27999
rect 3801 27965 3835 27999
rect 4169 27965 4203 27999
rect 4997 27965 5031 27999
rect 7205 27965 7239 27999
rect 7389 27965 7423 27999
rect 7665 27965 7699 27999
rect 8493 27965 8527 27999
rect 10241 27965 10275 27999
rect 12449 27965 12483 27999
rect 12633 27965 12667 27999
rect 5318 27897 5352 27931
rect 6653 27897 6687 27931
rect 8401 27897 8435 27931
rect 8855 27897 8889 27931
rect 10057 27897 10091 27931
rect 10562 27897 10596 27931
rect 6285 27829 6319 27863
rect 9413 27829 9447 27863
rect 12173 27829 12207 27863
rect 12725 27829 12759 27863
rect 3525 27625 3559 27659
rect 4721 27625 4755 27659
rect 5273 27625 5307 27659
rect 6653 27625 6687 27659
rect 8953 27625 8987 27659
rect 10977 27625 11011 27659
rect 12541 27625 12575 27659
rect 13231 27625 13265 27659
rect 7021 27557 7055 27591
rect 10149 27557 10183 27591
rect 10701 27557 10735 27591
rect 11345 27557 11379 27591
rect 11713 27557 11747 27591
rect 12265 27557 12299 27591
rect 4169 27489 4203 27523
rect 4997 27489 5031 27523
rect 5181 27489 5215 27523
rect 5641 27489 5675 27523
rect 6009 27489 6043 27523
rect 7941 27489 7975 27523
rect 8401 27489 8435 27523
rect 13128 27489 13162 27523
rect 8493 27421 8527 27455
rect 10057 27421 10091 27455
rect 11621 27421 11655 27455
rect 4353 27353 4387 27387
rect 9505 27285 9539 27319
rect 4169 27081 4203 27115
rect 5917 27081 5951 27115
rect 6193 27081 6227 27115
rect 7021 27081 7055 27115
rect 10057 27081 10091 27115
rect 11621 27081 11655 27115
rect 12587 27081 12621 27115
rect 13093 27081 13127 27115
rect 7757 27013 7791 27047
rect 8677 26945 8711 26979
rect 10517 26945 10551 26979
rect 4997 26877 5031 26911
rect 6837 26877 6871 26911
rect 7941 26877 7975 26911
rect 8493 26877 8527 26911
rect 12173 26877 12207 26911
rect 12484 26877 12518 26911
rect 5318 26809 5352 26843
rect 6561 26809 6595 26843
rect 10609 26809 10643 26843
rect 11161 26809 11195 26843
rect 4905 26741 4939 26775
rect 7389 26741 7423 26775
rect 8953 26741 8987 26775
rect 9321 26741 9355 26775
rect 10057 26537 10091 26571
rect 10425 26537 10459 26571
rect 11529 26537 11563 26571
rect 12219 26537 12253 26571
rect 5549 26469 5583 26503
rect 10701 26469 10735 26503
rect 11253 26469 11287 26503
rect 4905 26401 4939 26435
rect 7021 26401 7055 26435
rect 8125 26401 8159 26435
rect 8585 26401 8619 26435
rect 12116 26401 12150 26435
rect 7849 26333 7883 26367
rect 8769 26333 8803 26367
rect 10609 26333 10643 26367
rect 4721 26265 4755 26299
rect 6837 26265 6871 26299
rect 5825 26197 5859 26231
rect 9413 26197 9447 26231
rect 4905 25993 4939 26027
rect 6469 25993 6503 26027
rect 10241 25993 10275 26027
rect 10885 25993 10919 26027
rect 11483 25993 11517 26027
rect 12081 25993 12115 26027
rect 5917 25857 5951 25891
rect 9321 25857 9355 25891
rect 4537 25789 4571 25823
rect 5549 25789 5583 25823
rect 7665 25789 7699 25823
rect 8033 25789 8067 25823
rect 8309 25789 8343 25823
rect 11380 25789 11414 25823
rect 5365 25721 5399 25755
rect 8493 25721 8527 25755
rect 9683 25721 9717 25755
rect 5273 25653 5307 25687
rect 8861 25653 8895 25687
rect 9229 25653 9263 25687
rect 10609 25653 10643 25687
rect 5549 25449 5583 25483
rect 6653 25449 6687 25483
rect 7021 25449 7055 25483
rect 9045 25449 9079 25483
rect 9413 25449 9447 25483
rect 10609 25449 10643 25483
rect 11437 25449 11471 25483
rect 5181 25381 5215 25415
rect 10051 25381 10085 25415
rect 10885 25381 10919 25415
rect 11897 25381 11931 25415
rect 5549 25313 5583 25347
rect 6101 25313 6135 25347
rect 7205 25313 7239 25347
rect 7297 25313 7331 25347
rect 9689 25313 9723 25347
rect 6193 25245 6227 25279
rect 4445 25177 4479 25211
rect 4813 25109 4847 25143
rect 8309 25109 8343 25143
rect 7159 24905 7193 24939
rect 8033 24905 8067 24939
rect 5457 24837 5491 24871
rect 5089 24769 5123 24803
rect 5549 24769 5583 24803
rect 6653 24769 6687 24803
rect 7389 24769 7423 24803
rect 7757 24769 7791 24803
rect 9045 24769 9079 24803
rect 10885 24769 10919 24803
rect 11253 24769 11287 24803
rect 3985 24701 4019 24735
rect 4353 24701 4387 24735
rect 5328 24701 5362 24735
rect 7251 24701 7285 24735
rect 9965 24701 9999 24735
rect 10609 24701 10643 24735
rect 3709 24633 3743 24667
rect 3801 24633 3835 24667
rect 5181 24633 5215 24667
rect 5917 24633 5951 24667
rect 6285 24633 6319 24667
rect 7021 24633 7055 24667
rect 9407 24633 9441 24667
rect 10241 24633 10275 24667
rect 10977 24633 11011 24667
rect 4721 24565 4755 24599
rect 8493 24565 8527 24599
rect 8953 24565 8987 24599
rect 3157 24361 3191 24395
rect 3525 24361 3559 24395
rect 5273 24361 5307 24395
rect 6653 24361 6687 24395
rect 7205 24361 7239 24395
rect 9781 24361 9815 24395
rect 11253 24293 11287 24327
rect 2973 24225 3007 24259
rect 4261 24225 4295 24259
rect 5733 24225 5767 24259
rect 6193 24225 6227 24259
rect 6745 24225 6779 24259
rect 7021 24225 7055 24259
rect 7849 24225 7883 24259
rect 8309 24225 8343 24259
rect 9689 24225 9723 24259
rect 10149 24225 10183 24259
rect 11345 24225 11379 24259
rect 4169 24157 4203 24191
rect 9137 24157 9171 24191
rect 5641 24089 5675 24123
rect 6837 24089 6871 24123
rect 8493 24089 8527 24123
rect 11161 24089 11195 24123
rect 5917 24021 5951 24055
rect 8769 24021 8803 24055
rect 10701 24021 10735 24055
rect 12541 24021 12575 24055
rect 2789 23817 2823 23851
rect 4353 23817 4387 23851
rect 6653 23817 6687 23851
rect 7389 23817 7423 23851
rect 8217 23817 8251 23851
rect 8953 23817 8987 23851
rect 10149 23817 10183 23851
rect 11437 23817 11471 23851
rect 12725 23817 12759 23851
rect 3341 23749 3375 23783
rect 7278 23749 7312 23783
rect 8493 23749 8527 23783
rect 8815 23749 8849 23783
rect 12614 23749 12648 23783
rect 3985 23681 4019 23715
rect 4721 23681 4755 23715
rect 5549 23681 5583 23715
rect 6285 23681 6319 23715
rect 7481 23681 7515 23715
rect 9045 23681 9079 23715
rect 10517 23681 10551 23715
rect 11897 23681 11931 23715
rect 12817 23681 12851 23715
rect 3157 23613 3191 23647
rect 3249 23613 3283 23647
rect 3525 23613 3559 23647
rect 4997 23613 5031 23647
rect 5641 23613 5675 23647
rect 7113 23613 7147 23647
rect 8677 23613 8711 23647
rect 12173 23613 12207 23647
rect 12449 23613 12483 23647
rect 9413 23545 9447 23579
rect 10609 23545 10643 23579
rect 11161 23545 11195 23579
rect 4905 23477 4939 23511
rect 7757 23477 7791 23511
rect 9689 23477 9723 23511
rect 13093 23477 13127 23511
rect 3893 23273 3927 23307
rect 5549 23273 5583 23307
rect 6837 23273 6871 23307
rect 7205 23273 7239 23307
rect 7573 23273 7607 23307
rect 9045 23273 9079 23307
rect 12725 23273 12759 23307
rect 10517 23205 10551 23239
rect 11897 23205 11931 23239
rect 2605 23137 2639 23171
rect 2789 23137 2823 23171
rect 4144 23137 4178 23171
rect 4905 23137 4939 23171
rect 5549 23137 5583 23171
rect 6101 23137 6135 23171
rect 6285 23137 6319 23171
rect 8033 23137 8067 23171
rect 8493 23137 8527 23171
rect 12081 23137 12115 23171
rect 8769 23069 8803 23103
rect 10241 23069 10275 23103
rect 10425 23069 10459 23103
rect 11069 23069 11103 23103
rect 4215 23001 4249 23035
rect 2881 22933 2915 22967
rect 3525 22933 3559 22967
rect 12173 22933 12207 22967
rect 2237 22729 2271 22763
rect 5825 22729 5859 22763
rect 6101 22729 6135 22763
rect 6469 22729 6503 22763
rect 8033 22729 8067 22763
rect 11989 22729 12023 22763
rect 12587 22729 12621 22763
rect 13599 22729 13633 22763
rect 2513 22661 2547 22695
rect 3985 22661 4019 22695
rect 8401 22661 8435 22695
rect 4905 22593 4939 22627
rect 7205 22593 7239 22627
rect 9045 22593 9079 22627
rect 10885 22593 10919 22627
rect 11161 22593 11195 22627
rect 2329 22525 2363 22559
rect 10333 22525 10367 22559
rect 12484 22525 12518 22559
rect 12909 22525 12943 22559
rect 13496 22525 13530 22559
rect 13921 22525 13955 22559
rect 2881 22457 2915 22491
rect 3433 22457 3467 22491
rect 3525 22457 3559 22491
rect 4813 22457 4847 22491
rect 5226 22457 5260 22491
rect 6929 22457 6963 22491
rect 7021 22457 7055 22491
rect 9366 22457 9400 22491
rect 10977 22457 11011 22491
rect 3249 22389 3283 22423
rect 4445 22389 4479 22423
rect 8861 22389 8895 22423
rect 9965 22389 9999 22423
rect 2697 22185 2731 22219
rect 3111 22185 3145 22219
rect 3433 22185 3467 22219
rect 4537 22185 4571 22219
rect 6653 22185 6687 22219
rect 7665 22185 7699 22219
rect 9045 22185 9079 22219
rect 10977 22185 11011 22219
rect 5318 22117 5352 22151
rect 8170 22117 8204 22151
rect 10010 22117 10044 22151
rect 11621 22117 11655 22151
rect 13185 22117 13219 22151
rect 3040 22049 3074 22083
rect 6837 22049 6871 22083
rect 8769 22049 8803 22083
rect 12449 22049 12483 22083
rect 4997 21981 5031 22015
rect 7389 21981 7423 22015
rect 7849 21981 7883 22015
rect 9689 21981 9723 22015
rect 11529 21981 11563 22015
rect 12173 21981 12207 22015
rect 13093 21981 13127 22015
rect 4905 21913 4939 21947
rect 6285 21913 6319 21947
rect 7021 21913 7055 21947
rect 11345 21913 11379 21947
rect 13645 21913 13679 21947
rect 5917 21845 5951 21879
rect 10609 21845 10643 21879
rect 4169 21641 4203 21675
rect 5641 21641 5675 21675
rect 7757 21641 7791 21675
rect 9045 21641 9079 21675
rect 9413 21641 9447 21675
rect 10517 21641 10551 21675
rect 11253 21641 11287 21675
rect 12173 21641 12207 21675
rect 13461 21641 13495 21675
rect 13829 21641 13863 21675
rect 10793 21573 10827 21607
rect 11483 21573 11517 21607
rect 3801 21505 3835 21539
rect 4721 21505 4755 21539
rect 4997 21505 5031 21539
rect 12817 21505 12851 21539
rect 6964 21437 6998 21471
rect 7389 21437 7423 21471
rect 7941 21437 7975 21471
rect 8401 21437 8435 21471
rect 9597 21437 9631 21471
rect 11391 21437 11425 21471
rect 11805 21437 11839 21471
rect 4537 21369 4571 21403
rect 4813 21369 4847 21403
rect 8677 21369 8711 21403
rect 9918 21369 9952 21403
rect 12541 21369 12575 21403
rect 12633 21369 12667 21403
rect 3065 21301 3099 21335
rect 6561 21301 6595 21335
rect 7067 21301 7101 21335
rect 7849 21097 7883 21131
rect 8125 21097 8159 21131
rect 9045 21097 9079 21131
rect 10609 21097 10643 21131
rect 12541 21097 12575 21131
rect 13139 21097 13173 21131
rect 7205 21029 7239 21063
rect 10010 21029 10044 21063
rect 11621 21029 11655 21063
rect 4813 20961 4847 20995
rect 6469 20961 6503 20995
rect 7021 20961 7055 20995
rect 8033 20961 8067 20995
rect 8493 20961 8527 20995
rect 13068 20961 13102 20995
rect 4445 20893 4479 20927
rect 7573 20893 7607 20927
rect 9689 20893 9723 20927
rect 11529 20893 11563 20927
rect 12173 20893 12207 20927
rect 12817 20893 12851 20927
rect 9505 20757 9539 20791
rect 10977 20757 11011 20791
rect 4261 20553 4295 20587
rect 5365 20553 5399 20587
rect 6561 20553 6595 20587
rect 7205 20553 7239 20587
rect 8401 20553 8435 20587
rect 8769 20553 8803 20587
rect 10149 20553 10183 20587
rect 11713 20553 11747 20587
rect 12587 20553 12621 20587
rect 13277 20553 13311 20587
rect 4997 20485 5031 20519
rect 13599 20485 13633 20519
rect 8953 20417 8987 20451
rect 10793 20417 10827 20451
rect 11161 20417 11195 20451
rect 12081 20417 12115 20451
rect 5825 20349 5859 20383
rect 7665 20349 7699 20383
rect 7849 20349 7883 20383
rect 8125 20349 8159 20383
rect 12500 20349 12534 20383
rect 12909 20349 12943 20383
rect 13496 20349 13530 20383
rect 13921 20349 13955 20383
rect 3341 20281 3375 20315
rect 3893 20281 3927 20315
rect 4445 20281 4479 20315
rect 4537 20281 4571 20315
rect 6101 20281 6135 20315
rect 9315 20281 9349 20315
rect 10609 20281 10643 20315
rect 10885 20281 10919 20315
rect 9873 20213 9907 20247
rect 3111 20009 3145 20043
rect 6929 20009 6963 20043
rect 7205 20009 7239 20043
rect 9505 20009 9539 20043
rect 11897 20009 11931 20043
rect 10425 19941 10459 19975
rect 10517 19941 10551 19975
rect 3040 19873 3074 19907
rect 4905 19873 4939 19907
rect 6469 19873 6503 19907
rect 7389 19873 7423 19907
rect 7665 19873 7699 19907
rect 9965 19873 9999 19907
rect 4997 19805 5031 19839
rect 7481 19805 7515 19839
rect 7849 19805 7883 19839
rect 10885 19805 10919 19839
rect 8401 19737 8435 19771
rect 5273 19669 5307 19703
rect 6101 19669 6135 19703
rect 8769 19669 8803 19703
rect 3065 19465 3099 19499
rect 6285 19465 6319 19499
rect 10977 19465 11011 19499
rect 5273 19397 5307 19431
rect 8493 19397 8527 19431
rect 4077 19329 4111 19363
rect 4721 19329 4755 19363
rect 6929 19329 6963 19363
rect 3709 19261 3743 19295
rect 4169 19261 4203 19295
rect 5089 19261 5123 19295
rect 5181 19261 5215 19295
rect 5457 19261 5491 19295
rect 6837 19261 6871 19295
rect 7113 19261 7147 19295
rect 7849 19261 7883 19295
rect 8309 19261 8343 19295
rect 8401 19261 8435 19295
rect 8677 19261 8711 19295
rect 9965 19261 9999 19295
rect 10425 19261 10459 19295
rect 7573 19193 7607 19227
rect 4353 19125 4387 19159
rect 5641 19125 5675 19159
rect 6561 19125 6595 19159
rect 8861 19125 8895 19159
rect 9781 19125 9815 19159
rect 10057 19125 10091 19159
rect 5181 18921 5215 18955
rect 6101 18921 6135 18955
rect 7389 18921 7423 18955
rect 10333 18921 10367 18955
rect 4629 18853 4663 18887
rect 4721 18785 4755 18819
rect 4997 18785 5031 18819
rect 6285 18785 6319 18819
rect 6561 18785 6595 18819
rect 8217 18785 8251 18819
rect 8585 18785 8619 18819
rect 9689 18785 9723 18819
rect 10701 18785 10735 18819
rect 6745 18717 6779 18751
rect 8769 18717 8803 18751
rect 11713 18717 11747 18751
rect 4813 18649 4847 18683
rect 6377 18649 6411 18683
rect 7941 18649 7975 18683
rect 9873 18649 9907 18683
rect 5825 18581 5859 18615
rect 10885 18581 10919 18615
rect 2881 18377 2915 18411
rect 3893 18377 3927 18411
rect 6377 18377 6411 18411
rect 8861 18377 8895 18411
rect 9321 18377 9355 18411
rect 10701 18377 10735 18411
rect 3157 18309 3191 18343
rect 4813 18309 4847 18343
rect 7021 18309 7055 18343
rect 2973 18173 3007 18207
rect 3525 18173 3559 18207
rect 3985 18173 4019 18207
rect 5273 18173 5307 18207
rect 5457 18173 5491 18207
rect 6837 18173 6871 18207
rect 7757 18173 7791 18207
rect 8033 18173 8067 18207
rect 8401 18173 8435 18207
rect 8585 18173 8619 18207
rect 9413 18173 9447 18207
rect 10333 18173 10367 18207
rect 11161 18173 11195 18207
rect 11621 18173 11655 18207
rect 7389 18105 7423 18139
rect 9775 18105 9809 18139
rect 4169 18037 4203 18071
rect 5089 18037 5123 18071
rect 11345 18037 11379 18071
rect 6285 17833 6319 17867
rect 6745 17833 6779 17867
rect 8585 17833 8619 17867
rect 9413 17833 9447 17867
rect 5267 17765 5301 17799
rect 10051 17765 10085 17799
rect 11529 17765 11563 17799
rect 11621 17765 11655 17799
rect 2973 17697 3007 17731
rect 4905 17697 4939 17731
rect 7481 17697 7515 17731
rect 7941 17697 7975 17731
rect 9689 17697 9723 17731
rect 8033 17629 8067 17663
rect 12173 17629 12207 17663
rect 3157 17493 3191 17527
rect 4813 17493 4847 17527
rect 5825 17493 5859 17527
rect 7113 17493 7147 17527
rect 10609 17493 10643 17527
rect 12541 17493 12575 17527
rect 3065 17289 3099 17323
rect 4261 17289 4295 17323
rect 4629 17289 4663 17323
rect 6561 17289 6595 17323
rect 7389 17289 7423 17323
rect 8953 17289 8987 17323
rect 10333 17289 10367 17323
rect 11345 17289 11379 17323
rect 11713 17289 11747 17323
rect 12173 17289 12207 17323
rect 4905 17221 4939 17255
rect 7113 17221 7147 17255
rect 5273 17153 5307 17187
rect 12541 17153 12575 17187
rect 12817 17153 12851 17187
rect 3709 17085 3743 17119
rect 4721 17085 4755 17119
rect 5733 17085 5767 17119
rect 6193 17085 6227 17119
rect 7573 17085 7607 17119
rect 8033 17085 8067 17119
rect 8309 17085 8343 17119
rect 9137 17085 9171 17119
rect 10952 17085 10986 17119
rect 5549 17017 5583 17051
rect 9499 17017 9533 17051
rect 12633 17017 12667 17051
rect 3893 16949 3927 16983
rect 5917 16949 5951 16983
rect 10057 16949 10091 16983
rect 11023 16949 11057 16983
rect 3157 16745 3191 16779
rect 5825 16745 5859 16779
rect 6561 16745 6595 16779
rect 9137 16745 9171 16779
rect 9873 16745 9907 16779
rect 11529 16745 11563 16779
rect 7573 16677 7607 16711
rect 8211 16677 8245 16711
rect 10701 16677 10735 16711
rect 12265 16677 12299 16711
rect 12817 16677 12851 16711
rect 2973 16609 3007 16643
rect 4997 16609 5031 16643
rect 5273 16609 5307 16643
rect 5457 16609 5491 16643
rect 6561 16609 6595 16643
rect 6837 16609 6871 16643
rect 7849 16609 7883 16643
rect 8769 16609 8803 16643
rect 10609 16541 10643 16575
rect 12173 16541 12207 16575
rect 11161 16473 11195 16507
rect 4629 16405 4663 16439
rect 2973 16201 3007 16235
rect 3985 16201 4019 16235
rect 4813 16201 4847 16235
rect 6377 16201 6411 16235
rect 7389 16201 7423 16235
rect 8585 16201 8619 16235
rect 8953 16201 8987 16235
rect 11023 16201 11057 16235
rect 11713 16201 11747 16235
rect 12173 16201 12207 16235
rect 12909 16201 12943 16235
rect 9137 16065 9171 16099
rect 12587 16065 12621 16099
rect 4077 15997 4111 16031
rect 5365 15997 5399 16031
rect 5641 15997 5675 16031
rect 7849 15997 7883 16031
rect 8033 15997 8067 16031
rect 10952 15997 10986 16031
rect 12500 15997 12534 16031
rect 13277 15997 13311 16031
rect 5825 15929 5859 15963
rect 7113 15929 7147 15963
rect 8309 15929 8343 15963
rect 9458 15929 9492 15963
rect 4261 15861 4295 15895
rect 10057 15861 10091 15895
rect 10609 15861 10643 15895
rect 11345 15861 11379 15895
rect 4813 15657 4847 15691
rect 6837 15657 6871 15691
rect 7021 15657 7055 15691
rect 7941 15657 7975 15691
rect 8309 15657 8343 15691
rect 8677 15657 8711 15691
rect 9137 15657 9171 15691
rect 5503 15589 5537 15623
rect 10010 15589 10044 15623
rect 11529 15589 11563 15623
rect 11621 15589 11655 15623
rect 7113 15521 7147 15555
rect 7389 15521 7423 15555
rect 8493 15521 8527 15555
rect 9689 15521 9723 15555
rect 13036 15521 13070 15555
rect 5181 15453 5215 15487
rect 12173 15453 12207 15487
rect 6101 15317 6135 15351
rect 10609 15317 10643 15351
rect 10977 15317 11011 15351
rect 13139 15317 13173 15351
rect 6009 15113 6043 15147
rect 6561 15113 6595 15147
rect 8033 15113 8067 15147
rect 8493 15113 8527 15147
rect 8769 15113 8803 15147
rect 10149 15113 10183 15147
rect 10609 15113 10643 15147
rect 11713 15113 11747 15147
rect 13921 15113 13955 15147
rect 6837 14977 6871 15011
rect 8953 14977 8987 15011
rect 10793 14977 10827 15011
rect 13599 14977 13633 15011
rect 4905 14909 4939 14943
rect 5273 14909 5307 14943
rect 5457 14909 5491 14943
rect 12265 14909 12299 14943
rect 12500 14909 12534 14943
rect 13512 14909 13546 14943
rect 7158 14841 7192 14875
rect 9274 14841 9308 14875
rect 10885 14841 10919 14875
rect 11437 14841 11471 14875
rect 4537 14773 4571 14807
rect 5273 14773 5307 14807
rect 7757 14773 7791 14807
rect 9873 14773 9907 14807
rect 12587 14773 12621 14807
rect 13001 14773 13035 14807
rect 5457 14569 5491 14603
rect 5825 14569 5859 14603
rect 7389 14569 7423 14603
rect 7849 14569 7883 14603
rect 8953 14569 8987 14603
rect 9965 14569 9999 14603
rect 11529 14569 11563 14603
rect 6561 14501 6595 14535
rect 10517 14501 10551 14535
rect 12081 14501 12115 14535
rect 12633 14501 12667 14535
rect 5064 14433 5098 14467
rect 8125 14433 8159 14467
rect 8401 14433 8435 14467
rect 11069 14433 11103 14467
rect 6469 14365 6503 14399
rect 7113 14365 7147 14399
rect 8493 14365 8527 14399
rect 10425 14365 10459 14399
rect 11989 14365 12023 14399
rect 5135 14229 5169 14263
rect 3019 14025 3053 14059
rect 4445 14025 4479 14059
rect 4813 14025 4847 14059
rect 6285 14025 6319 14059
rect 6653 14025 6687 14059
rect 8033 14025 8067 14059
rect 10057 14025 10091 14059
rect 11161 14025 11195 14059
rect 11621 14025 11655 14059
rect 12725 14025 12759 14059
rect 3433 13957 3467 13991
rect 11897 13957 11931 13991
rect 4905 13889 4939 13923
rect 9413 13889 9447 13923
rect 10885 13889 10919 13923
rect 2948 13821 2982 13855
rect 3928 13821 3962 13855
rect 4031 13821 4065 13855
rect 5825 13821 5859 13855
rect 7573 13821 7607 13855
rect 8401 13821 8435 13855
rect 8861 13821 8895 13855
rect 5267 13753 5301 13787
rect 6929 13753 6963 13787
rect 7021 13753 7055 13787
rect 10241 13753 10275 13787
rect 10333 13753 10367 13787
rect 8677 13685 8711 13719
rect 5273 13481 5307 13515
rect 6745 13481 6779 13515
rect 7113 13481 7147 13515
rect 8861 13481 8895 13515
rect 10701 13481 10735 13515
rect 11391 13481 11425 13515
rect 4261 13413 4295 13447
rect 4353 13413 4387 13447
rect 5825 13413 5859 13447
rect 5917 13413 5951 13447
rect 7986 13413 8020 13447
rect 9873 13413 9907 13447
rect 11288 13345 11322 13379
rect 4905 13277 4939 13311
rect 6469 13277 6503 13311
rect 7665 13277 7699 13311
rect 9781 13277 9815 13311
rect 10425 13277 10459 13311
rect 8585 13141 8619 13175
rect 3709 12937 3743 12971
rect 6193 12937 6227 12971
rect 7665 12937 7699 12971
rect 8953 12937 8987 12971
rect 10885 12937 10919 12971
rect 11897 12937 11931 12971
rect 4077 12869 4111 12903
rect 5825 12869 5859 12903
rect 6561 12801 6595 12835
rect 7297 12801 7331 12835
rect 7757 12801 7791 12835
rect 10517 12801 10551 12835
rect 4220 12733 4254 12767
rect 4629 12733 4663 12767
rect 11136 12733 11170 12767
rect 11529 12733 11563 12767
rect 4307 12665 4341 12699
rect 5273 12665 5307 12699
rect 5365 12665 5399 12699
rect 8078 12665 8112 12699
rect 9321 12665 9355 12699
rect 9597 12665 9631 12699
rect 9689 12665 9723 12699
rect 10241 12665 10275 12699
rect 5089 12597 5123 12631
rect 8677 12597 8711 12631
rect 11207 12597 11241 12631
rect 5043 12393 5077 12427
rect 5365 12393 5399 12427
rect 7849 12393 7883 12427
rect 6101 12325 6135 12359
rect 6653 12325 6687 12359
rect 8217 12325 8251 12359
rect 9873 12325 9907 12359
rect 11437 12325 11471 12359
rect 11989 12325 12023 12359
rect 4940 12257 4974 12291
rect 12852 12257 12886 12291
rect 6009 12189 6043 12223
rect 8125 12189 8159 12223
rect 9781 12189 9815 12223
rect 11345 12189 11379 12223
rect 12955 12189 12989 12223
rect 8677 12121 8711 12155
rect 10333 12121 10367 12155
rect 9505 12053 9539 12087
rect 4905 11849 4939 11883
rect 5641 11849 5675 11883
rect 6561 11849 6595 11883
rect 7297 11849 7331 11883
rect 8677 11849 8711 11883
rect 9505 11849 9539 11883
rect 11161 11849 11195 11883
rect 12081 11849 12115 11883
rect 13277 11849 13311 11883
rect 5181 11781 5215 11815
rect 7665 11781 7699 11815
rect 9781 11713 9815 11747
rect 11391 11713 11425 11747
rect 4721 11645 4755 11679
rect 5800 11645 5834 11679
rect 6193 11645 6227 11679
rect 7757 11645 7791 11679
rect 8953 11645 8987 11679
rect 11288 11645 11322 11679
rect 11713 11645 11747 11679
rect 12516 11645 12550 11679
rect 12909 11645 12943 11679
rect 8078 11577 8112 11611
rect 9873 11577 9907 11611
rect 10425 11577 10459 11611
rect 5871 11509 5905 11543
rect 10701 11509 10735 11543
rect 12587 11509 12621 11543
rect 5733 11305 5767 11339
rect 7297 11305 7331 11339
rect 9137 11305 9171 11339
rect 9413 11305 9447 11339
rect 11391 11305 11425 11339
rect 7021 11237 7055 11271
rect 8170 11237 8204 11271
rect 9873 11237 9907 11271
rect 10425 11237 10459 11271
rect 4721 11169 4755 11203
rect 5273 11169 5307 11203
rect 6561 11169 6595 11203
rect 6745 11169 6779 11203
rect 11288 11169 11322 11203
rect 12332 11169 12366 11203
rect 5457 11101 5491 11135
rect 7849 11101 7883 11135
rect 9781 11101 9815 11135
rect 7757 11033 7791 11067
rect 6101 10965 6135 10999
rect 8769 10965 8803 10999
rect 12403 10965 12437 10999
rect 4077 10761 4111 10795
rect 4813 10761 4847 10795
rect 6377 10761 6411 10795
rect 7941 10761 7975 10795
rect 9505 10761 9539 10795
rect 11437 10761 11471 10795
rect 12633 10761 12667 10795
rect 9137 10693 9171 10727
rect 5549 10625 5583 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 8585 10625 8619 10659
rect 10425 10625 10459 10659
rect 11805 10625 11839 10659
rect 4169 10489 4203 10523
rect 5273 10489 5307 10523
rect 5365 10489 5399 10523
rect 7021 10489 7055 10523
rect 8677 10489 8711 10523
rect 9965 10489 9999 10523
rect 10149 10489 10183 10523
rect 10241 10489 10275 10523
rect 8401 10421 8435 10455
rect 11069 10421 11103 10455
rect 5273 10217 5307 10251
rect 6745 10217 6779 10251
rect 8309 10217 8343 10251
rect 8769 10217 8803 10251
rect 10609 10217 10643 10251
rect 5911 10149 5945 10183
rect 7481 10149 7515 10183
rect 8033 10149 8067 10183
rect 10051 10149 10085 10183
rect 11437 10149 11471 10183
rect 4537 10081 4571 10115
rect 6469 10081 6503 10115
rect 7113 10081 7147 10115
rect 5549 10013 5583 10047
rect 7389 10013 7423 10047
rect 9045 10013 9079 10047
rect 9689 10013 9723 10047
rect 4721 9877 4755 9911
rect 4537 9673 4571 9707
rect 6285 9673 6319 9707
rect 9781 9673 9815 9707
rect 5917 9605 5951 9639
rect 7849 9605 7883 9639
rect 10701 9537 10735 9571
rect 11345 9537 11379 9571
rect 4169 9469 4203 9503
rect 4997 9469 5031 9503
rect 7113 9469 7147 9503
rect 7297 9469 7331 9503
rect 8585 9469 8619 9503
rect 8861 9469 8895 9503
rect 10241 9469 10275 9503
rect 10425 9469 10459 9503
rect 4905 9401 4939 9435
rect 5359 9401 5393 9435
rect 8309 9401 8343 9435
rect 9137 9401 9171 9435
rect 10977 9401 11011 9435
rect 6561 9333 6595 9367
rect 6929 9333 6963 9367
rect 5181 9129 5215 9163
rect 5457 9129 5491 9163
rect 6469 9129 6503 9163
rect 8493 9129 8527 9163
rect 8769 9129 8803 9163
rect 9827 9129 9861 9163
rect 7475 9061 7509 9095
rect 10517 9061 10551 9095
rect 4388 8993 4422 9027
rect 5549 8993 5583 9027
rect 5825 8993 5859 9027
rect 6929 8993 6963 9027
rect 9756 8993 9790 9027
rect 10701 8993 10735 9027
rect 7113 8925 7147 8959
rect 10241 8857 10275 8891
rect 10885 8857 10919 8891
rect 4491 8789 4525 8823
rect 8033 8789 8067 8823
rect 4353 8585 4387 8619
rect 4629 8585 4663 8619
rect 4997 8585 5031 8619
rect 6193 8585 6227 8619
rect 9229 8585 9263 8619
rect 9505 8585 9539 8619
rect 10793 8585 10827 8619
rect 7757 8517 7791 8551
rect 5917 8449 5951 8483
rect 7021 8449 7055 8483
rect 8125 8449 8159 8483
rect 5181 8381 5215 8415
rect 5641 8381 5675 8415
rect 8493 8381 8527 8415
rect 8769 8381 8803 8415
rect 9505 8381 9539 8415
rect 9781 8381 9815 8415
rect 10241 8381 10275 8415
rect 7205 8313 7239 8347
rect 8953 8313 8987 8347
rect 9689 8313 9723 8347
rect 9873 8245 9907 8279
rect 6561 7973 6595 8007
rect 8125 7973 8159 8007
rect 10051 7973 10085 8007
rect 5089 7905 5123 7939
rect 5365 7905 5399 7939
rect 9689 7905 9723 7939
rect 5549 7837 5583 7871
rect 6469 7837 6503 7871
rect 7113 7837 7147 7871
rect 8033 7837 8067 7871
rect 8677 7837 8711 7871
rect 11437 7837 11471 7871
rect 6193 7701 6227 7735
rect 10609 7701 10643 7735
rect 4905 7497 4939 7531
rect 7757 7497 7791 7531
rect 8125 7497 8159 7531
rect 10793 7497 10827 7531
rect 4537 7429 4571 7463
rect 9137 7429 9171 7463
rect 10425 7429 10459 7463
rect 11115 7429 11149 7463
rect 6837 7361 6871 7395
rect 9229 7361 9263 7395
rect 5457 7293 5491 7327
rect 5641 7293 5675 7327
rect 11044 7293 11078 7327
rect 11437 7293 11471 7327
rect 5917 7225 5951 7259
rect 7199 7225 7233 7259
rect 9591 7225 9625 7259
rect 6193 7157 6227 7191
rect 6653 7157 6687 7191
rect 8401 7157 8435 7191
rect 10149 7157 10183 7191
rect 5365 6953 5399 6987
rect 9229 6953 9263 6987
rect 10885 6953 10919 6987
rect 6187 6885 6221 6919
rect 8078 6885 8112 6919
rect 10051 6885 10085 6919
rect 11621 6885 11655 6919
rect 4848 6817 4882 6851
rect 4951 6817 4985 6851
rect 5733 6817 5767 6851
rect 7573 6817 7607 6851
rect 7757 6817 7791 6851
rect 9689 6817 9723 6851
rect 10609 6817 10643 6851
rect 5825 6749 5859 6783
rect 7021 6749 7055 6783
rect 11529 6749 11563 6783
rect 11989 6749 12023 6783
rect 6745 6613 6779 6647
rect 8677 6613 8711 6647
rect 4813 6409 4847 6443
rect 6561 6409 6595 6443
rect 7849 6409 7883 6443
rect 8401 6409 8435 6443
rect 9781 6409 9815 6443
rect 11437 6409 11471 6443
rect 11805 6409 11839 6443
rect 7205 6273 7239 6307
rect 8677 6273 8711 6307
rect 8953 6273 8987 6307
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 5768 6205 5802 6239
rect 6193 6205 6227 6239
rect 5871 6137 5905 6171
rect 6929 6137 6963 6171
rect 7021 6137 7055 6171
rect 8769 6137 8803 6171
rect 10425 6137 10459 6171
rect 10977 6137 11011 6171
rect 5641 6069 5675 6103
rect 6101 5865 6135 5899
rect 7389 5865 7423 5899
rect 8769 5865 8803 5899
rect 9873 5865 9907 5899
rect 7021 5797 7055 5831
rect 7757 5797 7791 5831
rect 7849 5797 7883 5831
rect 8401 5797 8435 5831
rect 10241 5797 10275 5831
rect 6285 5729 6319 5763
rect 6469 5729 6503 5763
rect 10793 5729 10827 5763
rect 11688 5729 11722 5763
rect 10149 5661 10183 5695
rect 11759 5525 11793 5559
rect 5641 5321 5675 5355
rect 6285 5321 6319 5355
rect 6561 5321 6595 5355
rect 7205 5321 7239 5355
rect 10333 5321 10367 5355
rect 11713 5321 11747 5355
rect 12909 5321 12943 5355
rect 7573 5253 7607 5287
rect 9045 5253 9079 5287
rect 11253 5253 11287 5287
rect 8677 5185 8711 5219
rect 9781 5185 9815 5219
rect 10609 5185 10643 5219
rect 5800 5117 5834 5151
rect 7665 5117 7699 5151
rect 8125 5117 8159 5151
rect 9229 5117 9263 5151
rect 9689 5117 9723 5151
rect 10839 5117 10873 5151
rect 12516 5117 12550 5151
rect 8401 5049 8435 5083
rect 5871 4981 5905 5015
rect 10931 4981 10965 5015
rect 12587 4981 12621 5015
rect 5273 4777 5307 4811
rect 7665 4777 7699 4811
rect 9229 4777 9263 4811
rect 6653 4709 6687 4743
rect 9873 4709 9907 4743
rect 5508 4641 5542 4675
rect 8033 4641 8067 4675
rect 8585 4641 8619 4675
rect 11253 4641 11287 4675
rect 12357 4641 12391 4675
rect 13461 4641 13495 4675
rect 5595 4573 5629 4607
rect 6009 4573 6043 4607
rect 6561 4573 6595 4607
rect 8769 4573 8803 4607
rect 9781 4573 9815 4607
rect 10149 4573 10183 4607
rect 7113 4505 7147 4539
rect 12541 4505 12575 4539
rect 6285 4437 6319 4471
rect 10793 4437 10827 4471
rect 11437 4437 11471 4471
rect 13645 4437 13679 4471
rect 7941 4233 7975 4267
rect 11253 4233 11287 4267
rect 12265 4233 12299 4267
rect 13369 4233 13403 4267
rect 5089 4097 5123 4131
rect 7205 4097 7239 4131
rect 8217 4097 8251 4131
rect 9689 4097 9723 4131
rect 10241 4097 10275 4131
rect 10885 4097 10919 4131
rect 11621 4097 11655 4131
rect 4220 4029 4254 4063
rect 5273 4029 5307 4063
rect 5641 4029 5675 4063
rect 8401 4029 8435 4063
rect 12449 4029 12483 4063
rect 13001 4029 13035 4063
rect 13588 4029 13622 4063
rect 14013 4029 14047 4063
rect 4307 3961 4341 3995
rect 5917 3961 5951 3995
rect 6929 3961 6963 3995
rect 7021 3961 7055 3995
rect 8722 3961 8756 3995
rect 10333 3961 10367 3995
rect 4721 3893 4755 3927
rect 6193 3893 6227 3927
rect 6653 3893 6687 3927
rect 9321 3893 9355 3927
rect 10057 3893 10091 3927
rect 12633 3893 12667 3927
rect 13691 3893 13725 3927
rect 9413 3689 9447 3723
rect 11161 3689 11195 3723
rect 6279 3621 6313 3655
rect 8170 3621 8204 3655
rect 9045 3621 9079 3655
rect 9873 3621 9907 3655
rect 11437 3621 11471 3655
rect 4629 3553 4663 3587
rect 4905 3553 4939 3587
rect 5089 3553 5123 3587
rect 7113 3553 7147 3587
rect 7849 3553 7883 3587
rect 10701 3553 10735 3587
rect 13461 3553 13495 3587
rect 5917 3485 5951 3519
rect 9781 3485 9815 3519
rect 11345 3485 11379 3519
rect 6837 3417 6871 3451
rect 8769 3417 8803 3451
rect 10333 3417 10367 3451
rect 11897 3417 11931 3451
rect 5365 3349 5399 3383
rect 5733 3349 5767 3383
rect 7481 3349 7515 3383
rect 13645 3349 13679 3383
rect 4307 3145 4341 3179
rect 6285 3145 6319 3179
rect 6561 3145 6595 3179
rect 7757 3145 7791 3179
rect 8033 3145 8067 3179
rect 8401 3145 8435 3179
rect 9505 3145 9539 3179
rect 9873 3145 9907 3179
rect 11437 3145 11471 3179
rect 11805 3145 11839 3179
rect 13001 3145 13035 3179
rect 13691 3145 13725 3179
rect 4077 3077 4111 3111
rect 4997 3077 5031 3111
rect 10977 3077 11011 3111
rect 12633 3077 12667 3111
rect 13461 3077 13495 3111
rect 5273 3009 5307 3043
rect 5917 3009 5951 3043
rect 6837 3009 6871 3043
rect 8585 3009 8619 3043
rect 10425 3009 10459 3043
rect 3224 2941 3258 2975
rect 3709 2941 3743 2975
rect 4220 2941 4254 2975
rect 12449 2941 12483 2975
rect 13588 2941 13622 2975
rect 14013 2941 14047 2975
rect 4629 2873 4663 2907
rect 5365 2873 5399 2907
rect 7199 2873 7233 2907
rect 8906 2873 8940 2907
rect 10241 2873 10275 2907
rect 10517 2873 10551 2907
rect 3295 2805 3329 2839
rect 4399 2601 4433 2635
rect 6285 2601 6319 2635
rect 6745 2601 6779 2635
rect 8033 2601 8067 2635
rect 9505 2601 9539 2635
rect 11161 2601 11195 2635
rect 13185 2601 13219 2635
rect 6009 2533 6043 2567
rect 7205 2533 7239 2567
rect 7757 2533 7791 2567
rect 9965 2533 9999 2567
rect 10517 2533 10551 2567
rect 4296 2465 4330 2499
rect 4721 2465 4755 2499
rect 5181 2465 5215 2499
rect 5917 2465 5951 2499
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 11345 2465 11379 2499
rect 11897 2465 11931 2499
rect 12633 2465 12667 2499
rect 7113 2397 7147 2431
rect 8401 2397 8435 2431
rect 9873 2397 9907 2431
rect 10793 2397 10827 2431
rect 8769 2261 8803 2295
rect 11529 2261 11563 2295
rect 12817 2261 12851 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 8113 37315 8171 37321
rect 8113 37281 8125 37315
rect 8159 37312 8171 37315
rect 8570 37312 8576 37324
rect 8159 37284 8576 37312
rect 8159 37281 8171 37284
rect 8113 37275 8171 37281
rect 8570 37272 8576 37284
rect 8628 37272 8634 37324
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 10962 36904 10968 36916
rect 10923 36876 10968 36904
rect 10962 36864 10968 36876
rect 11020 36864 11026 36916
rect 6984 36703 7042 36709
rect 6984 36669 6996 36703
rect 7030 36700 7042 36703
rect 8021 36703 8079 36709
rect 8021 36700 8033 36703
rect 7030 36672 7328 36700
rect 7030 36669 7042 36672
rect 6984 36663 7042 36669
rect 7300 36576 7328 36672
rect 7852 36672 8033 36700
rect 7055 36567 7113 36573
rect 7055 36533 7067 36567
rect 7101 36564 7113 36567
rect 7190 36564 7196 36576
rect 7101 36536 7196 36564
rect 7101 36533 7113 36536
rect 7055 36527 7113 36533
rect 7190 36524 7196 36536
rect 7248 36524 7254 36576
rect 7282 36524 7288 36576
rect 7340 36564 7346 36576
rect 7377 36567 7435 36573
rect 7377 36564 7389 36567
rect 7340 36536 7389 36564
rect 7340 36524 7346 36536
rect 7377 36533 7389 36536
rect 7423 36533 7435 36567
rect 7377 36527 7435 36533
rect 7558 36524 7564 36576
rect 7616 36564 7622 36576
rect 7852 36573 7880 36672
rect 8021 36669 8033 36672
rect 8067 36669 8079 36703
rect 8570 36700 8576 36712
rect 8531 36672 8576 36700
rect 8021 36663 8079 36669
rect 8570 36660 8576 36672
rect 8628 36660 8634 36712
rect 10781 36703 10839 36709
rect 10781 36669 10793 36703
rect 10827 36700 10839 36703
rect 10827 36672 11192 36700
rect 10827 36669 10839 36672
rect 10781 36663 10839 36669
rect 11164 36576 11192 36672
rect 7837 36567 7895 36573
rect 7837 36564 7849 36567
rect 7616 36536 7849 36564
rect 7616 36524 7622 36536
rect 7837 36533 7849 36536
rect 7883 36533 7895 36567
rect 7837 36527 7895 36533
rect 8297 36567 8355 36573
rect 8297 36533 8309 36567
rect 8343 36564 8355 36567
rect 8386 36564 8392 36576
rect 8343 36536 8392 36564
rect 8343 36533 8355 36536
rect 8297 36527 8355 36533
rect 8386 36524 8392 36536
rect 8444 36524 8450 36576
rect 11146 36524 11152 36576
rect 11204 36564 11210 36576
rect 11333 36567 11391 36573
rect 11333 36564 11345 36567
rect 11204 36536 11345 36564
rect 11204 36524 11210 36536
rect 11333 36533 11345 36536
rect 11379 36533 11391 36567
rect 11333 36527 11391 36533
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 9861 36363 9919 36369
rect 9861 36329 9873 36363
rect 9907 36360 9919 36363
rect 10686 36360 10692 36372
rect 9907 36332 10692 36360
rect 9907 36329 9919 36332
rect 9861 36323 9919 36329
rect 10686 36320 10692 36332
rect 10744 36320 10750 36372
rect 11425 36363 11483 36369
rect 11425 36329 11437 36363
rect 11471 36360 11483 36363
rect 12342 36360 12348 36372
rect 11471 36332 12348 36360
rect 11471 36329 11483 36332
rect 11425 36323 11483 36329
rect 12342 36320 12348 36332
rect 12400 36320 12406 36372
rect 6914 36252 6920 36304
rect 6972 36292 6978 36304
rect 7285 36295 7343 36301
rect 7285 36292 7297 36295
rect 6972 36264 7297 36292
rect 6972 36252 6978 36264
rect 7285 36261 7297 36264
rect 7331 36261 7343 36295
rect 7285 36255 7343 36261
rect 9677 36227 9735 36233
rect 9677 36193 9689 36227
rect 9723 36224 9735 36227
rect 9766 36224 9772 36236
rect 9723 36196 9772 36224
rect 9723 36193 9735 36196
rect 9677 36187 9735 36193
rect 9766 36184 9772 36196
rect 9824 36184 9830 36236
rect 11238 36224 11244 36236
rect 11199 36196 11244 36224
rect 11238 36184 11244 36196
rect 11296 36184 11302 36236
rect 7190 36156 7196 36168
rect 7151 36128 7196 36156
rect 7190 36116 7196 36128
rect 7248 36116 7254 36168
rect 7742 36088 7748 36100
rect 7703 36060 7748 36088
rect 7742 36048 7748 36060
rect 7800 36048 7806 36100
rect 8570 35980 8576 36032
rect 8628 36020 8634 36032
rect 8757 36023 8815 36029
rect 8757 36020 8769 36023
rect 8628 35992 8769 36020
rect 8628 35980 8634 35992
rect 8757 35989 8769 35992
rect 8803 36020 8815 36023
rect 9582 36020 9588 36032
rect 8803 35992 9588 36020
rect 8803 35989 8815 35992
rect 8757 35983 8815 35989
rect 9582 35980 9588 35992
rect 9640 35980 9646 36032
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 7190 35776 7196 35828
rect 7248 35816 7254 35828
rect 8113 35819 8171 35825
rect 8113 35816 8125 35819
rect 7248 35788 8125 35816
rect 7248 35776 7254 35788
rect 8113 35785 8125 35788
rect 8159 35785 8171 35819
rect 8113 35779 8171 35785
rect 10413 35819 10471 35825
rect 10413 35785 10425 35819
rect 10459 35816 10471 35819
rect 11330 35816 11336 35828
rect 10459 35788 11336 35816
rect 10459 35785 10471 35788
rect 10413 35779 10471 35785
rect 11330 35776 11336 35788
rect 11388 35776 11394 35828
rect 11471 35819 11529 35825
rect 11471 35785 11483 35819
rect 11517 35816 11529 35819
rect 12066 35816 12072 35828
rect 11517 35788 12072 35816
rect 11517 35785 11529 35788
rect 11471 35779 11529 35785
rect 12066 35776 12072 35788
rect 12124 35776 12130 35828
rect 12621 35819 12679 35825
rect 12621 35785 12633 35819
rect 12667 35816 12679 35819
rect 13722 35816 13728 35828
rect 12667 35788 13728 35816
rect 12667 35785 12679 35788
rect 12621 35779 12679 35785
rect 13722 35776 13728 35788
rect 13780 35776 13786 35828
rect 7742 35748 7748 35760
rect 7703 35720 7748 35748
rect 7742 35708 7748 35720
rect 7800 35708 7806 35760
rect 6914 35640 6920 35692
rect 6972 35680 6978 35692
rect 7193 35683 7251 35689
rect 7193 35680 7205 35683
rect 6972 35652 7205 35680
rect 6972 35640 6978 35652
rect 7193 35649 7205 35652
rect 7239 35649 7251 35683
rect 7193 35643 7251 35649
rect 8665 35615 8723 35621
rect 8665 35612 8677 35615
rect 8496 35584 8677 35612
rect 6273 35547 6331 35553
rect 6273 35513 6285 35547
rect 6319 35544 6331 35547
rect 7006 35544 7012 35556
rect 6319 35516 7012 35544
rect 6319 35513 6331 35516
rect 6273 35507 6331 35513
rect 7006 35504 7012 35516
rect 7064 35504 7070 35556
rect 7285 35547 7343 35553
rect 7285 35513 7297 35547
rect 7331 35513 7343 35547
rect 7285 35507 7343 35513
rect 6641 35479 6699 35485
rect 6641 35445 6653 35479
rect 6687 35476 6699 35479
rect 6730 35476 6736 35488
rect 6687 35448 6736 35476
rect 6687 35445 6699 35448
rect 6641 35439 6699 35445
rect 6730 35436 6736 35448
rect 6788 35436 6794 35488
rect 7024 35476 7052 35504
rect 7300 35476 7328 35507
rect 7024 35448 7328 35476
rect 7466 35436 7472 35488
rect 7524 35476 7530 35488
rect 8496 35485 8524 35584
rect 8665 35581 8677 35584
rect 8711 35581 8723 35615
rect 8665 35575 8723 35581
rect 9217 35615 9275 35621
rect 9217 35581 9229 35615
rect 9263 35612 9275 35615
rect 9490 35612 9496 35624
rect 9263 35584 9496 35612
rect 9263 35581 9275 35584
rect 9217 35575 9275 35581
rect 9490 35572 9496 35584
rect 9548 35572 9554 35624
rect 10226 35612 10232 35624
rect 10187 35584 10232 35612
rect 10226 35572 10232 35584
rect 10284 35612 10290 35624
rect 10781 35615 10839 35621
rect 10781 35612 10793 35615
rect 10284 35584 10793 35612
rect 10284 35572 10290 35584
rect 10781 35581 10793 35584
rect 10827 35581 10839 35615
rect 10781 35575 10839 35581
rect 11400 35615 11458 35621
rect 11400 35581 11412 35615
rect 11446 35612 11458 35615
rect 12437 35615 12495 35621
rect 11446 35584 12020 35612
rect 11446 35581 11458 35584
rect 11400 35575 11458 35581
rect 11992 35488 12020 35584
rect 12437 35581 12449 35615
rect 12483 35612 12495 35615
rect 12483 35584 13032 35612
rect 12483 35581 12495 35584
rect 12437 35575 12495 35581
rect 13004 35488 13032 35584
rect 8481 35479 8539 35485
rect 8481 35476 8493 35479
rect 7524 35448 8493 35476
rect 7524 35436 7530 35448
rect 8481 35445 8493 35448
rect 8527 35445 8539 35479
rect 8754 35476 8760 35488
rect 8715 35448 8760 35476
rect 8481 35439 8539 35445
rect 8754 35436 8760 35448
rect 8812 35436 8818 35488
rect 9766 35476 9772 35488
rect 9727 35448 9772 35476
rect 9766 35436 9772 35448
rect 9824 35436 9830 35488
rect 11330 35436 11336 35488
rect 11388 35476 11394 35488
rect 11793 35479 11851 35485
rect 11793 35476 11805 35479
rect 11388 35448 11805 35476
rect 11388 35436 11394 35448
rect 11793 35445 11805 35448
rect 11839 35445 11851 35479
rect 11793 35439 11851 35445
rect 11974 35436 11980 35488
rect 12032 35476 12038 35488
rect 12161 35479 12219 35485
rect 12161 35476 12173 35479
rect 12032 35448 12173 35476
rect 12032 35436 12038 35448
rect 12161 35445 12173 35448
rect 12207 35445 12219 35479
rect 12986 35476 12992 35488
rect 12947 35448 12992 35476
rect 12161 35439 12219 35445
rect 12986 35436 12992 35448
rect 13044 35436 13050 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 6914 35232 6920 35284
rect 6972 35272 6978 35284
rect 7837 35275 7895 35281
rect 7837 35272 7849 35275
rect 6972 35244 7849 35272
rect 6972 35232 6978 35244
rect 7837 35241 7849 35244
rect 7883 35241 7895 35275
rect 7837 35235 7895 35241
rect 11701 35275 11759 35281
rect 11701 35241 11713 35275
rect 11747 35272 11759 35275
rect 12066 35272 12072 35284
rect 11747 35244 12072 35272
rect 11747 35241 11759 35244
rect 11701 35235 11759 35241
rect 12066 35232 12072 35244
rect 12124 35232 12130 35284
rect 12897 35275 12955 35281
rect 12897 35241 12909 35275
rect 12943 35272 12955 35275
rect 14182 35272 14188 35284
rect 12943 35244 14188 35272
rect 12943 35241 12955 35244
rect 12897 35235 12955 35241
rect 14182 35232 14188 35244
rect 14240 35232 14246 35284
rect 7006 35204 7012 35216
rect 6967 35176 7012 35204
rect 7006 35164 7012 35176
rect 7064 35164 7070 35216
rect 9858 35164 9864 35216
rect 9916 35204 9922 35216
rect 9953 35207 10011 35213
rect 9953 35204 9965 35207
rect 9916 35176 9965 35204
rect 9916 35164 9922 35176
rect 9953 35173 9965 35176
rect 9999 35173 10011 35207
rect 9953 35167 10011 35173
rect 5880 35139 5938 35145
rect 5880 35105 5892 35139
rect 5926 35136 5938 35139
rect 6270 35136 6276 35148
rect 5926 35108 6276 35136
rect 5926 35105 5938 35108
rect 5880 35099 5938 35105
rect 6270 35096 6276 35108
rect 6328 35096 6334 35148
rect 8294 35096 8300 35148
rect 8352 35136 8358 35148
rect 8608 35139 8666 35145
rect 8608 35136 8620 35139
rect 8352 35108 8620 35136
rect 8352 35096 8358 35108
rect 8608 35105 8620 35108
rect 8654 35105 8666 35139
rect 8608 35099 8666 35105
rect 11238 35096 11244 35148
rect 11296 35136 11302 35148
rect 11517 35139 11575 35145
rect 11517 35136 11529 35139
rect 11296 35108 11529 35136
rect 11296 35096 11302 35108
rect 11517 35105 11529 35108
rect 11563 35105 11575 35139
rect 11517 35099 11575 35105
rect 12434 35096 12440 35148
rect 12492 35136 12498 35148
rect 12713 35139 12771 35145
rect 12713 35136 12725 35139
rect 12492 35108 12725 35136
rect 12492 35096 12498 35108
rect 12713 35105 12725 35108
rect 12759 35105 12771 35139
rect 12713 35099 12771 35105
rect 6917 35071 6975 35077
rect 6917 35037 6929 35071
rect 6963 35037 6975 35071
rect 6917 35031 6975 35037
rect 7561 35071 7619 35077
rect 7561 35037 7573 35071
rect 7607 35068 7619 35071
rect 7926 35068 7932 35080
rect 7607 35040 7932 35068
rect 7607 35037 7619 35040
rect 7561 35031 7619 35037
rect 5951 35003 6009 35009
rect 5951 34969 5963 35003
rect 5997 35000 6009 35003
rect 6641 35003 6699 35009
rect 6641 35000 6653 35003
rect 5997 34972 6653 35000
rect 5997 34969 6009 34972
rect 5951 34963 6009 34969
rect 6641 34969 6653 34972
rect 6687 35000 6699 35003
rect 6932 35000 6960 35031
rect 7926 35028 7932 35040
rect 7984 35028 7990 35080
rect 8711 35071 8769 35077
rect 8711 35037 8723 35071
rect 8757 35068 8769 35071
rect 9398 35068 9404 35080
rect 8757 35040 9404 35068
rect 8757 35037 8769 35040
rect 8711 35031 8769 35037
rect 9398 35028 9404 35040
rect 9456 35068 9462 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9456 35040 9873 35068
rect 9456 35028 9462 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 10505 35071 10563 35077
rect 10505 35037 10517 35071
rect 10551 35068 10563 35071
rect 11054 35068 11060 35080
rect 10551 35040 11060 35068
rect 10551 35037 10563 35040
rect 10505 35031 10563 35037
rect 11054 35028 11060 35040
rect 11112 35028 11118 35080
rect 6687 34972 6960 35000
rect 6687 34969 6699 34972
rect 6641 34963 6699 34969
rect 5258 34932 5264 34944
rect 5219 34904 5264 34932
rect 5258 34892 5264 34904
rect 5316 34892 5322 34944
rect 10873 34935 10931 34941
rect 10873 34901 10885 34935
rect 10919 34932 10931 34935
rect 10962 34932 10968 34944
rect 10919 34904 10968 34932
rect 10919 34901 10931 34904
rect 10873 34895 10931 34901
rect 10962 34892 10968 34904
rect 11020 34892 11026 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 4295 34731 4353 34737
rect 4295 34697 4307 34731
rect 4341 34728 4353 34731
rect 5442 34728 5448 34740
rect 4341 34700 5448 34728
rect 4341 34697 4353 34700
rect 4295 34691 4353 34697
rect 5442 34688 5448 34700
rect 5500 34688 5506 34740
rect 6270 34728 6276 34740
rect 6231 34700 6276 34728
rect 6270 34688 6276 34700
rect 6328 34688 6334 34740
rect 7006 34688 7012 34740
rect 7064 34728 7070 34740
rect 7745 34731 7803 34737
rect 7745 34728 7757 34731
rect 7064 34700 7757 34728
rect 7064 34688 7070 34700
rect 7745 34697 7757 34700
rect 7791 34697 7803 34731
rect 7745 34691 7803 34697
rect 8294 34688 8300 34740
rect 8352 34728 8358 34740
rect 8478 34728 8484 34740
rect 8352 34700 8484 34728
rect 8352 34688 8358 34700
rect 8478 34688 8484 34700
rect 8536 34688 8542 34740
rect 13630 34728 13636 34740
rect 13591 34700 13636 34728
rect 13630 34688 13636 34700
rect 13688 34688 13694 34740
rect 10962 34660 10968 34672
rect 10520 34632 10968 34660
rect 8205 34595 8263 34601
rect 8205 34561 8217 34595
rect 8251 34592 8263 34595
rect 8665 34595 8723 34601
rect 8665 34592 8677 34595
rect 8251 34564 8677 34592
rect 8251 34561 8263 34564
rect 8205 34555 8263 34561
rect 8665 34561 8677 34564
rect 8711 34592 8723 34595
rect 8754 34592 8760 34604
rect 8711 34564 8760 34592
rect 8711 34561 8723 34564
rect 8665 34555 8723 34561
rect 8754 34552 8760 34564
rect 8812 34552 8818 34604
rect 10520 34601 10548 34632
rect 10962 34620 10968 34632
rect 11020 34620 11026 34672
rect 10505 34595 10563 34601
rect 10505 34561 10517 34595
rect 10551 34561 10563 34595
rect 10870 34592 10876 34604
rect 10831 34564 10876 34592
rect 10505 34555 10563 34561
rect 10870 34552 10876 34564
rect 10928 34552 10934 34604
rect 12342 34552 12348 34604
rect 12400 34592 12406 34604
rect 12575 34595 12633 34601
rect 12575 34592 12587 34595
rect 12400 34564 12587 34592
rect 12400 34552 12406 34564
rect 12575 34561 12587 34564
rect 12621 34561 12633 34595
rect 12575 34555 12633 34561
rect 4154 34484 4160 34536
rect 4212 34533 4218 34536
rect 4212 34527 4250 34533
rect 4238 34524 4250 34527
rect 4617 34527 4675 34533
rect 4617 34524 4629 34527
rect 4238 34496 4629 34524
rect 4238 34493 4250 34496
rect 4212 34487 4250 34493
rect 4617 34493 4629 34496
rect 4663 34493 4675 34527
rect 4617 34487 4675 34493
rect 5077 34527 5135 34533
rect 5077 34493 5089 34527
rect 5123 34524 5135 34527
rect 5166 34524 5172 34536
rect 5123 34496 5172 34524
rect 5123 34493 5135 34496
rect 5077 34487 5135 34493
rect 4212 34484 4218 34487
rect 5166 34484 5172 34496
rect 5224 34484 5230 34536
rect 5258 34484 5264 34536
rect 5316 34524 5322 34536
rect 5626 34524 5632 34536
rect 5316 34496 5632 34524
rect 5316 34484 5322 34496
rect 5626 34484 5632 34496
rect 5684 34484 5690 34536
rect 5905 34527 5963 34533
rect 5905 34493 5917 34527
rect 5951 34524 5963 34527
rect 6822 34524 6828 34536
rect 5951 34496 6828 34524
rect 5951 34493 5963 34496
rect 5905 34487 5963 34493
rect 6822 34484 6828 34496
rect 6880 34484 6886 34536
rect 9585 34527 9643 34533
rect 9585 34493 9597 34527
rect 9631 34524 9643 34527
rect 9858 34524 9864 34536
rect 9631 34496 9864 34524
rect 9631 34493 9643 34496
rect 9585 34487 9643 34493
rect 9858 34484 9864 34496
rect 9916 34484 9922 34536
rect 11238 34484 11244 34536
rect 11296 34524 11302 34536
rect 11517 34527 11575 34533
rect 11517 34524 11529 34527
rect 11296 34496 11529 34524
rect 11296 34484 11302 34496
rect 11517 34493 11529 34496
rect 11563 34493 11575 34527
rect 11517 34487 11575 34493
rect 12434 34484 12440 34536
rect 12492 34533 12498 34536
rect 12492 34527 12530 34533
rect 12518 34524 12530 34527
rect 12897 34527 12955 34533
rect 12897 34524 12909 34527
rect 12518 34496 12909 34524
rect 12518 34493 12530 34496
rect 12492 34487 12530 34493
rect 12897 34493 12909 34496
rect 12943 34524 12955 34527
rect 13265 34527 13323 34533
rect 13265 34524 13277 34527
rect 12943 34496 13277 34524
rect 12943 34493 12955 34496
rect 12897 34487 12955 34493
rect 13265 34493 13277 34496
rect 13311 34493 13323 34527
rect 13265 34487 13323 34493
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13906 34524 13912 34536
rect 13495 34496 13912 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 12492 34484 12498 34487
rect 13906 34484 13912 34496
rect 13964 34524 13970 34536
rect 14001 34527 14059 34533
rect 14001 34524 14013 34527
rect 13964 34496 14013 34524
rect 13964 34484 13970 34496
rect 14001 34493 14013 34496
rect 14047 34493 14059 34527
rect 14001 34487 14059 34493
rect 9030 34465 9036 34468
rect 7146 34459 7204 34465
rect 7146 34456 7158 34459
rect 6564 34428 7158 34456
rect 6178 34348 6184 34400
rect 6236 34388 6242 34400
rect 6564 34397 6592 34428
rect 7146 34425 7158 34428
rect 7192 34425 7204 34459
rect 9027 34456 9036 34465
rect 8991 34428 9036 34456
rect 7146 34419 7204 34425
rect 9027 34419 9036 34428
rect 9030 34416 9036 34419
rect 9088 34416 9094 34468
rect 10597 34459 10655 34465
rect 10597 34425 10609 34459
rect 10643 34425 10655 34459
rect 10597 34419 10655 34425
rect 6549 34391 6607 34397
rect 6549 34388 6561 34391
rect 6236 34360 6561 34388
rect 6236 34348 6242 34360
rect 6549 34357 6561 34360
rect 6595 34357 6607 34391
rect 10318 34388 10324 34400
rect 10279 34360 10324 34388
rect 6549 34351 6607 34357
rect 10318 34348 10324 34360
rect 10376 34388 10382 34400
rect 10612 34388 10640 34419
rect 10376 34360 10640 34388
rect 10376 34348 10382 34360
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 6914 34144 6920 34196
rect 6972 34184 6978 34196
rect 7377 34187 7435 34193
rect 7377 34184 7389 34187
rect 6972 34156 7389 34184
rect 6972 34144 6978 34156
rect 7377 34153 7389 34156
rect 7423 34153 7435 34187
rect 9398 34184 9404 34196
rect 9359 34156 9404 34184
rect 7377 34147 7435 34153
rect 9398 34144 9404 34156
rect 9456 34144 9462 34196
rect 10597 34187 10655 34193
rect 10597 34153 10609 34187
rect 10643 34184 10655 34187
rect 13538 34184 13544 34196
rect 10643 34156 11652 34184
rect 13499 34156 13544 34184
rect 10643 34153 10655 34156
rect 10597 34147 10655 34153
rect 6178 34125 6184 34128
rect 6175 34116 6184 34125
rect 6139 34088 6184 34116
rect 6175 34079 6184 34088
rect 6178 34076 6184 34079
rect 6236 34076 6242 34128
rect 7006 34116 7012 34128
rect 6967 34088 7012 34116
rect 7006 34076 7012 34088
rect 7064 34076 7070 34128
rect 7745 34119 7803 34125
rect 7745 34116 7757 34119
rect 7208 34088 7757 34116
rect 4522 34008 4528 34060
rect 4580 34048 4586 34060
rect 4836 34051 4894 34057
rect 4836 34048 4848 34051
rect 4580 34020 4848 34048
rect 4580 34008 4586 34020
rect 4836 34017 4848 34020
rect 4882 34017 4894 34051
rect 6730 34048 6736 34060
rect 6643 34020 6736 34048
rect 4836 34011 4894 34017
rect 6730 34008 6736 34020
rect 6788 34048 6794 34060
rect 7208 34048 7236 34088
rect 7745 34085 7757 34088
rect 7791 34116 7803 34119
rect 7834 34116 7840 34128
rect 7791 34088 7840 34116
rect 7791 34085 7803 34088
rect 7745 34079 7803 34085
rect 7834 34076 7840 34088
rect 7892 34076 7898 34128
rect 9030 34116 9036 34128
rect 8680 34088 9036 34116
rect 6788 34020 7236 34048
rect 6788 34008 6794 34020
rect 5813 33983 5871 33989
rect 5813 33949 5825 33983
rect 5859 33980 5871 33983
rect 5902 33980 5908 33992
rect 5859 33952 5908 33980
rect 5859 33949 5871 33952
rect 5813 33943 5871 33949
rect 5902 33940 5908 33952
rect 5960 33940 5966 33992
rect 7653 33983 7711 33989
rect 7653 33949 7665 33983
rect 7699 33949 7711 33983
rect 7926 33980 7932 33992
rect 7887 33952 7932 33980
rect 7653 33943 7711 33949
rect 4939 33915 4997 33921
rect 4939 33881 4951 33915
rect 4985 33912 4997 33915
rect 7668 33912 7696 33943
rect 7926 33940 7932 33952
rect 7984 33940 7990 33992
rect 8294 33912 8300 33924
rect 4985 33884 8300 33912
rect 4985 33881 4997 33884
rect 4939 33875 4997 33881
rect 8294 33872 8300 33884
rect 8352 33872 8358 33924
rect 5258 33844 5264 33856
rect 5219 33816 5264 33844
rect 5258 33804 5264 33816
rect 5316 33804 5322 33856
rect 5534 33804 5540 33856
rect 5592 33844 5598 33856
rect 5629 33847 5687 33853
rect 5629 33844 5641 33847
rect 5592 33816 5641 33844
rect 5592 33804 5598 33816
rect 5629 33813 5641 33816
rect 5675 33813 5687 33847
rect 5629 33807 5687 33813
rect 8202 33804 8208 33856
rect 8260 33844 8266 33856
rect 8680 33853 8708 34088
rect 9030 34076 9036 34088
rect 9088 34116 9094 34128
rect 10039 34119 10097 34125
rect 10039 34116 10051 34119
rect 9088 34088 10051 34116
rect 9088 34076 9094 34088
rect 10039 34085 10051 34088
rect 10085 34116 10097 34119
rect 10134 34116 10140 34128
rect 10085 34088 10140 34116
rect 10085 34085 10097 34088
rect 10039 34079 10097 34085
rect 10134 34076 10140 34088
rect 10192 34076 10198 34128
rect 11054 34076 11060 34128
rect 11112 34116 11118 34128
rect 11514 34116 11520 34128
rect 11112 34088 11520 34116
rect 11112 34076 11118 34088
rect 11514 34076 11520 34088
rect 11572 34076 11578 34128
rect 11624 34125 11652 34156
rect 13538 34144 13544 34156
rect 13596 34144 13602 34196
rect 11609 34119 11667 34125
rect 11609 34085 11621 34119
rect 11655 34116 11667 34119
rect 11698 34116 11704 34128
rect 11655 34088 11704 34116
rect 11655 34085 11667 34088
rect 11609 34079 11667 34085
rect 11698 34076 11704 34088
rect 11756 34076 11762 34128
rect 13357 34051 13415 34057
rect 13357 34017 13369 34051
rect 13403 34048 13415 34051
rect 13538 34048 13544 34060
rect 13403 34020 13544 34048
rect 13403 34017 13415 34020
rect 13357 34011 13415 34017
rect 13538 34008 13544 34020
rect 13596 34008 13602 34060
rect 9674 33980 9680 33992
rect 9635 33952 9680 33980
rect 9674 33940 9680 33952
rect 9732 33940 9738 33992
rect 11974 33980 11980 33992
rect 11935 33952 11980 33980
rect 11974 33940 11980 33952
rect 12032 33940 12038 33992
rect 8665 33847 8723 33853
rect 8665 33844 8677 33847
rect 8260 33816 8677 33844
rect 8260 33804 8266 33816
rect 8665 33813 8677 33816
rect 8711 33813 8723 33847
rect 8665 33807 8723 33813
rect 10502 33804 10508 33856
rect 10560 33844 10566 33856
rect 10873 33847 10931 33853
rect 10873 33844 10885 33847
rect 10560 33816 10885 33844
rect 10560 33804 10566 33816
rect 10873 33813 10885 33816
rect 10919 33813 10931 33847
rect 12526 33844 12532 33856
rect 12487 33816 12532 33844
rect 10873 33807 10931 33813
rect 12526 33804 12532 33816
rect 12584 33804 12590 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 4522 33600 4528 33652
rect 4580 33640 4586 33652
rect 4801 33643 4859 33649
rect 4801 33640 4813 33643
rect 4580 33612 4813 33640
rect 4580 33600 4586 33612
rect 4801 33609 4813 33612
rect 4847 33640 4859 33643
rect 5350 33640 5356 33652
rect 4847 33612 5356 33640
rect 4847 33609 4859 33612
rect 4801 33603 4859 33609
rect 5350 33600 5356 33612
rect 5408 33600 5414 33652
rect 7834 33640 7840 33652
rect 7795 33612 7840 33640
rect 7834 33600 7840 33612
rect 7892 33600 7898 33652
rect 8297 33643 8355 33649
rect 8297 33609 8309 33643
rect 8343 33640 8355 33643
rect 8386 33640 8392 33652
rect 8343 33612 8392 33640
rect 8343 33609 8355 33612
rect 8297 33603 8355 33609
rect 8386 33600 8392 33612
rect 8444 33600 8450 33652
rect 10045 33643 10103 33649
rect 10045 33609 10057 33643
rect 10091 33640 10103 33643
rect 10134 33640 10140 33652
rect 10091 33612 10140 33640
rect 10091 33609 10103 33612
rect 10045 33603 10103 33609
rect 10134 33600 10140 33612
rect 10192 33640 10198 33652
rect 10413 33643 10471 33649
rect 10413 33640 10425 33643
rect 10192 33612 10425 33640
rect 10192 33600 10198 33612
rect 10413 33609 10425 33612
rect 10459 33609 10471 33643
rect 11698 33640 11704 33652
rect 11659 33612 11704 33640
rect 10413 33603 10471 33609
rect 11698 33600 11704 33612
rect 11756 33600 11762 33652
rect 5902 33504 5908 33516
rect 5815 33476 5908 33504
rect 5902 33464 5908 33476
rect 5960 33504 5966 33516
rect 6549 33507 6607 33513
rect 6549 33504 6561 33507
rect 5960 33476 6561 33504
rect 5960 33464 5966 33476
rect 6549 33473 6561 33476
rect 6595 33473 6607 33507
rect 6549 33467 6607 33473
rect 7561 33507 7619 33513
rect 7561 33473 7573 33507
rect 7607 33504 7619 33507
rect 7926 33504 7932 33516
rect 7607 33476 7932 33504
rect 7607 33473 7619 33476
rect 7561 33467 7619 33473
rect 7926 33464 7932 33476
rect 7984 33464 7990 33516
rect 8404 33504 8432 33600
rect 9677 33575 9735 33581
rect 9677 33541 9689 33575
rect 9723 33572 9735 33575
rect 10318 33572 10324 33584
rect 9723 33544 10324 33572
rect 9723 33541 9735 33544
rect 9677 33535 9735 33541
rect 10318 33532 10324 33544
rect 10376 33572 10382 33584
rect 10376 33544 12204 33572
rect 10376 33532 10382 33544
rect 8757 33507 8815 33513
rect 8757 33504 8769 33507
rect 8404 33476 8769 33504
rect 8757 33473 8769 33476
rect 8803 33473 8815 33507
rect 10502 33504 10508 33516
rect 10463 33476 10508 33504
rect 8757 33467 8815 33473
rect 10502 33464 10508 33476
rect 10560 33464 10566 33516
rect 3881 33439 3939 33445
rect 3881 33405 3893 33439
rect 3927 33405 3939 33439
rect 4062 33436 4068 33448
rect 4023 33408 4068 33436
rect 3881 33399 3939 33405
rect 3513 33371 3571 33377
rect 3513 33337 3525 33371
rect 3559 33368 3571 33371
rect 3896 33368 3924 33399
rect 4062 33396 4068 33408
rect 4120 33396 4126 33448
rect 5258 33436 5264 33448
rect 5219 33408 5264 33436
rect 5258 33396 5264 33408
rect 5316 33396 5322 33448
rect 5626 33436 5632 33448
rect 5587 33408 5632 33436
rect 5626 33396 5632 33408
rect 5684 33396 5690 33448
rect 5166 33368 5172 33380
rect 3559 33340 5172 33368
rect 3559 33337 3571 33340
rect 3513 33331 3571 33337
rect 5166 33328 5172 33340
rect 5224 33328 5230 33380
rect 5534 33328 5540 33380
rect 5592 33368 5598 33380
rect 6917 33371 6975 33377
rect 6917 33368 6929 33371
rect 5592 33340 6929 33368
rect 5592 33328 5598 33340
rect 6917 33337 6929 33340
rect 6963 33337 6975 33371
rect 6917 33331 6975 33337
rect 7006 33328 7012 33380
rect 7064 33368 7070 33380
rect 8665 33371 8723 33377
rect 7064 33340 7109 33368
rect 7064 33328 7070 33340
rect 8665 33337 8677 33371
rect 8711 33368 8723 33371
rect 9078 33371 9136 33377
rect 9078 33368 9090 33371
rect 8711 33340 9090 33368
rect 8711 33337 8723 33340
rect 8665 33331 8723 33337
rect 9078 33337 9090 33340
rect 9124 33368 9136 33371
rect 10134 33368 10140 33380
rect 9124 33340 10140 33368
rect 9124 33337 9136 33340
rect 9078 33331 9136 33337
rect 10134 33328 10140 33340
rect 10192 33368 10198 33380
rect 10826 33371 10884 33377
rect 10826 33368 10838 33371
rect 10192 33340 10838 33368
rect 10192 33328 10198 33340
rect 10826 33337 10838 33340
rect 10872 33337 10884 33371
rect 10826 33331 10884 33337
rect 3878 33300 3884 33312
rect 3839 33272 3884 33300
rect 3878 33260 3884 33272
rect 3936 33260 3942 33312
rect 6178 33300 6184 33312
rect 6139 33272 6184 33300
rect 6178 33260 6184 33272
rect 6236 33260 6242 33312
rect 11422 33300 11428 33312
rect 11383 33272 11428 33300
rect 11422 33260 11428 33272
rect 11480 33260 11486 33312
rect 12176 33309 12204 33544
rect 12250 33464 12256 33516
rect 12308 33504 12314 33516
rect 12805 33507 12863 33513
rect 12805 33504 12817 33507
rect 12308 33476 12817 33504
rect 12308 33464 12314 33476
rect 12805 33473 12817 33476
rect 12851 33473 12863 33507
rect 12805 33467 12863 33473
rect 12250 33328 12256 33380
rect 12308 33368 12314 33380
rect 12526 33368 12532 33380
rect 12308 33340 12532 33368
rect 12308 33328 12314 33340
rect 12526 33328 12532 33340
rect 12584 33328 12590 33380
rect 12621 33371 12679 33377
rect 12621 33337 12633 33371
rect 12667 33337 12679 33371
rect 12621 33331 12679 33337
rect 12161 33303 12219 33309
rect 12161 33269 12173 33303
rect 12207 33300 12219 33303
rect 12636 33300 12664 33331
rect 13538 33300 13544 33312
rect 12207 33272 12664 33300
rect 13499 33272 13544 33300
rect 12207 33269 12219 33272
rect 12161 33263 12219 33269
rect 13538 33260 13544 33272
rect 13596 33260 13602 33312
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 3697 33099 3755 33105
rect 3697 33065 3709 33099
rect 3743 33096 3755 33099
rect 4062 33096 4068 33108
rect 3743 33068 4068 33096
rect 3743 33065 3755 33068
rect 3697 33059 3755 33065
rect 4062 33056 4068 33068
rect 4120 33056 4126 33108
rect 4847 33099 4905 33105
rect 4847 33065 4859 33099
rect 4893 33096 4905 33099
rect 5442 33096 5448 33108
rect 4893 33068 5448 33096
rect 4893 33065 4905 33068
rect 4847 33059 4905 33065
rect 5442 33056 5448 33068
rect 5500 33056 5506 33108
rect 5626 33096 5632 33108
rect 5587 33068 5632 33096
rect 5626 33056 5632 33068
rect 5684 33056 5690 33108
rect 8294 33056 8300 33108
rect 8352 33096 8358 33108
rect 8849 33099 8907 33105
rect 8849 33096 8861 33099
rect 8352 33068 8861 33096
rect 8352 33056 8358 33068
rect 8849 33065 8861 33068
rect 8895 33065 8907 33099
rect 8849 33059 8907 33065
rect 9674 33056 9680 33108
rect 9732 33096 9738 33108
rect 9861 33099 9919 33105
rect 9861 33096 9873 33099
rect 9732 33068 9873 33096
rect 9732 33056 9738 33068
rect 9861 33065 9873 33068
rect 9907 33065 9919 33099
rect 11514 33096 11520 33108
rect 11475 33068 11520 33096
rect 9861 33059 9919 33065
rect 11514 33056 11520 33068
rect 11572 33056 11578 33108
rect 12342 33096 12348 33108
rect 11808 33068 12348 33096
rect 6083 33031 6141 33037
rect 6083 32997 6095 33031
rect 6129 33028 6141 33031
rect 6178 33028 6184 33040
rect 6129 33000 6184 33028
rect 6129 32997 6141 33000
rect 6083 32991 6141 32997
rect 6178 32988 6184 33000
rect 6236 32988 6242 33040
rect 8018 33028 8024 33040
rect 7979 33000 8024 33028
rect 8018 32988 8024 33000
rect 8076 32988 8082 33040
rect 10318 33028 10324 33040
rect 10279 33000 10324 33028
rect 10318 32988 10324 33000
rect 10376 32988 10382 33040
rect 10870 33028 10876 33040
rect 10831 33000 10876 33028
rect 10870 32988 10876 33000
rect 10928 32988 10934 33040
rect 11808 33037 11836 33068
rect 12342 33056 12348 33068
rect 12400 33056 12406 33108
rect 11793 33031 11851 33037
rect 11793 32997 11805 33031
rect 11839 32997 11851 33031
rect 11793 32991 11851 32997
rect 11882 32988 11888 33040
rect 11940 33028 11946 33040
rect 11940 33000 11985 33028
rect 11940 32988 11946 33000
rect 4338 32920 4344 32972
rect 4396 32960 4402 32972
rect 4744 32963 4802 32969
rect 4744 32960 4756 32963
rect 4396 32932 4756 32960
rect 4396 32920 4402 32932
rect 4744 32929 4756 32932
rect 4790 32960 4802 32963
rect 4982 32960 4988 32972
rect 4790 32932 4988 32960
rect 4790 32929 4802 32932
rect 4744 32923 4802 32929
rect 4982 32920 4988 32932
rect 5040 32920 5046 32972
rect 13332 32963 13390 32969
rect 13332 32929 13344 32963
rect 13378 32960 13390 32963
rect 13538 32960 13544 32972
rect 13378 32932 13544 32960
rect 13378 32929 13390 32932
rect 13332 32923 13390 32929
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32892 5779 32895
rect 6086 32892 6092 32904
rect 5767 32864 6092 32892
rect 5767 32861 5779 32864
rect 5721 32855 5779 32861
rect 6086 32852 6092 32864
rect 6144 32852 6150 32904
rect 7742 32852 7748 32904
rect 7800 32892 7806 32904
rect 7929 32895 7987 32901
rect 7929 32892 7941 32895
rect 7800 32864 7941 32892
rect 7800 32852 7806 32864
rect 7929 32861 7941 32864
rect 7975 32861 7987 32895
rect 8294 32892 8300 32904
rect 8255 32864 8300 32892
rect 7929 32855 7987 32861
rect 8294 32852 8300 32864
rect 8352 32852 8358 32904
rect 9582 32852 9588 32904
rect 9640 32892 9646 32904
rect 10229 32895 10287 32901
rect 10229 32892 10241 32895
rect 9640 32864 10241 32892
rect 9640 32852 9646 32864
rect 10229 32861 10241 32864
rect 10275 32861 10287 32895
rect 10229 32855 10287 32861
rect 11514 32852 11520 32904
rect 11572 32892 11578 32904
rect 12069 32895 12127 32901
rect 12069 32892 12081 32895
rect 11572 32864 12081 32892
rect 11572 32852 11578 32864
rect 12069 32861 12081 32864
rect 12115 32892 12127 32895
rect 12158 32892 12164 32904
rect 12115 32864 12164 32892
rect 12115 32861 12127 32864
rect 12069 32855 12127 32861
rect 12158 32852 12164 32864
rect 12216 32852 12222 32904
rect 5166 32756 5172 32768
rect 5127 32728 5172 32756
rect 5166 32716 5172 32728
rect 5224 32716 5230 32768
rect 6641 32759 6699 32765
rect 6641 32725 6653 32759
rect 6687 32756 6699 32759
rect 7006 32756 7012 32768
rect 6687 32728 7012 32756
rect 6687 32725 6699 32728
rect 6641 32719 6699 32725
rect 7006 32716 7012 32728
rect 7064 32716 7070 32768
rect 7374 32756 7380 32768
rect 7335 32728 7380 32756
rect 7374 32716 7380 32728
rect 7432 32716 7438 32768
rect 12894 32716 12900 32768
rect 12952 32756 12958 32768
rect 13403 32759 13461 32765
rect 13403 32756 13415 32759
rect 12952 32728 13415 32756
rect 12952 32716 12958 32728
rect 13403 32725 13415 32728
rect 13449 32725 13461 32759
rect 13403 32719 13461 32725
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 4982 32552 4988 32564
rect 4943 32524 4988 32552
rect 4982 32512 4988 32524
rect 5040 32512 5046 32564
rect 8018 32512 8024 32564
rect 8076 32552 8082 32564
rect 8297 32555 8355 32561
rect 8297 32552 8309 32555
rect 8076 32524 8309 32552
rect 8076 32512 8082 32524
rect 8297 32521 8309 32524
rect 8343 32552 8355 32555
rect 8573 32555 8631 32561
rect 8573 32552 8585 32555
rect 8343 32524 8585 32552
rect 8343 32521 8355 32524
rect 8297 32515 8355 32521
rect 8573 32521 8585 32524
rect 8619 32521 8631 32555
rect 8573 32515 8631 32521
rect 10318 32512 10324 32564
rect 10376 32552 10382 32564
rect 10965 32555 11023 32561
rect 10965 32552 10977 32555
rect 10376 32524 10977 32552
rect 10376 32512 10382 32524
rect 10965 32521 10977 32524
rect 11011 32552 11023 32555
rect 11422 32552 11428 32564
rect 11011 32524 11428 32552
rect 11011 32521 11023 32524
rect 10965 32515 11023 32521
rect 11422 32512 11428 32524
rect 11480 32552 11486 32564
rect 11701 32555 11759 32561
rect 11701 32552 11713 32555
rect 11480 32524 11713 32552
rect 11480 32512 11486 32524
rect 11701 32521 11713 32524
rect 11747 32552 11759 32555
rect 11882 32552 11888 32564
rect 11747 32524 11888 32552
rect 11747 32521 11759 32524
rect 11701 32515 11759 32521
rect 11882 32512 11888 32524
rect 11940 32512 11946 32564
rect 12161 32555 12219 32561
rect 12161 32521 12173 32555
rect 12207 32552 12219 32555
rect 12342 32552 12348 32564
rect 12207 32524 12348 32552
rect 12207 32521 12219 32524
rect 12161 32515 12219 32521
rect 12342 32512 12348 32524
rect 12400 32512 12406 32564
rect 12618 32561 12624 32564
rect 12575 32555 12624 32561
rect 12575 32521 12587 32555
rect 12621 32521 12624 32555
rect 12575 32515 12624 32521
rect 12618 32512 12624 32515
rect 12676 32512 12682 32564
rect 6549 32419 6607 32425
rect 6549 32416 6561 32419
rect 5644 32388 6561 32416
rect 5644 32360 5672 32388
rect 6549 32385 6561 32388
rect 6595 32385 6607 32419
rect 6549 32379 6607 32385
rect 9493 32419 9551 32425
rect 9493 32385 9505 32419
rect 9539 32416 9551 32419
rect 10042 32416 10048 32428
rect 9539 32388 10048 32416
rect 9539 32385 9551 32388
rect 9493 32379 9551 32385
rect 10042 32376 10048 32388
rect 10100 32376 10106 32428
rect 10689 32419 10747 32425
rect 10689 32385 10701 32419
rect 10735 32416 10747 32419
rect 10870 32416 10876 32428
rect 10735 32388 10876 32416
rect 10735 32385 10747 32388
rect 10689 32379 10747 32385
rect 10870 32376 10876 32388
rect 10928 32376 10934 32428
rect 4224 32351 4282 32357
rect 4224 32317 4236 32351
rect 4270 32348 4282 32351
rect 4522 32348 4528 32360
rect 4270 32320 4528 32348
rect 4270 32317 4282 32320
rect 4224 32311 4282 32317
rect 4522 32308 4528 32320
rect 4580 32348 4586 32360
rect 4617 32351 4675 32357
rect 4617 32348 4629 32351
rect 4580 32320 4629 32348
rect 4580 32308 4586 32320
rect 4617 32317 4629 32320
rect 4663 32317 4675 32351
rect 5166 32348 5172 32360
rect 5127 32320 5172 32348
rect 4617 32311 4675 32317
rect 5166 32308 5172 32320
rect 5224 32308 5230 32360
rect 5626 32348 5632 32360
rect 5587 32320 5632 32348
rect 5626 32308 5632 32320
rect 5684 32308 5690 32360
rect 5994 32308 6000 32360
rect 6052 32348 6058 32360
rect 7374 32348 7380 32360
rect 6052 32320 7380 32348
rect 6052 32308 6058 32320
rect 7374 32308 7380 32320
rect 7432 32308 7438 32360
rect 12434 32308 12440 32360
rect 12492 32357 12498 32360
rect 12492 32351 12530 32357
rect 12518 32348 12530 32351
rect 12897 32351 12955 32357
rect 12897 32348 12909 32351
rect 12518 32320 12909 32348
rect 12518 32317 12530 32320
rect 12492 32311 12530 32317
rect 12897 32317 12909 32320
rect 12943 32317 12955 32351
rect 12897 32311 12955 32317
rect 12492 32308 12498 32311
rect 5905 32283 5963 32289
rect 5905 32249 5917 32283
rect 5951 32280 5963 32283
rect 6086 32280 6092 32292
rect 5951 32252 6092 32280
rect 5951 32249 5963 32252
rect 5905 32243 5963 32249
rect 6086 32240 6092 32252
rect 6144 32240 6150 32292
rect 7699 32283 7757 32289
rect 7699 32249 7711 32283
rect 7745 32280 7757 32283
rect 8202 32280 8208 32292
rect 7745 32252 8208 32280
rect 7745 32249 7757 32252
rect 7699 32243 7757 32249
rect 4295 32215 4353 32221
rect 4295 32181 4307 32215
rect 4341 32212 4353 32215
rect 5534 32212 5540 32224
rect 4341 32184 5540 32212
rect 4341 32181 4353 32184
rect 4295 32175 4353 32181
rect 5534 32172 5540 32184
rect 5592 32172 5598 32224
rect 6178 32172 6184 32224
rect 6236 32212 6242 32224
rect 6273 32215 6331 32221
rect 6273 32212 6285 32215
rect 6236 32184 6285 32212
rect 6236 32172 6242 32184
rect 6273 32181 6285 32184
rect 6319 32212 6331 32215
rect 7098 32212 7104 32224
rect 6319 32184 7104 32212
rect 6319 32181 6331 32184
rect 6273 32175 6331 32181
rect 7098 32172 7104 32184
rect 7156 32212 7162 32224
rect 7193 32215 7251 32221
rect 7193 32212 7205 32215
rect 7156 32184 7205 32212
rect 7156 32172 7162 32184
rect 7193 32181 7205 32184
rect 7239 32212 7251 32215
rect 7713 32212 7741 32243
rect 8202 32240 8208 32252
rect 8260 32240 8266 32292
rect 9858 32280 9864 32292
rect 9771 32252 9864 32280
rect 9858 32240 9864 32252
rect 9916 32280 9922 32292
rect 10137 32283 10195 32289
rect 10137 32280 10149 32283
rect 9916 32252 10149 32280
rect 9916 32240 9922 32252
rect 10137 32249 10149 32252
rect 10183 32249 10195 32283
rect 10137 32243 10195 32249
rect 7239 32184 7741 32212
rect 7239 32181 7251 32184
rect 7193 32175 7251 32181
rect 9582 32172 9588 32224
rect 9640 32212 9646 32224
rect 11333 32215 11391 32221
rect 11333 32212 11345 32215
rect 9640 32184 11345 32212
rect 9640 32172 9646 32184
rect 11333 32181 11345 32184
rect 11379 32181 11391 32215
rect 11333 32175 11391 32181
rect 13357 32215 13415 32221
rect 13357 32181 13369 32215
rect 13403 32212 13415 32215
rect 13538 32212 13544 32224
rect 13403 32184 13544 32212
rect 13403 32181 13415 32184
rect 13357 32175 13415 32181
rect 13538 32172 13544 32184
rect 13596 32172 13602 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 6086 31968 6092 32020
rect 6144 32008 6150 32020
rect 6273 32011 6331 32017
rect 6273 32008 6285 32011
rect 6144 31980 6285 32008
rect 6144 31968 6150 31980
rect 6273 31977 6285 31980
rect 6319 31977 6331 32011
rect 7742 32008 7748 32020
rect 6273 31971 6331 31977
rect 7576 31980 7748 32008
rect 5994 31940 6000 31952
rect 5955 31912 6000 31940
rect 5994 31900 6000 31912
rect 6052 31900 6058 31952
rect 7006 31940 7012 31952
rect 6967 31912 7012 31940
rect 7006 31900 7012 31912
rect 7064 31900 7070 31952
rect 7576 31949 7604 31980
rect 7742 31968 7748 31980
rect 7800 32008 7806 32020
rect 7837 32011 7895 32017
rect 7837 32008 7849 32011
rect 7800 31980 7849 32008
rect 7800 31968 7806 31980
rect 7837 31977 7849 31980
rect 7883 31977 7895 32011
rect 7837 31971 7895 31977
rect 7926 31968 7932 32020
rect 7984 32008 7990 32020
rect 8205 32011 8263 32017
rect 8205 32008 8217 32011
rect 7984 31980 8217 32008
rect 7984 31968 7990 31980
rect 8205 31977 8217 31980
rect 8251 31977 8263 32011
rect 8205 31971 8263 31977
rect 8711 32011 8769 32017
rect 8711 31977 8723 32011
rect 8757 32008 8769 32011
rect 9582 32008 9588 32020
rect 8757 31980 9588 32008
rect 8757 31977 8769 31980
rect 8711 31971 8769 31977
rect 9582 31968 9588 31980
rect 9640 31968 9646 32020
rect 9674 31968 9680 32020
rect 9732 32008 9738 32020
rect 9769 32011 9827 32017
rect 9769 32008 9781 32011
rect 9732 31980 9781 32008
rect 9732 31968 9738 31980
rect 9769 31977 9781 31980
rect 9815 31977 9827 32011
rect 9769 31971 9827 31977
rect 11379 32011 11437 32017
rect 11379 31977 11391 32011
rect 11425 32008 11437 32011
rect 12250 32008 12256 32020
rect 11425 31980 12256 32008
rect 11425 31977 11437 31980
rect 11379 31971 11437 31977
rect 12250 31968 12256 31980
rect 12308 31968 12314 32020
rect 7561 31943 7619 31949
rect 7561 31909 7573 31943
rect 7607 31909 7619 31943
rect 7561 31903 7619 31909
rect 4062 31832 4068 31884
rect 4120 31881 4126 31884
rect 4120 31875 4158 31881
rect 4146 31841 4158 31875
rect 5442 31872 5448 31884
rect 5403 31844 5448 31872
rect 4120 31835 4158 31841
rect 4120 31832 4126 31835
rect 5442 31832 5448 31844
rect 5500 31832 5506 31884
rect 5626 31832 5632 31884
rect 5684 31872 5690 31884
rect 5721 31875 5779 31881
rect 5721 31872 5733 31875
rect 5684 31844 5733 31872
rect 5684 31832 5690 31844
rect 5721 31841 5733 31844
rect 5767 31841 5779 31875
rect 5721 31835 5779 31841
rect 8640 31875 8698 31881
rect 8640 31841 8652 31875
rect 8686 31872 8698 31875
rect 8754 31872 8760 31884
rect 8686 31844 8760 31872
rect 8686 31841 8698 31844
rect 8640 31835 8698 31841
rect 8754 31832 8760 31844
rect 8812 31832 8818 31884
rect 9950 31872 9956 31884
rect 9911 31844 9956 31872
rect 9950 31832 9956 31844
rect 10008 31832 10014 31884
rect 10137 31875 10195 31881
rect 10137 31841 10149 31875
rect 10183 31841 10195 31875
rect 10137 31835 10195 31841
rect 4246 31813 4252 31816
rect 4203 31807 4252 31813
rect 4203 31773 4215 31807
rect 4249 31773 4252 31807
rect 4203 31767 4252 31773
rect 4246 31764 4252 31767
rect 4304 31764 4310 31816
rect 6906 31807 6964 31813
rect 6906 31773 6918 31807
rect 6952 31773 6964 31807
rect 10152 31804 10180 31835
rect 11146 31832 11152 31884
rect 11204 31872 11210 31884
rect 11308 31875 11366 31881
rect 11308 31872 11320 31875
rect 11204 31844 11320 31872
rect 11204 31832 11210 31844
rect 11308 31841 11320 31844
rect 11354 31872 11366 31875
rect 12158 31872 12164 31884
rect 11354 31844 12164 31872
rect 11354 31841 11366 31844
rect 11308 31835 11366 31841
rect 12158 31832 12164 31844
rect 12216 31832 12222 31884
rect 6906 31767 6964 31773
rect 9508 31776 10180 31804
rect 5534 31696 5540 31748
rect 5592 31736 5598 31748
rect 6546 31736 6552 31748
rect 5592 31708 6552 31736
rect 5592 31696 5598 31708
rect 6546 31696 6552 31708
rect 6604 31736 6610 31748
rect 6932 31736 6960 31767
rect 6604 31708 6960 31736
rect 6604 31696 6610 31708
rect 9508 31680 9536 31776
rect 9125 31671 9183 31677
rect 9125 31637 9137 31671
rect 9171 31668 9183 31671
rect 9490 31668 9496 31680
rect 9171 31640 9496 31668
rect 9171 31637 9183 31640
rect 9125 31631 9183 31637
rect 9490 31628 9496 31640
rect 9548 31628 9554 31680
rect 10594 31628 10600 31680
rect 10652 31668 10658 31680
rect 10689 31671 10747 31677
rect 10689 31668 10701 31671
rect 10652 31640 10701 31668
rect 10652 31628 10658 31640
rect 10689 31637 10701 31640
rect 10735 31637 10747 31671
rect 10689 31631 10747 31637
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 5718 31464 5724 31476
rect 5679 31436 5724 31464
rect 5718 31424 5724 31436
rect 5776 31424 5782 31476
rect 6546 31464 6552 31476
rect 6507 31436 6552 31464
rect 6546 31424 6552 31436
rect 6604 31424 6610 31476
rect 7006 31464 7012 31476
rect 6967 31436 7012 31464
rect 7006 31424 7012 31436
rect 7064 31424 7070 31476
rect 8113 31399 8171 31405
rect 8113 31365 8125 31399
rect 8159 31396 8171 31399
rect 8294 31396 8300 31408
rect 8159 31368 8300 31396
rect 8159 31365 8171 31368
rect 8113 31359 8171 31365
rect 8294 31356 8300 31368
rect 8352 31356 8358 31408
rect 7561 31331 7619 31337
rect 7561 31297 7573 31331
rect 7607 31328 7619 31331
rect 7926 31328 7932 31340
rect 7607 31300 7932 31328
rect 7607 31297 7619 31300
rect 7561 31291 7619 31297
rect 7926 31288 7932 31300
rect 7984 31288 7990 31340
rect 9582 31328 9588 31340
rect 9543 31300 9588 31328
rect 9582 31288 9588 31300
rect 9640 31288 9646 31340
rect 10778 31328 10784 31340
rect 10739 31300 10784 31328
rect 10778 31288 10784 31300
rect 10836 31288 10842 31340
rect 11425 31331 11483 31337
rect 11425 31297 11437 31331
rect 11471 31328 11483 31331
rect 11974 31328 11980 31340
rect 11471 31300 11980 31328
rect 11471 31297 11483 31300
rect 11425 31291 11483 31297
rect 11974 31288 11980 31300
rect 12032 31288 12038 31340
rect 4525 31263 4583 31269
rect 4525 31229 4537 31263
rect 4571 31260 4583 31263
rect 5166 31260 5172 31272
rect 4571 31232 5172 31260
rect 4571 31229 4583 31232
rect 4525 31223 4583 31229
rect 5166 31220 5172 31232
rect 5224 31220 5230 31272
rect 9030 31260 9036 31272
rect 8991 31232 9036 31260
rect 9030 31220 9036 31232
rect 9088 31220 9094 31272
rect 9490 31260 9496 31272
rect 9403 31232 9496 31260
rect 9490 31220 9496 31232
rect 9548 31260 9554 31272
rect 9548 31232 9812 31260
rect 9548 31220 9554 31232
rect 4062 31152 4068 31204
rect 4120 31192 4126 31204
rect 4157 31195 4215 31201
rect 4157 31192 4169 31195
rect 4120 31164 4169 31192
rect 4120 31152 4126 31164
rect 4157 31161 4169 31164
rect 4203 31192 4215 31195
rect 5350 31192 5356 31204
rect 4203 31164 5356 31192
rect 4203 31161 4215 31164
rect 4157 31155 4215 31161
rect 5350 31152 5356 31164
rect 5408 31152 5414 31204
rect 7653 31195 7711 31201
rect 7653 31161 7665 31195
rect 7699 31192 7711 31195
rect 7742 31192 7748 31204
rect 7699 31164 7748 31192
rect 7699 31161 7711 31164
rect 7653 31155 7711 31161
rect 7742 31152 7748 31164
rect 7800 31152 7806 31204
rect 9784 31136 9812 31232
rect 9950 31152 9956 31204
rect 10008 31192 10014 31204
rect 10413 31195 10471 31201
rect 10413 31192 10425 31195
rect 10008 31164 10425 31192
rect 10008 31152 10014 31164
rect 10413 31161 10425 31164
rect 10459 31161 10471 31195
rect 10413 31155 10471 31161
rect 10594 31152 10600 31204
rect 10652 31192 10658 31204
rect 10873 31195 10931 31201
rect 10873 31192 10885 31195
rect 10652 31164 10885 31192
rect 10652 31152 10658 31164
rect 10873 31161 10885 31164
rect 10919 31161 10931 31195
rect 10873 31155 10931 31161
rect 4890 31124 4896 31136
rect 4851 31096 4896 31124
rect 4890 31084 4896 31096
rect 4948 31084 4954 31136
rect 5442 31084 5448 31136
rect 5500 31124 5506 31136
rect 6086 31124 6092 31136
rect 5500 31096 6092 31124
rect 5500 31084 5506 31096
rect 6086 31084 6092 31096
rect 6144 31084 6150 31136
rect 8665 31127 8723 31133
rect 8665 31093 8677 31127
rect 8711 31124 8723 31127
rect 8754 31124 8760 31136
rect 8711 31096 8760 31124
rect 8711 31093 8723 31096
rect 8665 31087 8723 31093
rect 8754 31084 8760 31096
rect 8812 31084 8818 31136
rect 9766 31084 9772 31136
rect 9824 31124 9830 31136
rect 10045 31127 10103 31133
rect 10045 31124 10057 31127
rect 9824 31096 10057 31124
rect 9824 31084 9830 31096
rect 10045 31093 10057 31096
rect 10091 31093 10103 31127
rect 10045 31087 10103 31093
rect 11793 31127 11851 31133
rect 11793 31093 11805 31127
rect 11839 31124 11851 31127
rect 12158 31124 12164 31136
rect 11839 31096 12164 31124
rect 11839 31093 11851 31096
rect 11793 31087 11851 31093
rect 12158 31084 12164 31096
rect 12216 31084 12222 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 7006 30880 7012 30932
rect 7064 30920 7070 30932
rect 9030 30920 9036 30932
rect 7064 30892 9036 30920
rect 7064 30880 7070 30892
rect 9030 30880 9036 30892
rect 9088 30880 9094 30932
rect 10594 30920 10600 30932
rect 10555 30892 10600 30920
rect 10594 30880 10600 30892
rect 10652 30880 10658 30932
rect 10778 30880 10784 30932
rect 10836 30920 10842 30932
rect 10873 30923 10931 30929
rect 10873 30920 10885 30923
rect 10836 30892 10885 30920
rect 10836 30880 10842 30892
rect 10873 30889 10885 30892
rect 10919 30889 10931 30923
rect 10873 30883 10931 30889
rect 4801 30855 4859 30861
rect 4801 30821 4813 30855
rect 4847 30852 4859 30855
rect 4890 30852 4896 30864
rect 4847 30824 4896 30852
rect 4847 30821 4859 30824
rect 4801 30815 4859 30821
rect 4890 30812 4896 30824
rect 4948 30812 4954 30864
rect 7834 30852 7840 30864
rect 7795 30824 7840 30852
rect 7834 30812 7840 30824
rect 7892 30812 7898 30864
rect 10039 30855 10097 30861
rect 10039 30821 10051 30855
rect 10085 30852 10097 30855
rect 10134 30852 10140 30864
rect 10085 30824 10140 30852
rect 10085 30821 10097 30824
rect 10039 30815 10097 30821
rect 10134 30812 10140 30824
rect 10192 30812 10198 30864
rect 11606 30852 11612 30864
rect 11567 30824 11612 30852
rect 11606 30812 11612 30824
rect 11664 30812 11670 30864
rect 5626 30744 5632 30796
rect 5684 30784 5690 30796
rect 5810 30784 5816 30796
rect 5684 30756 5816 30784
rect 5684 30744 5690 30756
rect 5810 30744 5816 30756
rect 5868 30744 5874 30796
rect 6178 30744 6184 30796
rect 6236 30784 6242 30796
rect 6273 30787 6331 30793
rect 6273 30784 6285 30787
rect 6236 30756 6285 30784
rect 6236 30744 6242 30756
rect 6273 30753 6285 30756
rect 6319 30753 6331 30787
rect 6454 30784 6460 30796
rect 6415 30756 6460 30784
rect 6273 30747 6331 30753
rect 6454 30744 6460 30756
rect 6512 30744 6518 30796
rect 4062 30676 4068 30728
rect 4120 30716 4126 30728
rect 4709 30719 4767 30725
rect 4709 30716 4721 30719
rect 4120 30688 4721 30716
rect 4120 30676 4126 30688
rect 4709 30685 4721 30688
rect 4755 30685 4767 30719
rect 5350 30716 5356 30728
rect 5311 30688 5356 30716
rect 4709 30679 4767 30685
rect 5350 30676 5356 30688
rect 5408 30676 5414 30728
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30716 7803 30719
rect 8018 30716 8024 30728
rect 7791 30688 8024 30716
rect 7791 30685 7803 30688
rect 7745 30679 7803 30685
rect 8018 30676 8024 30688
rect 8076 30676 8082 30728
rect 9674 30716 9680 30728
rect 9635 30688 9680 30716
rect 9674 30676 9680 30688
rect 9732 30676 9738 30728
rect 11514 30716 11520 30728
rect 11475 30688 11520 30716
rect 11514 30676 11520 30688
rect 11572 30676 11578 30728
rect 11974 30716 11980 30728
rect 11935 30688 11980 30716
rect 11974 30676 11980 30688
rect 12032 30676 12038 30728
rect 5442 30608 5448 30660
rect 5500 30648 5506 30660
rect 8294 30648 8300 30660
rect 5500 30620 6592 30648
rect 8255 30620 8300 30648
rect 5500 30608 5506 30620
rect 5166 30540 5172 30592
rect 5224 30580 5230 30592
rect 5721 30583 5779 30589
rect 5721 30580 5733 30583
rect 5224 30552 5733 30580
rect 5224 30540 5230 30552
rect 5721 30549 5733 30552
rect 5767 30580 5779 30583
rect 5902 30580 5908 30592
rect 5767 30552 5908 30580
rect 5767 30549 5779 30552
rect 5721 30543 5779 30549
rect 5902 30540 5908 30552
rect 5960 30540 5966 30592
rect 6564 30589 6592 30620
rect 8294 30608 8300 30620
rect 8352 30648 8358 30660
rect 8665 30651 8723 30657
rect 8665 30648 8677 30651
rect 8352 30620 8677 30648
rect 8352 30608 8358 30620
rect 8665 30617 8677 30620
rect 8711 30617 8723 30651
rect 8665 30611 8723 30617
rect 6549 30583 6607 30589
rect 6549 30549 6561 30583
rect 6595 30549 6607 30583
rect 7098 30580 7104 30592
rect 7059 30552 7104 30580
rect 6549 30543 6607 30549
rect 7098 30540 7104 30552
rect 7156 30540 7162 30592
rect 7561 30583 7619 30589
rect 7561 30549 7573 30583
rect 7607 30580 7619 30583
rect 7742 30580 7748 30592
rect 7607 30552 7748 30580
rect 7607 30549 7619 30552
rect 7561 30543 7619 30549
rect 7742 30540 7748 30552
rect 7800 30540 7806 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 4709 30379 4767 30385
rect 4709 30345 4721 30379
rect 4755 30376 4767 30379
rect 4890 30376 4896 30388
rect 4755 30348 4896 30376
rect 4755 30345 4767 30348
rect 4709 30339 4767 30345
rect 4890 30336 4896 30348
rect 4948 30336 4954 30388
rect 6365 30379 6423 30385
rect 6365 30345 6377 30379
rect 6411 30376 6423 30379
rect 6454 30376 6460 30388
rect 6411 30348 6460 30376
rect 6411 30345 6423 30348
rect 6365 30339 6423 30345
rect 6454 30336 6460 30348
rect 6512 30336 6518 30388
rect 7742 30376 7748 30388
rect 7703 30348 7748 30376
rect 7742 30336 7748 30348
rect 7800 30336 7806 30388
rect 8018 30376 8024 30388
rect 7979 30348 8024 30376
rect 8018 30336 8024 30348
rect 8076 30336 8082 30388
rect 11514 30376 11520 30388
rect 11475 30348 11520 30376
rect 11514 30336 11520 30348
rect 11572 30336 11578 30388
rect 3881 30311 3939 30317
rect 3881 30277 3893 30311
rect 3927 30308 3939 30311
rect 4062 30308 4068 30320
rect 3927 30280 4068 30308
rect 3927 30277 3939 30280
rect 3881 30271 3939 30277
rect 3988 30249 4016 30280
rect 4062 30268 4068 30280
rect 4120 30268 4126 30320
rect 8846 30317 8852 30320
rect 8803 30311 8852 30317
rect 8803 30277 8815 30311
rect 8849 30277 8852 30311
rect 8803 30271 8852 30277
rect 8846 30268 8852 30271
rect 8904 30268 8910 30320
rect 10597 30311 10655 30317
rect 10597 30277 10609 30311
rect 10643 30308 10655 30311
rect 11606 30308 11612 30320
rect 10643 30280 11612 30308
rect 10643 30277 10655 30280
rect 10597 30271 10655 30277
rect 11606 30268 11612 30280
rect 11664 30308 11670 30320
rect 11793 30311 11851 30317
rect 11793 30308 11805 30311
rect 11664 30280 11805 30308
rect 11664 30268 11670 30280
rect 11793 30277 11805 30280
rect 11839 30277 11851 30311
rect 11793 30271 11851 30277
rect 3973 30243 4031 30249
rect 3973 30209 3985 30243
rect 4019 30240 4031 30243
rect 5350 30240 5356 30252
rect 4019 30212 4053 30240
rect 5311 30212 5356 30240
rect 4019 30209 4031 30212
rect 3973 30203 4031 30209
rect 5350 30200 5356 30212
rect 5408 30200 5414 30252
rect 9582 30200 9588 30252
rect 9640 30240 9646 30252
rect 9677 30243 9735 30249
rect 9677 30240 9689 30243
rect 9640 30212 9689 30240
rect 9640 30200 9646 30212
rect 9677 30209 9689 30212
rect 9723 30209 9735 30243
rect 9677 30203 9735 30209
rect 6822 30172 6828 30184
rect 6783 30144 6828 30172
rect 6822 30132 6828 30144
rect 6880 30132 6886 30184
rect 8294 30132 8300 30184
rect 8352 30172 8358 30184
rect 8700 30175 8758 30181
rect 8700 30172 8712 30175
rect 8352 30144 8712 30172
rect 8352 30132 8358 30144
rect 8700 30141 8712 30144
rect 8746 30141 8758 30175
rect 8700 30135 8758 30141
rect 5074 30104 5080 30116
rect 5035 30076 5080 30104
rect 5074 30064 5080 30076
rect 5132 30064 5138 30116
rect 5166 30064 5172 30116
rect 5224 30104 5230 30116
rect 5224 30076 5269 30104
rect 5224 30064 5230 30076
rect 7098 30064 7104 30116
rect 7156 30113 7162 30116
rect 7156 30107 7204 30113
rect 7156 30073 7158 30107
rect 7192 30104 7204 30107
rect 9125 30107 9183 30113
rect 9125 30104 9137 30107
rect 7192 30076 9137 30104
rect 7192 30073 7204 30076
rect 7156 30067 7204 30073
rect 9125 30073 9137 30076
rect 9171 30104 9183 30107
rect 9493 30107 9551 30113
rect 9493 30104 9505 30107
rect 9171 30076 9505 30104
rect 9171 30073 9183 30076
rect 9125 30067 9183 30073
rect 9493 30073 9505 30076
rect 9539 30104 9551 30107
rect 9998 30107 10056 30113
rect 9998 30104 10010 30107
rect 9539 30076 10010 30104
rect 9539 30073 9551 30076
rect 9493 30067 9551 30073
rect 9998 30073 10010 30076
rect 10044 30073 10056 30107
rect 9998 30067 10056 30073
rect 7156 30064 7162 30067
rect 8386 30036 8392 30048
rect 8347 30008 8392 30036
rect 8386 29996 8392 30008
rect 8444 29996 8450 30048
rect 9674 29996 9680 30048
rect 9732 30036 9738 30048
rect 10873 30039 10931 30045
rect 10873 30036 10885 30039
rect 9732 30008 10885 30036
rect 9732 29996 9738 30008
rect 10873 30005 10885 30008
rect 10919 30005 10931 30039
rect 10873 29999 10931 30005
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 4617 29835 4675 29841
rect 4617 29801 4629 29835
rect 4663 29832 4675 29835
rect 5074 29832 5080 29844
rect 4663 29804 5080 29832
rect 4663 29801 4675 29804
rect 4617 29795 4675 29801
rect 5074 29792 5080 29804
rect 5132 29832 5138 29844
rect 5350 29832 5356 29844
rect 5132 29804 5356 29832
rect 5132 29792 5138 29804
rect 5350 29792 5356 29804
rect 5408 29792 5414 29844
rect 7561 29835 7619 29841
rect 7561 29801 7573 29835
rect 7607 29832 7619 29835
rect 7834 29832 7840 29844
rect 7607 29804 7840 29832
rect 7607 29801 7619 29804
rect 7561 29795 7619 29801
rect 7834 29792 7840 29804
rect 7892 29792 7898 29844
rect 8018 29792 8024 29844
rect 8076 29832 8082 29844
rect 8389 29835 8447 29841
rect 8389 29832 8401 29835
rect 8076 29804 8401 29832
rect 8076 29792 8082 29804
rect 8389 29801 8401 29804
rect 8435 29801 8447 29835
rect 8389 29795 8447 29801
rect 9493 29835 9551 29841
rect 9493 29801 9505 29835
rect 9539 29832 9551 29835
rect 9582 29832 9588 29844
rect 9539 29804 9588 29832
rect 9539 29801 9551 29804
rect 9493 29795 9551 29801
rect 9582 29792 9588 29804
rect 9640 29792 9646 29844
rect 11241 29835 11299 29841
rect 11241 29801 11253 29835
rect 11287 29832 11299 29835
rect 11514 29832 11520 29844
rect 11287 29804 11520 29832
rect 11287 29801 11299 29804
rect 11241 29795 11299 29801
rect 11514 29792 11520 29804
rect 11572 29792 11578 29844
rect 12391 29835 12449 29841
rect 12391 29801 12403 29835
rect 12437 29801 12449 29835
rect 12391 29795 12449 29801
rect 4798 29724 4804 29776
rect 4856 29764 4862 29776
rect 4893 29767 4951 29773
rect 4893 29764 4905 29767
rect 4856 29736 4905 29764
rect 4856 29724 4862 29736
rect 4893 29733 4905 29736
rect 4939 29733 4951 29767
rect 4893 29727 4951 29733
rect 6546 29724 6552 29776
rect 6604 29764 6610 29776
rect 6962 29767 7020 29773
rect 6962 29764 6974 29767
rect 6604 29736 6974 29764
rect 6604 29724 6610 29736
rect 6962 29733 6974 29736
rect 7008 29764 7020 29767
rect 7098 29764 7104 29776
rect 7008 29736 7104 29764
rect 7008 29733 7020 29736
rect 6962 29727 7020 29733
rect 7098 29724 7104 29736
rect 7156 29724 7162 29776
rect 9861 29767 9919 29773
rect 9861 29733 9873 29767
rect 9907 29764 9919 29767
rect 10042 29764 10048 29776
rect 9907 29736 10048 29764
rect 9907 29733 9919 29736
rect 9861 29727 9919 29733
rect 10042 29724 10048 29736
rect 10100 29724 10106 29776
rect 10686 29724 10692 29776
rect 10744 29764 10750 29776
rect 12406 29764 12434 29795
rect 10744 29736 12434 29764
rect 10744 29724 10750 29736
rect 3050 29705 3056 29708
rect 3028 29699 3056 29705
rect 3028 29665 3040 29699
rect 3028 29659 3056 29665
rect 3050 29656 3056 29659
rect 3108 29656 3114 29708
rect 12342 29705 12348 29708
rect 12320 29699 12348 29705
rect 12320 29665 12332 29699
rect 12320 29659 12348 29665
rect 12342 29656 12348 29659
rect 12400 29656 12406 29708
rect 4798 29628 4804 29640
rect 4759 29600 4804 29628
rect 4798 29588 4804 29600
rect 4856 29588 4862 29640
rect 6178 29588 6184 29640
rect 6236 29628 6242 29640
rect 6641 29631 6699 29637
rect 6641 29628 6653 29631
rect 6236 29600 6653 29628
rect 6236 29588 6242 29600
rect 6641 29597 6653 29600
rect 6687 29628 6699 29631
rect 7374 29628 7380 29640
rect 6687 29600 7380 29628
rect 6687 29597 6699 29600
rect 6641 29591 6699 29597
rect 7374 29588 7380 29600
rect 7432 29588 7438 29640
rect 9769 29631 9827 29637
rect 9769 29597 9781 29631
rect 9815 29628 9827 29631
rect 9950 29628 9956 29640
rect 9815 29600 9956 29628
rect 9815 29597 9827 29600
rect 9769 29591 9827 29597
rect 9950 29588 9956 29600
rect 10008 29588 10014 29640
rect 10413 29631 10471 29637
rect 10413 29597 10425 29631
rect 10459 29628 10471 29631
rect 10778 29628 10784 29640
rect 10459 29600 10784 29628
rect 10459 29597 10471 29600
rect 10413 29591 10471 29597
rect 10778 29588 10784 29600
rect 10836 29588 10842 29640
rect 5350 29560 5356 29572
rect 4448 29532 4660 29560
rect 5311 29532 5356 29560
rect 4448 29504 4476 29532
rect 3099 29495 3157 29501
rect 3099 29461 3111 29495
rect 3145 29492 3157 29495
rect 4430 29492 4436 29504
rect 3145 29464 4436 29492
rect 3145 29461 3157 29464
rect 3099 29455 3157 29461
rect 4430 29452 4436 29464
rect 4488 29452 4494 29504
rect 4632 29492 4660 29532
rect 5350 29520 5356 29532
rect 5408 29520 5414 29572
rect 5721 29495 5779 29501
rect 5721 29492 5733 29495
rect 4632 29464 5733 29492
rect 5721 29461 5733 29464
rect 5767 29461 5779 29495
rect 6362 29492 6368 29504
rect 6323 29464 6368 29492
rect 5721 29455 5779 29461
rect 6362 29452 6368 29464
rect 6420 29452 6426 29504
rect 10781 29495 10839 29501
rect 10781 29461 10793 29495
rect 10827 29492 10839 29495
rect 10962 29492 10968 29504
rect 10827 29464 10968 29492
rect 10827 29461 10839 29464
rect 10781 29455 10839 29461
rect 10962 29452 10968 29464
rect 11020 29452 11026 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 11054 29248 11060 29300
rect 11112 29288 11118 29300
rect 12342 29288 12348 29300
rect 11112 29260 12348 29288
rect 11112 29248 11118 29260
rect 12342 29248 12348 29260
rect 12400 29288 12406 29300
rect 12986 29288 12992 29300
rect 12400 29260 12992 29288
rect 12400 29248 12406 29260
rect 12986 29248 12992 29260
rect 13044 29248 13050 29300
rect 5166 29180 5172 29232
rect 5224 29220 5230 29232
rect 6546 29220 6552 29232
rect 5224 29192 6552 29220
rect 5224 29180 5230 29192
rect 6546 29180 6552 29192
rect 6604 29220 6610 29232
rect 10962 29220 10968 29232
rect 6604 29192 8708 29220
rect 6604 29180 6610 29192
rect 4430 29112 4436 29164
rect 4488 29152 4494 29164
rect 4985 29155 5043 29161
rect 4985 29152 4997 29155
rect 4488 29124 4997 29152
rect 4488 29112 4494 29124
rect 4985 29121 4997 29124
rect 5031 29121 5043 29155
rect 5350 29152 5356 29164
rect 5311 29124 5356 29152
rect 4985 29115 5043 29121
rect 5350 29112 5356 29124
rect 5408 29112 5414 29164
rect 7374 29152 7380 29164
rect 7335 29124 7380 29152
rect 7374 29112 7380 29124
rect 7432 29112 7438 29164
rect 3510 29044 3516 29096
rect 3568 29084 3574 29096
rect 3932 29087 3990 29093
rect 3932 29084 3944 29087
rect 3568 29056 3944 29084
rect 3568 29044 3574 29056
rect 3932 29053 3944 29056
rect 3978 29084 3990 29087
rect 4246 29084 4252 29096
rect 3978 29056 4252 29084
rect 3978 29053 3990 29056
rect 3932 29047 3990 29053
rect 4246 29044 4252 29056
rect 4304 29084 4310 29096
rect 4341 29087 4399 29093
rect 4341 29084 4353 29087
rect 4304 29056 4353 29084
rect 4304 29044 4310 29056
rect 4341 29053 4353 29056
rect 4387 29053 4399 29087
rect 4341 29047 4399 29053
rect 6273 29087 6331 29093
rect 6273 29053 6285 29087
rect 6319 29084 6331 29087
rect 7006 29084 7012 29096
rect 6319 29056 7012 29084
rect 6319 29053 6331 29056
rect 6273 29047 6331 29053
rect 7006 29044 7012 29056
rect 7064 29044 7070 29096
rect 7282 29084 7288 29096
rect 7243 29056 7288 29084
rect 7282 29044 7288 29056
rect 7340 29044 7346 29096
rect 8573 29087 8631 29093
rect 8573 29053 8585 29087
rect 8619 29053 8631 29087
rect 8573 29047 8631 29053
rect 3050 29016 3056 29028
rect 3011 28988 3056 29016
rect 3050 28976 3056 28988
rect 3108 28976 3114 29028
rect 4019 29019 4077 29025
rect 4019 28985 4031 29019
rect 4065 29016 4077 29019
rect 4798 29016 4804 29028
rect 4065 28988 4804 29016
rect 4065 28985 4077 28988
rect 4019 28979 4077 28985
rect 4798 28976 4804 28988
rect 4856 28976 4862 29028
rect 5077 29019 5135 29025
rect 5077 29016 5089 29019
rect 4908 28988 5089 29016
rect 4908 28960 4936 28988
rect 5077 28985 5089 28988
rect 5123 28985 5135 29019
rect 6362 29016 6368 29028
rect 5077 28979 5135 28985
rect 5368 28988 6368 29016
rect 4706 28948 4712 28960
rect 4667 28920 4712 28948
rect 4706 28908 4712 28920
rect 4764 28908 4770 28960
rect 4890 28908 4896 28960
rect 4948 28908 4954 28960
rect 5368 28948 5396 28988
rect 6362 28976 6368 28988
rect 6420 28976 6426 29028
rect 8113 29019 8171 29025
rect 8113 28985 8125 29019
rect 8159 29016 8171 29019
rect 8294 29016 8300 29028
rect 8159 28988 8300 29016
rect 8159 28985 8171 28988
rect 8113 28979 8171 28985
rect 8294 28976 8300 28988
rect 8352 29016 8358 29028
rect 8588 29016 8616 29047
rect 8680 29016 8708 29192
rect 10428 29192 10968 29220
rect 10428 29161 10456 29192
rect 10962 29180 10968 29192
rect 11020 29180 11026 29232
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29121 10471 29155
rect 10870 29152 10876 29164
rect 10831 29124 10876 29152
rect 10413 29115 10471 29121
rect 10870 29112 10876 29124
rect 10928 29112 10934 29164
rect 9493 29087 9551 29093
rect 9493 29053 9505 29087
rect 9539 29084 9551 29087
rect 9539 29056 10272 29084
rect 9539 29053 9551 29056
rect 9493 29047 9551 29053
rect 8894 29019 8952 29025
rect 8894 29016 8906 29019
rect 8352 28988 8616 29016
rect 8655 28988 8906 29016
rect 8352 28976 8358 28988
rect 5534 28948 5540 28960
rect 5368 28920 5540 28948
rect 5534 28908 5540 28920
rect 5592 28908 5598 28960
rect 8386 28948 8392 28960
rect 8347 28920 8392 28948
rect 8386 28908 8392 28920
rect 8444 28948 8450 28960
rect 8655 28948 8683 28988
rect 8894 28985 8906 28988
rect 8940 28985 8952 29019
rect 8894 28979 8952 28985
rect 9861 29019 9919 29025
rect 9861 28985 9873 29019
rect 9907 29016 9919 29019
rect 10042 29016 10048 29028
rect 9907 28988 10048 29016
rect 9907 28985 9919 28988
rect 9861 28979 9919 28985
rect 10042 28976 10048 28988
rect 10100 28976 10106 29028
rect 10244 29025 10272 29056
rect 12434 29044 12440 29096
rect 12492 29084 12498 29096
rect 13265 29087 13323 29093
rect 13265 29084 13277 29087
rect 12492 29056 13277 29084
rect 12492 29044 12498 29056
rect 13265 29053 13277 29056
rect 13311 29053 13323 29087
rect 13265 29047 13323 29053
rect 13446 29044 13452 29096
rect 13504 29093 13510 29096
rect 13504 29087 13542 29093
rect 13530 29084 13542 29087
rect 13909 29087 13967 29093
rect 13909 29084 13921 29087
rect 13530 29056 13921 29084
rect 13530 29053 13542 29056
rect 13504 29047 13542 29053
rect 13909 29053 13921 29056
rect 13955 29053 13967 29087
rect 13909 29047 13967 29053
rect 13504 29044 13510 29047
rect 10229 29019 10287 29025
rect 10229 28985 10241 29019
rect 10275 29016 10287 29019
rect 10505 29019 10563 29025
rect 10505 29016 10517 29019
rect 10275 28988 10517 29016
rect 10275 28985 10287 28988
rect 10229 28979 10287 28985
rect 10505 28985 10517 28988
rect 10551 29016 10563 29019
rect 11054 29016 11060 29028
rect 10551 28988 11060 29016
rect 10551 28985 10563 28988
rect 10505 28979 10563 28985
rect 11054 28976 11060 28988
rect 11112 28976 11118 29028
rect 12986 28976 12992 29028
rect 13044 29016 13050 29028
rect 13587 29019 13645 29025
rect 13587 29016 13599 29019
rect 13044 28988 13599 29016
rect 13044 28976 13050 28988
rect 13587 28985 13599 28988
rect 13633 28985 13645 29019
rect 13587 28979 13645 28985
rect 8444 28920 8683 28948
rect 8444 28908 8450 28920
rect 9766 28908 9772 28960
rect 9824 28948 9830 28960
rect 12621 28951 12679 28957
rect 12621 28948 12633 28951
rect 9824 28920 12633 28948
rect 9824 28908 9830 28920
rect 12621 28917 12633 28920
rect 12667 28917 12679 28951
rect 12621 28911 12679 28917
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 4617 28747 4675 28753
rect 4617 28713 4629 28747
rect 4663 28744 4675 28747
rect 4798 28744 4804 28756
rect 4663 28716 4804 28744
rect 4663 28713 4675 28716
rect 4617 28707 4675 28713
rect 4798 28704 4804 28716
rect 4856 28704 4862 28756
rect 5718 28704 5724 28756
rect 5776 28704 5782 28756
rect 6178 28744 6184 28756
rect 6139 28716 6184 28744
rect 6178 28704 6184 28716
rect 6236 28704 6242 28756
rect 9950 28744 9956 28756
rect 9911 28716 9956 28744
rect 9950 28704 9956 28716
rect 10008 28704 10014 28756
rect 11238 28704 11244 28756
rect 11296 28744 11302 28756
rect 11296 28716 12480 28744
rect 11296 28704 11302 28716
rect 4706 28676 4712 28688
rect 4667 28648 4712 28676
rect 4706 28636 4712 28648
rect 4764 28636 4770 28688
rect 5736 28676 5764 28704
rect 7282 28676 7288 28688
rect 5736 28648 7288 28676
rect 6748 28620 6776 28648
rect 7282 28636 7288 28648
rect 7340 28636 7346 28688
rect 8757 28679 8815 28685
rect 8757 28645 8769 28679
rect 8803 28676 8815 28679
rect 9582 28676 9588 28688
rect 8803 28648 9588 28676
rect 8803 28645 8815 28648
rect 8757 28639 8815 28645
rect 9582 28636 9588 28648
rect 9640 28636 9646 28688
rect 10321 28679 10379 28685
rect 10321 28645 10333 28679
rect 10367 28676 10379 28679
rect 11146 28676 11152 28688
rect 10367 28648 11152 28676
rect 10367 28645 10379 28648
rect 10321 28639 10379 28645
rect 11146 28636 11152 28648
rect 11204 28676 11210 28688
rect 11885 28679 11943 28685
rect 11885 28676 11897 28679
rect 11204 28648 11897 28676
rect 11204 28636 11210 28648
rect 11885 28645 11897 28648
rect 11931 28645 11943 28679
rect 11885 28639 11943 28645
rect 4798 28608 4804 28620
rect 4759 28580 4804 28608
rect 4798 28568 4804 28580
rect 4856 28608 4862 28620
rect 5721 28611 5779 28617
rect 5721 28608 5733 28611
rect 4856 28580 5733 28608
rect 4856 28568 4862 28580
rect 5721 28577 5733 28580
rect 5767 28577 5779 28611
rect 6546 28608 6552 28620
rect 6507 28580 6552 28608
rect 5721 28571 5779 28577
rect 6546 28568 6552 28580
rect 6604 28568 6610 28620
rect 6730 28608 6736 28620
rect 6643 28580 6736 28608
rect 6730 28568 6736 28580
rect 6788 28568 6794 28620
rect 8018 28608 8024 28620
rect 7979 28580 8024 28608
rect 8018 28568 8024 28580
rect 8076 28568 8082 28620
rect 8573 28611 8631 28617
rect 8573 28577 8585 28611
rect 8619 28608 8631 28611
rect 9766 28608 9772 28620
rect 8619 28580 9772 28608
rect 8619 28577 8631 28580
rect 8573 28571 8631 28577
rect 9766 28568 9772 28580
rect 9824 28568 9830 28620
rect 10870 28568 10876 28620
rect 10928 28608 10934 28620
rect 12452 28608 12480 28716
rect 13300 28611 13358 28617
rect 13300 28608 13312 28611
rect 10928 28580 10973 28608
rect 12452 28580 13312 28608
rect 10928 28568 10934 28580
rect 13300 28577 13312 28580
rect 13346 28608 13358 28611
rect 13630 28608 13636 28620
rect 13346 28580 13636 28608
rect 13346 28577 13358 28580
rect 13300 28571 13358 28577
rect 13630 28568 13636 28580
rect 13688 28568 13694 28620
rect 6822 28540 6828 28552
rect 6783 28512 6828 28540
rect 6822 28500 6828 28512
rect 6880 28500 6886 28552
rect 10226 28540 10232 28552
rect 10187 28512 10232 28540
rect 10226 28500 10232 28512
rect 10284 28500 10290 28552
rect 11793 28543 11851 28549
rect 11793 28509 11805 28543
rect 11839 28540 11851 28543
rect 12526 28540 12532 28552
rect 11839 28512 12532 28540
rect 11839 28509 11851 28512
rect 11793 28503 11851 28509
rect 12526 28500 12532 28512
rect 12584 28540 12590 28552
rect 12584 28512 12848 28540
rect 12584 28500 12590 28512
rect 10778 28432 10784 28484
rect 10836 28472 10842 28484
rect 12342 28472 12348 28484
rect 10836 28444 12348 28472
rect 10836 28432 10842 28444
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 12820 28472 12848 28512
rect 13403 28475 13461 28481
rect 13403 28472 13415 28475
rect 12820 28444 13415 28472
rect 13403 28441 13415 28444
rect 13449 28441 13461 28475
rect 13403 28435 13461 28441
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 4525 28203 4583 28209
rect 4525 28169 4537 28203
rect 4571 28200 4583 28203
rect 4798 28200 4804 28212
rect 4571 28172 4804 28200
rect 4571 28169 4583 28172
rect 4525 28163 4583 28169
rect 4798 28160 4804 28172
rect 4856 28200 4862 28212
rect 5905 28203 5963 28209
rect 5905 28200 5917 28203
rect 4856 28172 5917 28200
rect 4856 28160 4862 28172
rect 5905 28169 5917 28172
rect 5951 28169 5963 28203
rect 9766 28200 9772 28212
rect 9727 28172 9772 28200
rect 5905 28163 5963 28169
rect 9766 28160 9772 28172
rect 9824 28160 9830 28212
rect 11146 28200 11152 28212
rect 11107 28172 11152 28200
rect 11146 28160 11152 28172
rect 11204 28200 11210 28212
rect 11425 28203 11483 28209
rect 11425 28200 11437 28203
rect 11204 28172 11437 28200
rect 11204 28160 11210 28172
rect 11425 28169 11437 28172
rect 11471 28200 11483 28203
rect 11793 28203 11851 28209
rect 11793 28200 11805 28203
rect 11471 28172 11805 28200
rect 11471 28169 11483 28172
rect 11425 28163 11483 28169
rect 11793 28169 11805 28172
rect 11839 28169 11851 28203
rect 13630 28200 13636 28212
rect 13591 28172 13636 28200
rect 11793 28163 11851 28169
rect 13630 28160 13636 28172
rect 13688 28160 13694 28212
rect 8662 28132 8668 28144
rect 4724 28104 8668 28132
rect 3329 28067 3387 28073
rect 3329 28033 3341 28067
rect 3375 28064 3387 28067
rect 3375 28036 4200 28064
rect 3375 28033 3387 28036
rect 3329 28027 3387 28033
rect 3697 27999 3755 28005
rect 3697 27965 3709 27999
rect 3743 27965 3755 27999
rect 3697 27959 3755 27965
rect 3789 27999 3847 28005
rect 3789 27965 3801 27999
rect 3835 27996 3847 27999
rect 3878 27996 3884 28008
rect 3835 27968 3884 27996
rect 3835 27965 3847 27968
rect 3789 27959 3847 27965
rect 3510 27820 3516 27872
rect 3568 27860 3574 27872
rect 3712 27860 3740 27959
rect 3878 27956 3884 27968
rect 3936 27956 3942 28008
rect 4172 28005 4200 28036
rect 4157 27999 4215 28005
rect 4157 27965 4169 27999
rect 4203 27996 4215 27999
rect 4724 27996 4752 28104
rect 8662 28092 8668 28104
rect 8720 28092 8726 28144
rect 10962 28092 10968 28144
rect 11020 28132 11026 28144
rect 13170 28132 13176 28144
rect 11020 28104 13176 28132
rect 11020 28092 11026 28104
rect 13170 28092 13176 28104
rect 13228 28092 13234 28144
rect 4890 28064 4896 28076
rect 4803 28036 4896 28064
rect 4890 28024 4896 28036
rect 4948 28064 4954 28076
rect 5166 28064 5172 28076
rect 4948 28036 5172 28064
rect 4948 28024 4954 28036
rect 5166 28024 5172 28036
rect 5224 28024 5230 28076
rect 6546 28024 6552 28076
rect 6604 28064 6610 28076
rect 6822 28064 6828 28076
rect 6604 28036 6828 28064
rect 6604 28024 6610 28036
rect 6822 28024 6828 28036
rect 6880 28064 6886 28076
rect 7929 28067 7987 28073
rect 7929 28064 7941 28067
rect 6880 28036 7941 28064
rect 6880 28024 6886 28036
rect 7929 28033 7941 28036
rect 7975 28064 7987 28067
rect 8018 28064 8024 28076
rect 7975 28036 8024 28064
rect 7975 28033 7987 28036
rect 7929 28027 7987 28033
rect 8018 28024 8024 28036
rect 8076 28024 8082 28076
rect 11974 28024 11980 28076
rect 12032 28064 12038 28076
rect 13265 28067 13323 28073
rect 13265 28064 13277 28067
rect 12032 28036 13277 28064
rect 12032 28024 12038 28036
rect 4982 27996 4988 28008
rect 4203 27968 4752 27996
rect 4943 27968 4988 27996
rect 4203 27965 4215 27968
rect 4157 27959 4215 27965
rect 4982 27956 4988 27968
rect 5040 27956 5046 28008
rect 5184 27928 5212 28024
rect 7193 27999 7251 28005
rect 7193 27965 7205 27999
rect 7239 27965 7251 27999
rect 7193 27959 7251 27965
rect 5306 27931 5364 27937
rect 5306 27928 5318 27931
rect 5184 27900 5318 27928
rect 5306 27897 5318 27900
rect 5352 27897 5364 27931
rect 5306 27891 5364 27897
rect 6641 27931 6699 27937
rect 6641 27897 6653 27931
rect 6687 27928 6699 27931
rect 7208 27928 7236 27959
rect 7282 27956 7288 28008
rect 7340 27996 7346 28008
rect 7377 27999 7435 28005
rect 7377 27996 7389 27999
rect 7340 27968 7389 27996
rect 7340 27956 7346 27968
rect 7377 27965 7389 27968
rect 7423 27965 7435 27999
rect 7377 27959 7435 27965
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27996 7711 27999
rect 8481 27999 8539 28005
rect 8481 27996 8493 27999
rect 7699 27968 8493 27996
rect 7699 27965 7711 27968
rect 7653 27959 7711 27965
rect 8481 27965 8493 27968
rect 8527 27996 8539 27999
rect 8938 27996 8944 28008
rect 8527 27968 8944 27996
rect 8527 27965 8539 27968
rect 8481 27959 8539 27965
rect 8938 27956 8944 27968
rect 8996 27956 9002 28008
rect 9674 27956 9680 28008
rect 9732 27996 9738 28008
rect 12636 28005 12664 28036
rect 13265 28033 13277 28036
rect 13311 28033 13323 28067
rect 13265 28027 13323 28033
rect 10229 27999 10287 28005
rect 10229 27996 10241 27999
rect 9732 27968 10241 27996
rect 9732 27956 9738 27968
rect 10229 27965 10241 27968
rect 10275 27965 10287 27999
rect 12437 27999 12495 28005
rect 12437 27996 12449 27999
rect 10229 27959 10287 27965
rect 12176 27968 12449 27996
rect 7466 27928 7472 27940
rect 6687 27900 7472 27928
rect 6687 27897 6699 27900
rect 6641 27891 6699 27897
rect 7466 27888 7472 27900
rect 7524 27928 7530 27940
rect 8386 27928 8392 27940
rect 7524 27900 7696 27928
rect 8299 27900 8392 27928
rect 7524 27888 7530 27900
rect 7668 27872 7696 27900
rect 8386 27888 8392 27900
rect 8444 27928 8450 27940
rect 8843 27931 8901 27937
rect 8843 27928 8855 27931
rect 8444 27900 8855 27928
rect 8444 27888 8450 27900
rect 8843 27897 8855 27900
rect 8889 27928 8901 27931
rect 9766 27928 9772 27940
rect 8889 27900 9772 27928
rect 8889 27897 8901 27900
rect 8843 27891 8901 27897
rect 9766 27888 9772 27900
rect 9824 27928 9830 27940
rect 10045 27931 10103 27937
rect 10045 27928 10057 27931
rect 9824 27900 10057 27928
rect 9824 27888 9830 27900
rect 10045 27897 10057 27900
rect 10091 27928 10103 27931
rect 10550 27931 10608 27937
rect 10550 27928 10562 27931
rect 10091 27900 10562 27928
rect 10091 27897 10103 27900
rect 10045 27891 10103 27897
rect 10550 27897 10562 27900
rect 10596 27897 10608 27931
rect 10550 27891 10608 27897
rect 5534 27860 5540 27872
rect 3568 27832 5540 27860
rect 3568 27820 3574 27832
rect 5534 27820 5540 27832
rect 5592 27820 5598 27872
rect 6273 27863 6331 27869
rect 6273 27829 6285 27863
rect 6319 27860 6331 27863
rect 6822 27860 6828 27872
rect 6319 27832 6828 27860
rect 6319 27829 6331 27832
rect 6273 27823 6331 27829
rect 6822 27820 6828 27832
rect 6880 27820 6886 27872
rect 7650 27820 7656 27872
rect 7708 27820 7714 27872
rect 9398 27860 9404 27872
rect 9359 27832 9404 27860
rect 9398 27820 9404 27832
rect 9456 27820 9462 27872
rect 10134 27820 10140 27872
rect 10192 27860 10198 27872
rect 10318 27860 10324 27872
rect 10192 27832 10324 27860
rect 10192 27820 10198 27832
rect 10318 27820 10324 27832
rect 10376 27820 10382 27872
rect 11422 27820 11428 27872
rect 11480 27860 11486 27872
rect 12176 27869 12204 27968
rect 12437 27965 12449 27968
rect 12483 27965 12495 27999
rect 12437 27959 12495 27965
rect 12621 27999 12679 28005
rect 12621 27965 12633 27999
rect 12667 27965 12679 27999
rect 12621 27959 12679 27965
rect 12161 27863 12219 27869
rect 12161 27860 12173 27863
rect 11480 27832 12173 27860
rect 11480 27820 11486 27832
rect 12161 27829 12173 27832
rect 12207 27829 12219 27863
rect 12710 27860 12716 27872
rect 12671 27832 12716 27860
rect 12161 27823 12219 27829
rect 12710 27820 12716 27832
rect 12768 27820 12774 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 3510 27656 3516 27668
rect 3471 27628 3516 27656
rect 3510 27616 3516 27628
rect 3568 27616 3574 27668
rect 4709 27659 4767 27665
rect 4709 27625 4721 27659
rect 4755 27656 4767 27659
rect 4982 27656 4988 27668
rect 4755 27628 4988 27656
rect 4755 27625 4767 27628
rect 4709 27619 4767 27625
rect 4982 27616 4988 27628
rect 5040 27656 5046 27668
rect 5261 27659 5319 27665
rect 5261 27656 5273 27659
rect 5040 27628 5273 27656
rect 5040 27616 5046 27628
rect 5261 27625 5273 27628
rect 5307 27625 5319 27659
rect 5261 27619 5319 27625
rect 6641 27659 6699 27665
rect 6641 27625 6653 27659
rect 6687 27656 6699 27659
rect 6730 27656 6736 27668
rect 6687 27628 6736 27656
rect 6687 27625 6699 27628
rect 6641 27619 6699 27625
rect 6730 27616 6736 27628
rect 6788 27616 6794 27668
rect 8938 27656 8944 27668
rect 8899 27628 8944 27656
rect 8938 27616 8944 27628
rect 8996 27616 9002 27668
rect 9398 27616 9404 27668
rect 9456 27656 9462 27668
rect 9456 27628 9628 27656
rect 9456 27616 9462 27628
rect 5442 27588 5448 27600
rect 4172 27560 5448 27588
rect 4172 27532 4200 27560
rect 5442 27548 5448 27560
rect 5500 27548 5506 27600
rect 7009 27591 7067 27597
rect 7009 27557 7021 27591
rect 7055 27588 7067 27591
rect 7282 27588 7288 27600
rect 7055 27560 7288 27588
rect 7055 27557 7067 27560
rect 7009 27551 7067 27557
rect 7282 27548 7288 27560
rect 7340 27588 7346 27600
rect 9600 27588 9628 27628
rect 9674 27616 9680 27668
rect 9732 27656 9738 27668
rect 10965 27659 11023 27665
rect 10965 27656 10977 27659
rect 9732 27628 10977 27656
rect 9732 27616 9738 27628
rect 10965 27625 10977 27628
rect 11011 27625 11023 27659
rect 12526 27656 12532 27668
rect 12487 27628 12532 27656
rect 10965 27619 11023 27625
rect 12526 27616 12532 27628
rect 12584 27616 12590 27668
rect 13170 27616 13176 27668
rect 13228 27665 13234 27668
rect 13228 27659 13277 27665
rect 13228 27625 13231 27659
rect 13265 27625 13277 27659
rect 13228 27619 13277 27625
rect 13228 27616 13234 27619
rect 10042 27588 10048 27600
rect 7340 27560 8432 27588
rect 9600 27560 10048 27588
rect 7340 27548 7346 27560
rect 8404 27532 8432 27560
rect 10042 27548 10048 27560
rect 10100 27588 10106 27600
rect 10137 27591 10195 27597
rect 10137 27588 10149 27591
rect 10100 27560 10149 27588
rect 10100 27548 10106 27560
rect 10137 27557 10149 27560
rect 10183 27557 10195 27591
rect 10137 27551 10195 27557
rect 10689 27591 10747 27597
rect 10689 27557 10701 27591
rect 10735 27588 10747 27591
rect 10870 27588 10876 27600
rect 10735 27560 10876 27588
rect 10735 27557 10747 27560
rect 10689 27551 10747 27557
rect 10870 27548 10876 27560
rect 10928 27588 10934 27600
rect 11333 27591 11391 27597
rect 11333 27588 11345 27591
rect 10928 27560 11345 27588
rect 10928 27548 10934 27560
rect 11333 27557 11345 27560
rect 11379 27557 11391 27591
rect 11606 27588 11612 27600
rect 11333 27551 11391 27557
rect 11440 27560 11612 27588
rect 4154 27520 4160 27532
rect 4067 27492 4160 27520
rect 4154 27480 4160 27492
rect 4212 27480 4218 27532
rect 4890 27480 4896 27532
rect 4948 27520 4954 27532
rect 4985 27523 5043 27529
rect 4985 27520 4997 27523
rect 4948 27492 4997 27520
rect 4948 27480 4954 27492
rect 4985 27489 4997 27492
rect 5031 27489 5043 27523
rect 5166 27520 5172 27532
rect 5127 27492 5172 27520
rect 4985 27483 5043 27489
rect 5166 27480 5172 27492
rect 5224 27480 5230 27532
rect 5629 27523 5687 27529
rect 5629 27520 5641 27523
rect 5552 27492 5641 27520
rect 5552 27452 5580 27492
rect 5629 27489 5641 27492
rect 5675 27489 5687 27523
rect 5994 27520 6000 27532
rect 5955 27492 6000 27520
rect 5629 27483 5687 27489
rect 5994 27480 6000 27492
rect 6052 27480 6058 27532
rect 7374 27480 7380 27532
rect 7432 27520 7438 27532
rect 7558 27520 7564 27532
rect 7432 27492 7564 27520
rect 7432 27480 7438 27492
rect 7558 27480 7564 27492
rect 7616 27520 7622 27532
rect 7929 27523 7987 27529
rect 7929 27520 7941 27523
rect 7616 27492 7941 27520
rect 7616 27480 7622 27492
rect 7929 27489 7941 27492
rect 7975 27489 7987 27523
rect 8386 27520 8392 27532
rect 8347 27492 8392 27520
rect 7929 27483 7987 27489
rect 8386 27480 8392 27492
rect 8444 27480 8450 27532
rect 11054 27480 11060 27532
rect 11112 27520 11118 27532
rect 11440 27520 11468 27560
rect 11606 27548 11612 27560
rect 11664 27588 11670 27600
rect 11701 27591 11759 27597
rect 11701 27588 11713 27591
rect 11664 27560 11713 27588
rect 11664 27548 11670 27560
rect 11701 27557 11713 27560
rect 11747 27557 11759 27591
rect 11701 27551 11759 27557
rect 12253 27591 12311 27597
rect 12253 27557 12265 27591
rect 12299 27588 12311 27591
rect 12342 27588 12348 27600
rect 12299 27560 12348 27588
rect 12299 27557 12311 27560
rect 12253 27551 12311 27557
rect 12342 27548 12348 27560
rect 12400 27548 12406 27600
rect 11112 27492 11468 27520
rect 11112 27480 11118 27492
rect 13078 27480 13084 27532
rect 13136 27529 13142 27532
rect 13136 27523 13174 27529
rect 13162 27489 13174 27523
rect 13136 27483 13174 27489
rect 13136 27480 13142 27483
rect 6178 27452 6184 27464
rect 5552 27424 6184 27452
rect 4341 27387 4399 27393
rect 4341 27353 4353 27387
rect 4387 27384 4399 27387
rect 5552 27384 5580 27424
rect 6178 27412 6184 27424
rect 6236 27412 6242 27464
rect 8294 27412 8300 27464
rect 8352 27452 8358 27464
rect 8481 27455 8539 27461
rect 8481 27452 8493 27455
rect 8352 27424 8493 27452
rect 8352 27412 8358 27424
rect 8481 27421 8493 27424
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 10045 27455 10103 27461
rect 10045 27421 10057 27455
rect 10091 27452 10103 27455
rect 10134 27452 10140 27464
rect 10091 27424 10140 27452
rect 10091 27421 10103 27424
rect 10045 27415 10103 27421
rect 10134 27412 10140 27424
rect 10192 27452 10198 27464
rect 10686 27452 10692 27464
rect 10192 27424 10692 27452
rect 10192 27412 10198 27424
rect 10686 27412 10692 27424
rect 10744 27412 10750 27464
rect 11609 27455 11667 27461
rect 11609 27421 11621 27455
rect 11655 27421 11667 27455
rect 11609 27415 11667 27421
rect 4387 27356 5580 27384
rect 4387 27353 4399 27356
rect 4341 27347 4399 27353
rect 11514 27344 11520 27396
rect 11572 27384 11578 27396
rect 11624 27384 11652 27415
rect 11572 27356 11652 27384
rect 11572 27344 11578 27356
rect 9490 27316 9496 27328
rect 9451 27288 9496 27316
rect 9490 27276 9496 27288
rect 9548 27276 9554 27328
rect 11330 27276 11336 27328
rect 11388 27316 11394 27328
rect 12158 27316 12164 27328
rect 11388 27288 12164 27316
rect 11388 27276 11394 27288
rect 12158 27276 12164 27288
rect 12216 27276 12222 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 4154 27112 4160 27124
rect 4115 27084 4160 27112
rect 4154 27072 4160 27084
rect 4212 27072 4218 27124
rect 5902 27112 5908 27124
rect 5863 27084 5908 27112
rect 5902 27072 5908 27084
rect 5960 27072 5966 27124
rect 6178 27112 6184 27124
rect 6139 27084 6184 27112
rect 6178 27072 6184 27084
rect 6236 27072 6242 27124
rect 6730 27072 6736 27124
rect 6788 27112 6794 27124
rect 7009 27115 7067 27121
rect 7009 27112 7021 27115
rect 6788 27084 7021 27112
rect 6788 27072 6794 27084
rect 7009 27081 7021 27084
rect 7055 27081 7067 27115
rect 10042 27112 10048 27124
rect 10003 27084 10048 27112
rect 7009 27075 7067 27081
rect 10042 27072 10048 27084
rect 10100 27072 10106 27124
rect 11606 27112 11612 27124
rect 11567 27084 11612 27112
rect 11606 27072 11612 27084
rect 11664 27072 11670 27124
rect 12434 27072 12440 27124
rect 12492 27112 12498 27124
rect 12575 27115 12633 27121
rect 12575 27112 12587 27115
rect 12492 27084 12587 27112
rect 12492 27072 12498 27084
rect 12575 27081 12587 27084
rect 12621 27081 12633 27115
rect 13078 27112 13084 27124
rect 13039 27084 13084 27112
rect 12575 27075 12633 27081
rect 13078 27072 13084 27084
rect 13136 27072 13142 27124
rect 5258 27004 5264 27056
rect 5316 27044 5322 27056
rect 7745 27047 7803 27053
rect 7745 27044 7757 27047
rect 5316 27016 7757 27044
rect 5316 27004 5322 27016
rect 7745 27013 7757 27016
rect 7791 27013 7803 27047
rect 7745 27007 7803 27013
rect 4982 26908 4988 26920
rect 4943 26880 4988 26908
rect 4982 26868 4988 26880
rect 5040 26868 5046 26920
rect 6825 26911 6883 26917
rect 6825 26908 6837 26911
rect 6564 26880 6837 26908
rect 4798 26800 4804 26852
rect 4856 26840 4862 26852
rect 5306 26843 5364 26849
rect 5306 26840 5318 26843
rect 4856 26812 5318 26840
rect 4856 26800 4862 26812
rect 5306 26809 5318 26812
rect 5352 26809 5364 26843
rect 5306 26803 5364 26809
rect 6086 26800 6092 26852
rect 6144 26840 6150 26852
rect 6564 26849 6592 26880
rect 6825 26877 6837 26880
rect 6871 26877 6883 26911
rect 7760 26908 7788 27007
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26976 8723 26979
rect 9674 26976 9680 26988
rect 8711 26948 9680 26976
rect 8711 26945 8723 26948
rect 8665 26939 8723 26945
rect 9674 26936 9680 26948
rect 9732 26936 9738 26988
rect 10505 26979 10563 26985
rect 10505 26945 10517 26979
rect 10551 26976 10563 26979
rect 10870 26976 10876 26988
rect 10551 26948 10876 26976
rect 10551 26945 10563 26948
rect 10505 26939 10563 26945
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 7926 26908 7932 26920
rect 7760 26880 7932 26908
rect 6825 26871 6883 26877
rect 7926 26868 7932 26880
rect 7984 26868 7990 26920
rect 8386 26868 8392 26920
rect 8444 26908 8450 26920
rect 8481 26911 8539 26917
rect 8481 26908 8493 26911
rect 8444 26880 8493 26908
rect 8444 26868 8450 26880
rect 8481 26877 8493 26880
rect 8527 26908 8539 26911
rect 8527 26880 8892 26908
rect 8527 26877 8539 26880
rect 8481 26871 8539 26877
rect 6549 26843 6607 26849
rect 6549 26840 6561 26843
rect 6144 26812 6561 26840
rect 6144 26800 6150 26812
rect 6549 26809 6561 26812
rect 6595 26809 6607 26843
rect 6549 26803 6607 26809
rect 8864 26784 8892 26880
rect 11422 26868 11428 26920
rect 11480 26908 11486 26920
rect 12161 26911 12219 26917
rect 12161 26908 12173 26911
rect 11480 26880 12173 26908
rect 11480 26868 11486 26880
rect 12161 26877 12173 26880
rect 12207 26908 12219 26911
rect 12472 26911 12530 26917
rect 12472 26908 12484 26911
rect 12207 26880 12484 26908
rect 12207 26877 12219 26880
rect 12161 26871 12219 26877
rect 12472 26877 12484 26880
rect 12518 26877 12530 26911
rect 12472 26871 12530 26877
rect 10594 26800 10600 26852
rect 10652 26840 10658 26852
rect 11149 26843 11207 26849
rect 10652 26812 10697 26840
rect 10652 26800 10658 26812
rect 11149 26809 11161 26843
rect 11195 26840 11207 26843
rect 11238 26840 11244 26852
rect 11195 26812 11244 26840
rect 11195 26809 11207 26812
rect 11149 26803 11207 26809
rect 11238 26800 11244 26812
rect 11296 26800 11302 26852
rect 4706 26732 4712 26784
rect 4764 26772 4770 26784
rect 4893 26775 4951 26781
rect 4893 26772 4905 26775
rect 4764 26744 4905 26772
rect 4764 26732 4770 26744
rect 4893 26741 4905 26744
rect 4939 26772 4951 26775
rect 5994 26772 6000 26784
rect 4939 26744 6000 26772
rect 4939 26741 4951 26744
rect 4893 26735 4951 26741
rect 5994 26732 6000 26744
rect 6052 26772 6058 26784
rect 7098 26772 7104 26784
rect 6052 26744 7104 26772
rect 6052 26732 6058 26744
rect 7098 26732 7104 26744
rect 7156 26732 7162 26784
rect 7374 26772 7380 26784
rect 7335 26744 7380 26772
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 8846 26732 8852 26784
rect 8904 26772 8910 26784
rect 8941 26775 8999 26781
rect 8941 26772 8953 26775
rect 8904 26744 8953 26772
rect 8904 26732 8910 26744
rect 8941 26741 8953 26744
rect 8987 26772 8999 26775
rect 9309 26775 9367 26781
rect 9309 26772 9321 26775
rect 8987 26744 9321 26772
rect 8987 26741 8999 26744
rect 8941 26735 8999 26741
rect 9309 26741 9321 26744
rect 9355 26741 9367 26775
rect 9309 26735 9367 26741
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 10045 26571 10103 26577
rect 10045 26537 10057 26571
rect 10091 26568 10103 26571
rect 10134 26568 10140 26580
rect 10091 26540 10140 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 10134 26528 10140 26540
rect 10192 26528 10198 26580
rect 10413 26571 10471 26577
rect 10413 26537 10425 26571
rect 10459 26568 10471 26571
rect 10594 26568 10600 26580
rect 10459 26540 10600 26568
rect 10459 26537 10471 26540
rect 10413 26531 10471 26537
rect 10594 26528 10600 26540
rect 10652 26528 10658 26580
rect 11514 26568 11520 26580
rect 11475 26540 11520 26568
rect 11514 26528 11520 26540
rect 11572 26568 11578 26580
rect 12207 26571 12265 26577
rect 12207 26568 12219 26571
rect 11572 26540 12219 26568
rect 11572 26528 11578 26540
rect 12207 26537 12219 26540
rect 12253 26537 12265 26571
rect 12207 26531 12265 26537
rect 5534 26500 5540 26512
rect 5495 26472 5540 26500
rect 5534 26460 5540 26472
rect 5592 26460 5598 26512
rect 10686 26500 10692 26512
rect 10647 26472 10692 26500
rect 10686 26460 10692 26472
rect 10744 26460 10750 26512
rect 11238 26500 11244 26512
rect 11199 26472 11244 26500
rect 11238 26460 11244 26472
rect 11296 26460 11302 26512
rect 4890 26432 4896 26444
rect 4851 26404 4896 26432
rect 4890 26392 4896 26404
rect 4948 26392 4954 26444
rect 6454 26392 6460 26444
rect 6512 26432 6518 26444
rect 7009 26435 7067 26441
rect 7009 26432 7021 26435
rect 6512 26404 7021 26432
rect 6512 26392 6518 26404
rect 7009 26401 7021 26404
rect 7055 26432 7067 26435
rect 7190 26432 7196 26444
rect 7055 26404 7196 26432
rect 7055 26401 7067 26404
rect 7009 26395 7067 26401
rect 7190 26392 7196 26404
rect 7248 26432 7254 26444
rect 7742 26432 7748 26444
rect 7248 26404 7748 26432
rect 7248 26392 7254 26404
rect 7742 26392 7748 26404
rect 7800 26392 7806 26444
rect 8110 26432 8116 26444
rect 8071 26404 8116 26432
rect 8110 26392 8116 26404
rect 8168 26392 8174 26444
rect 8573 26435 8631 26441
rect 8573 26401 8585 26435
rect 8619 26432 8631 26435
rect 8846 26432 8852 26444
rect 8619 26404 8852 26432
rect 8619 26401 8631 26404
rect 8573 26395 8631 26401
rect 7837 26367 7895 26373
rect 7837 26333 7849 26367
rect 7883 26364 7895 26367
rect 8588 26364 8616 26395
rect 8846 26392 8852 26404
rect 8904 26392 8910 26444
rect 12066 26392 12072 26444
rect 12124 26441 12130 26444
rect 12124 26435 12162 26441
rect 12150 26401 12162 26435
rect 12124 26395 12162 26401
rect 12124 26392 12130 26395
rect 8754 26364 8760 26376
rect 7883 26336 8616 26364
rect 8715 26336 8760 26364
rect 7883 26333 7895 26336
rect 7837 26327 7895 26333
rect 8754 26324 8760 26336
rect 8812 26324 8818 26376
rect 10597 26367 10655 26373
rect 10597 26333 10609 26367
rect 10643 26364 10655 26367
rect 10778 26364 10784 26376
rect 10643 26336 10784 26364
rect 10643 26333 10655 26336
rect 10597 26327 10655 26333
rect 10778 26324 10784 26336
rect 10836 26324 10842 26376
rect 4709 26299 4767 26305
rect 4709 26265 4721 26299
rect 4755 26296 4767 26299
rect 4982 26296 4988 26308
rect 4755 26268 4988 26296
rect 4755 26265 4767 26268
rect 4709 26259 4767 26265
rect 4982 26256 4988 26268
rect 5040 26296 5046 26308
rect 6822 26296 6828 26308
rect 5040 26268 5488 26296
rect 6783 26268 6828 26296
rect 5040 26256 5046 26268
rect 5460 26228 5488 26268
rect 6822 26256 6828 26268
rect 6880 26256 6886 26308
rect 5534 26228 5540 26240
rect 5460 26200 5540 26228
rect 5534 26188 5540 26200
rect 5592 26188 5598 26240
rect 5810 26228 5816 26240
rect 5771 26200 5816 26228
rect 5810 26188 5816 26200
rect 5868 26188 5874 26240
rect 9401 26231 9459 26237
rect 9401 26197 9413 26231
rect 9447 26228 9459 26231
rect 9582 26228 9588 26240
rect 9447 26200 9588 26228
rect 9447 26197 9459 26200
rect 9401 26191 9459 26197
rect 9582 26188 9588 26200
rect 9640 26188 9646 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 4890 26024 4896 26036
rect 4851 25996 4896 26024
rect 4890 25984 4896 25996
rect 4948 25984 4954 26036
rect 6454 26024 6460 26036
rect 6415 25996 6460 26024
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 10229 26027 10287 26033
rect 10229 25993 10241 26027
rect 10275 26024 10287 26027
rect 10594 26024 10600 26036
rect 10275 25996 10600 26024
rect 10275 25993 10287 25996
rect 10229 25987 10287 25993
rect 10594 25984 10600 25996
rect 10652 25984 10658 26036
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 10873 26027 10931 26033
rect 10873 26024 10885 26027
rect 10744 25996 10885 26024
rect 10744 25984 10750 25996
rect 10873 25993 10885 25996
rect 10919 25993 10931 26027
rect 10873 25987 10931 25993
rect 11471 26027 11529 26033
rect 11471 25993 11483 26027
rect 11517 26024 11529 26027
rect 11974 26024 11980 26036
rect 11517 25996 11980 26024
rect 11517 25993 11529 25996
rect 11471 25987 11529 25993
rect 11974 25984 11980 25996
rect 12032 25984 12038 26036
rect 12066 25984 12072 26036
rect 12124 26024 12130 26036
rect 12124 25996 12169 26024
rect 12124 25984 12130 25996
rect 5905 25891 5963 25897
rect 5905 25857 5917 25891
rect 5951 25888 5963 25891
rect 6086 25888 6092 25900
rect 5951 25860 6092 25888
rect 5951 25857 5963 25860
rect 5905 25851 5963 25857
rect 6086 25848 6092 25860
rect 6144 25848 6150 25900
rect 9309 25891 9367 25897
rect 9309 25857 9321 25891
rect 9355 25888 9367 25891
rect 9582 25888 9588 25900
rect 9355 25860 9588 25888
rect 9355 25857 9367 25860
rect 9309 25851 9367 25857
rect 9582 25848 9588 25860
rect 9640 25848 9646 25900
rect 11514 25848 11520 25900
rect 11572 25888 11578 25900
rect 12084 25888 12112 25984
rect 11572 25860 12112 25888
rect 11572 25848 11578 25860
rect 4525 25823 4583 25829
rect 4525 25789 4537 25823
rect 4571 25820 4583 25823
rect 5166 25820 5172 25832
rect 4571 25792 5172 25820
rect 4571 25789 4583 25792
rect 4525 25783 4583 25789
rect 5166 25780 5172 25792
rect 5224 25820 5230 25832
rect 5537 25823 5595 25829
rect 5537 25820 5549 25823
rect 5224 25792 5549 25820
rect 5224 25780 5230 25792
rect 5537 25789 5549 25792
rect 5583 25820 5595 25823
rect 5810 25820 5816 25832
rect 5583 25792 5816 25820
rect 5583 25789 5595 25792
rect 5537 25783 5595 25789
rect 5810 25780 5816 25792
rect 5868 25780 5874 25832
rect 6914 25780 6920 25832
rect 6972 25820 6978 25832
rect 7653 25823 7711 25829
rect 7653 25820 7665 25823
rect 6972 25792 7665 25820
rect 6972 25780 6978 25792
rect 7653 25789 7665 25792
rect 7699 25820 7711 25823
rect 8018 25820 8024 25832
rect 7699 25792 8024 25820
rect 7699 25789 7711 25792
rect 7653 25783 7711 25789
rect 8018 25780 8024 25792
rect 8076 25780 8082 25832
rect 8297 25823 8355 25829
rect 8297 25789 8309 25823
rect 8343 25789 8355 25823
rect 8297 25783 8355 25789
rect 5353 25755 5411 25761
rect 5353 25721 5365 25755
rect 5399 25721 5411 25755
rect 5353 25715 5411 25721
rect 5258 25684 5264 25696
rect 5219 25656 5264 25684
rect 5258 25644 5264 25656
rect 5316 25684 5322 25696
rect 5368 25684 5396 25715
rect 5316 25656 5396 25684
rect 8312 25684 8340 25783
rect 11238 25780 11244 25832
rect 11296 25820 11302 25832
rect 11368 25823 11426 25829
rect 11368 25820 11380 25823
rect 11296 25792 11380 25820
rect 11296 25780 11302 25792
rect 11368 25789 11380 25792
rect 11414 25789 11426 25823
rect 11368 25783 11426 25789
rect 8481 25755 8539 25761
rect 8481 25721 8493 25755
rect 8527 25752 8539 25755
rect 9398 25752 9404 25764
rect 8527 25724 9404 25752
rect 8527 25721 8539 25724
rect 8481 25715 8539 25721
rect 9398 25712 9404 25724
rect 9456 25712 9462 25764
rect 9671 25755 9729 25761
rect 9671 25721 9683 25755
rect 9717 25721 9729 25755
rect 9671 25715 9729 25721
rect 8846 25684 8852 25696
rect 8312 25656 8852 25684
rect 5316 25644 5322 25656
rect 8846 25644 8852 25656
rect 8904 25644 8910 25696
rect 9217 25687 9275 25693
rect 9217 25653 9229 25687
rect 9263 25684 9275 25687
rect 9692 25684 9720 25715
rect 9766 25684 9772 25696
rect 9263 25656 9772 25684
rect 9263 25653 9275 25656
rect 9217 25647 9275 25653
rect 9766 25644 9772 25656
rect 9824 25684 9830 25696
rect 10042 25684 10048 25696
rect 9824 25656 10048 25684
rect 9824 25644 9830 25656
rect 10042 25644 10048 25656
rect 10100 25644 10106 25696
rect 10597 25687 10655 25693
rect 10597 25653 10609 25687
rect 10643 25684 10655 25687
rect 10778 25684 10784 25696
rect 10643 25656 10784 25684
rect 10643 25653 10655 25656
rect 10597 25647 10655 25653
rect 10778 25644 10784 25656
rect 10836 25644 10842 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 5534 25480 5540 25492
rect 5495 25452 5540 25480
rect 5534 25440 5540 25452
rect 5592 25440 5598 25492
rect 5810 25440 5816 25492
rect 5868 25480 5874 25492
rect 6641 25483 6699 25489
rect 6641 25480 6653 25483
rect 5868 25452 6653 25480
rect 5868 25440 5874 25452
rect 6641 25449 6653 25452
rect 6687 25449 6699 25483
rect 6641 25443 6699 25449
rect 6914 25440 6920 25492
rect 6972 25480 6978 25492
rect 7009 25483 7067 25489
rect 7009 25480 7021 25483
rect 6972 25452 7021 25480
rect 6972 25440 6978 25452
rect 7009 25449 7021 25452
rect 7055 25449 7067 25483
rect 7009 25443 7067 25449
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 9033 25483 9091 25489
rect 9033 25480 9045 25483
rect 8812 25452 9045 25480
rect 8812 25440 8818 25452
rect 9033 25449 9045 25452
rect 9079 25449 9091 25483
rect 9398 25480 9404 25492
rect 9359 25452 9404 25480
rect 9033 25443 9091 25449
rect 9398 25440 9404 25452
rect 9456 25440 9462 25492
rect 10597 25483 10655 25489
rect 10597 25449 10609 25483
rect 10643 25480 10655 25483
rect 10686 25480 10692 25492
rect 10643 25452 10692 25480
rect 10643 25449 10655 25452
rect 10597 25443 10655 25449
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 10778 25440 10784 25492
rect 10836 25480 10842 25492
rect 11425 25483 11483 25489
rect 11425 25480 11437 25483
rect 10836 25452 11437 25480
rect 10836 25440 10842 25452
rect 11425 25449 11437 25452
rect 11471 25449 11483 25483
rect 11425 25443 11483 25449
rect 5169 25415 5227 25421
rect 5169 25381 5181 25415
rect 5215 25412 5227 25415
rect 5215 25384 6132 25412
rect 5215 25381 5227 25384
rect 5169 25375 5227 25381
rect 6104 25356 6132 25384
rect 7098 25372 7104 25424
rect 7156 25412 7162 25424
rect 7156 25384 7328 25412
rect 7156 25372 7162 25384
rect 7300 25356 7328 25384
rect 5537 25347 5595 25353
rect 5537 25313 5549 25347
rect 5583 25344 5595 25347
rect 5810 25344 5816 25356
rect 5583 25316 5816 25344
rect 5583 25313 5595 25316
rect 5537 25307 5595 25313
rect 5810 25304 5816 25316
rect 5868 25304 5874 25356
rect 6086 25344 6092 25356
rect 5999 25316 6092 25344
rect 6086 25304 6092 25316
rect 6144 25344 6150 25356
rect 7193 25347 7251 25353
rect 7193 25344 7205 25347
rect 6144 25316 7205 25344
rect 6144 25304 6150 25316
rect 7193 25313 7205 25316
rect 7239 25313 7251 25347
rect 7193 25307 7251 25313
rect 7282 25304 7288 25356
rect 7340 25344 7346 25356
rect 9416 25344 9444 25440
rect 10042 25421 10048 25424
rect 10039 25412 10048 25421
rect 10003 25384 10048 25412
rect 10039 25375 10048 25384
rect 10042 25372 10048 25375
rect 10100 25372 10106 25424
rect 10870 25412 10876 25424
rect 10831 25384 10876 25412
rect 10870 25372 10876 25384
rect 10928 25372 10934 25424
rect 11238 25372 11244 25424
rect 11296 25412 11302 25424
rect 11885 25415 11943 25421
rect 11885 25412 11897 25415
rect 11296 25384 11897 25412
rect 11296 25372 11302 25384
rect 11885 25381 11897 25384
rect 11931 25381 11943 25415
rect 11885 25375 11943 25381
rect 9677 25347 9735 25353
rect 9677 25344 9689 25347
rect 7340 25316 7433 25344
rect 9416 25316 9689 25344
rect 7340 25304 7346 25316
rect 9677 25313 9689 25316
rect 9723 25313 9735 25347
rect 9677 25307 9735 25313
rect 6178 25276 6184 25288
rect 6139 25248 6184 25276
rect 6178 25236 6184 25248
rect 6236 25236 6242 25288
rect 4430 25208 4436 25220
rect 4343 25180 4436 25208
rect 4430 25168 4436 25180
rect 4488 25208 4494 25220
rect 5442 25208 5448 25220
rect 4488 25180 5448 25208
rect 4488 25168 4494 25180
rect 5442 25168 5448 25180
rect 5500 25168 5506 25220
rect 4801 25143 4859 25149
rect 4801 25109 4813 25143
rect 4847 25140 4859 25143
rect 5166 25140 5172 25152
rect 4847 25112 5172 25140
rect 4847 25109 4859 25112
rect 4801 25103 4859 25109
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 7834 25100 7840 25152
rect 7892 25140 7898 25152
rect 8110 25140 8116 25152
rect 7892 25112 8116 25140
rect 7892 25100 7898 25112
rect 8110 25100 8116 25112
rect 8168 25140 8174 25152
rect 8297 25143 8355 25149
rect 8297 25140 8309 25143
rect 8168 25112 8309 25140
rect 8168 25100 8174 25112
rect 8297 25109 8309 25112
rect 8343 25109 8355 25143
rect 8297 25103 8355 25109
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 6914 24896 6920 24948
rect 6972 24936 6978 24948
rect 7147 24939 7205 24945
rect 7147 24936 7159 24939
rect 6972 24908 7159 24936
rect 6972 24896 6978 24908
rect 7147 24905 7159 24908
rect 7193 24905 7205 24939
rect 7147 24899 7205 24905
rect 7282 24896 7288 24948
rect 7340 24936 7346 24948
rect 8021 24939 8079 24945
rect 8021 24936 8033 24939
rect 7340 24908 8033 24936
rect 7340 24896 7346 24908
rect 8021 24905 8033 24908
rect 8067 24905 8079 24939
rect 8021 24899 8079 24905
rect 5442 24868 5448 24880
rect 5403 24840 5448 24868
rect 5442 24828 5448 24840
rect 5500 24828 5506 24880
rect 5077 24803 5135 24809
rect 5077 24769 5089 24803
rect 5123 24800 5135 24803
rect 5537 24803 5595 24809
rect 5537 24800 5549 24803
rect 5123 24772 5549 24800
rect 5123 24769 5135 24772
rect 5077 24763 5135 24769
rect 5537 24769 5549 24772
rect 5583 24800 5595 24803
rect 6641 24803 6699 24809
rect 6641 24800 6653 24803
rect 5583 24772 6653 24800
rect 5583 24769 5595 24772
rect 5537 24763 5595 24769
rect 6641 24769 6653 24772
rect 6687 24800 6699 24803
rect 7377 24803 7435 24809
rect 7377 24800 7389 24803
rect 6687 24772 7389 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 7377 24769 7389 24772
rect 7423 24800 7435 24803
rect 7558 24800 7564 24812
rect 7423 24772 7564 24800
rect 7423 24769 7435 24772
rect 7377 24763 7435 24769
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 7742 24800 7748 24812
rect 7703 24772 7748 24800
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 8202 24760 8208 24812
rect 8260 24800 8266 24812
rect 8570 24800 8576 24812
rect 8260 24772 8576 24800
rect 8260 24760 8266 24772
rect 8570 24760 8576 24772
rect 8628 24760 8634 24812
rect 8754 24760 8760 24812
rect 8812 24800 8818 24812
rect 9033 24803 9091 24809
rect 9033 24800 9045 24803
rect 8812 24772 9045 24800
rect 8812 24760 8818 24772
rect 9033 24769 9045 24772
rect 9079 24769 9091 24803
rect 10870 24800 10876 24812
rect 10831 24772 10876 24800
rect 9033 24763 9091 24769
rect 10870 24760 10876 24772
rect 10928 24760 10934 24812
rect 11238 24800 11244 24812
rect 11199 24772 11244 24800
rect 11238 24760 11244 24772
rect 11296 24760 11302 24812
rect 3970 24732 3976 24744
rect 3931 24704 3976 24732
rect 3970 24692 3976 24704
rect 4028 24692 4034 24744
rect 4338 24732 4344 24744
rect 4299 24704 4344 24732
rect 4338 24692 4344 24704
rect 4396 24692 4402 24744
rect 5350 24741 5356 24744
rect 5316 24735 5356 24741
rect 5316 24701 5328 24735
rect 5316 24695 5356 24701
rect 5350 24692 5356 24695
rect 5408 24692 5414 24744
rect 6914 24692 6920 24744
rect 6972 24732 6978 24744
rect 7239 24735 7297 24741
rect 7239 24732 7251 24735
rect 6972 24704 7251 24732
rect 6972 24692 6978 24704
rect 7239 24701 7251 24704
rect 7285 24732 7297 24735
rect 9953 24735 10011 24741
rect 7285 24704 8524 24732
rect 7285 24701 7297 24704
rect 7239 24695 7297 24701
rect 3142 24624 3148 24676
rect 3200 24664 3206 24676
rect 3697 24667 3755 24673
rect 3697 24664 3709 24667
rect 3200 24636 3709 24664
rect 3200 24624 3206 24636
rect 3697 24633 3709 24636
rect 3743 24664 3755 24667
rect 3789 24667 3847 24673
rect 3789 24664 3801 24667
rect 3743 24636 3801 24664
rect 3743 24633 3755 24636
rect 3697 24627 3755 24633
rect 3789 24633 3801 24636
rect 3835 24664 3847 24667
rect 4890 24664 4896 24676
rect 3835 24636 4896 24664
rect 3835 24633 3847 24636
rect 3789 24627 3847 24633
rect 4890 24624 4896 24636
rect 4948 24624 4954 24676
rect 5166 24664 5172 24676
rect 5127 24636 5172 24664
rect 5166 24624 5172 24636
rect 5224 24624 5230 24676
rect 5905 24667 5963 24673
rect 5905 24633 5917 24667
rect 5951 24664 5963 24667
rect 5994 24664 6000 24676
rect 5951 24636 6000 24664
rect 5951 24633 5963 24636
rect 5905 24627 5963 24633
rect 5994 24624 6000 24636
rect 6052 24624 6058 24676
rect 6273 24667 6331 24673
rect 6273 24633 6285 24667
rect 6319 24664 6331 24667
rect 7009 24667 7067 24673
rect 7009 24664 7021 24667
rect 6319 24636 7021 24664
rect 6319 24633 6331 24636
rect 6273 24627 6331 24633
rect 7009 24633 7021 24636
rect 7055 24664 7067 24667
rect 7098 24664 7104 24676
rect 7055 24636 7104 24664
rect 7055 24633 7067 24636
rect 7009 24627 7067 24633
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 4709 24599 4767 24605
rect 4709 24596 4721 24599
rect 4028 24568 4721 24596
rect 4028 24556 4034 24568
rect 4709 24565 4721 24568
rect 4755 24596 4767 24599
rect 5258 24596 5264 24608
rect 4755 24568 5264 24596
rect 4755 24565 4767 24568
rect 4709 24559 4767 24565
rect 5258 24556 5264 24568
rect 5316 24596 5322 24608
rect 6288 24596 6316 24627
rect 7098 24624 7104 24636
rect 7156 24624 7162 24676
rect 8496 24605 8524 24704
rect 9953 24701 9965 24735
rect 9999 24732 10011 24735
rect 10597 24735 10655 24741
rect 10597 24732 10609 24735
rect 9999 24704 10609 24732
rect 9999 24701 10011 24704
rect 9953 24695 10011 24701
rect 10597 24701 10609 24704
rect 10643 24701 10655 24735
rect 10597 24695 10655 24701
rect 9395 24667 9453 24673
rect 9395 24633 9407 24667
rect 9441 24664 9453 24667
rect 10042 24664 10048 24676
rect 9441 24636 10048 24664
rect 9441 24633 9453 24636
rect 9395 24627 9453 24633
rect 9508 24608 9536 24636
rect 10042 24624 10048 24636
rect 10100 24664 10106 24676
rect 10229 24667 10287 24673
rect 10229 24664 10241 24667
rect 10100 24636 10241 24664
rect 10100 24624 10106 24636
rect 10229 24633 10241 24636
rect 10275 24633 10287 24667
rect 10229 24627 10287 24633
rect 5316 24568 6316 24596
rect 8481 24599 8539 24605
rect 5316 24556 5322 24568
rect 8481 24565 8493 24599
rect 8527 24596 8539 24599
rect 8570 24596 8576 24608
rect 8527 24568 8576 24596
rect 8527 24565 8539 24568
rect 8481 24559 8539 24565
rect 8570 24556 8576 24568
rect 8628 24556 8634 24608
rect 8941 24599 8999 24605
rect 8941 24565 8953 24599
rect 8987 24596 8999 24599
rect 9490 24596 9496 24608
rect 8987 24568 9496 24596
rect 8987 24565 8999 24568
rect 8941 24559 8999 24565
rect 9490 24556 9496 24568
rect 9548 24556 9554 24608
rect 10612 24596 10640 24695
rect 10965 24667 11023 24673
rect 10965 24633 10977 24667
rect 11011 24633 11023 24667
rect 10965 24627 11023 24633
rect 10980 24596 11008 24627
rect 10612 24568 11008 24596
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 3142 24392 3148 24404
rect 2832 24364 3148 24392
rect 2832 24352 2838 24364
rect 3142 24352 3148 24364
rect 3200 24352 3206 24404
rect 3326 24352 3332 24404
rect 3384 24392 3390 24404
rect 3513 24395 3571 24401
rect 3513 24392 3525 24395
rect 3384 24364 3525 24392
rect 3384 24352 3390 24364
rect 3513 24361 3525 24364
rect 3559 24392 3571 24395
rect 4430 24392 4436 24404
rect 3559 24364 4436 24392
rect 3559 24361 3571 24364
rect 3513 24355 3571 24361
rect 4430 24352 4436 24364
rect 4488 24352 4494 24404
rect 5261 24395 5319 24401
rect 5261 24361 5273 24395
rect 5307 24392 5319 24395
rect 5350 24392 5356 24404
rect 5307 24364 5356 24392
rect 5307 24361 5319 24364
rect 5261 24355 5319 24361
rect 5350 24352 5356 24364
rect 5408 24392 5414 24404
rect 6641 24395 6699 24401
rect 6641 24392 6653 24395
rect 5408 24364 6653 24392
rect 5408 24352 5414 24364
rect 6641 24361 6653 24364
rect 6687 24392 6699 24395
rect 6822 24392 6828 24404
rect 6687 24364 6828 24392
rect 6687 24361 6699 24364
rect 6641 24355 6699 24361
rect 4154 24284 4160 24336
rect 4212 24324 4218 24336
rect 4212 24296 4292 24324
rect 4212 24284 4218 24296
rect 2958 24256 2964 24268
rect 2919 24228 2964 24256
rect 2958 24216 2964 24228
rect 3016 24216 3022 24268
rect 4264 24265 4292 24296
rect 4249 24259 4307 24265
rect 4249 24225 4261 24259
rect 4295 24225 4307 24259
rect 5718 24256 5724 24268
rect 5679 24228 5724 24256
rect 4249 24219 4307 24225
rect 5718 24216 5724 24228
rect 5776 24256 5782 24268
rect 6748 24265 6776 24364
rect 6822 24352 6828 24364
rect 6880 24352 6886 24404
rect 7190 24392 7196 24404
rect 7151 24364 7196 24392
rect 7190 24352 7196 24364
rect 7248 24352 7254 24404
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 9769 24395 9827 24401
rect 9769 24392 9781 24395
rect 9732 24364 9781 24392
rect 9732 24352 9738 24364
rect 9769 24361 9781 24364
rect 9815 24361 9827 24395
rect 9769 24355 9827 24361
rect 11238 24324 11244 24336
rect 11199 24296 11244 24324
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 6181 24259 6239 24265
rect 6181 24256 6193 24259
rect 5776 24228 6193 24256
rect 5776 24216 5782 24228
rect 6181 24225 6193 24228
rect 6227 24225 6239 24259
rect 6181 24219 6239 24225
rect 6733 24259 6791 24265
rect 6733 24225 6745 24259
rect 6779 24225 6791 24259
rect 6733 24219 6791 24225
rect 7009 24259 7067 24265
rect 7009 24225 7021 24259
rect 7055 24256 7067 24259
rect 7558 24256 7564 24268
rect 7055 24228 7564 24256
rect 7055 24225 7067 24228
rect 7009 24219 7067 24225
rect 7558 24216 7564 24228
rect 7616 24216 7622 24268
rect 7834 24256 7840 24268
rect 7795 24228 7840 24256
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 8294 24256 8300 24268
rect 8255 24228 8300 24256
rect 8294 24216 8300 24228
rect 8352 24216 8358 24268
rect 9674 24256 9680 24268
rect 9635 24228 9680 24256
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10134 24256 10140 24268
rect 10095 24228 10140 24256
rect 10134 24216 10140 24228
rect 10192 24216 10198 24268
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11333 24259 11391 24265
rect 11333 24256 11345 24259
rect 11112 24228 11345 24256
rect 11112 24216 11118 24228
rect 11333 24225 11345 24228
rect 11379 24256 11391 24259
rect 11379 24228 12572 24256
rect 11379 24225 11391 24228
rect 11333 24219 11391 24225
rect 4062 24148 4068 24200
rect 4120 24188 4126 24200
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 4120 24160 4169 24188
rect 4120 24148 4126 24160
rect 4157 24157 4169 24160
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 8570 24148 8576 24200
rect 8628 24188 8634 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 8628 24160 9137 24188
rect 8628 24148 8634 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 4338 24080 4344 24132
rect 4396 24120 4402 24132
rect 5534 24120 5540 24132
rect 4396 24092 5540 24120
rect 4396 24080 4402 24092
rect 5534 24080 5540 24092
rect 5592 24120 5598 24132
rect 5629 24123 5687 24129
rect 5629 24120 5641 24123
rect 5592 24092 5641 24120
rect 5592 24080 5598 24092
rect 5629 24089 5641 24092
rect 5675 24120 5687 24123
rect 6178 24120 6184 24132
rect 5675 24092 6184 24120
rect 5675 24089 5687 24092
rect 5629 24083 5687 24089
rect 6178 24080 6184 24092
rect 6236 24080 6242 24132
rect 6822 24120 6828 24132
rect 6783 24092 6828 24120
rect 6822 24080 6828 24092
rect 6880 24080 6886 24132
rect 8481 24123 8539 24129
rect 8481 24089 8493 24123
rect 8527 24120 8539 24123
rect 8846 24120 8852 24132
rect 8527 24092 8852 24120
rect 8527 24089 8539 24092
rect 8481 24083 8539 24089
rect 8846 24080 8852 24092
rect 8904 24120 8910 24132
rect 10134 24120 10140 24132
rect 8904 24092 10140 24120
rect 8904 24080 8910 24092
rect 10134 24080 10140 24092
rect 10192 24080 10198 24132
rect 10502 24080 10508 24132
rect 10560 24120 10566 24132
rect 11149 24123 11207 24129
rect 11149 24120 11161 24123
rect 10560 24092 11161 24120
rect 10560 24080 10566 24092
rect 11149 24089 11161 24092
rect 11195 24120 11207 24123
rect 12342 24120 12348 24132
rect 11195 24092 12348 24120
rect 11195 24089 11207 24092
rect 11149 24083 11207 24089
rect 12342 24080 12348 24092
rect 12400 24080 12406 24132
rect 5810 24012 5816 24064
rect 5868 24052 5874 24064
rect 5905 24055 5963 24061
rect 5905 24052 5917 24055
rect 5868 24024 5917 24052
rect 5868 24012 5874 24024
rect 5905 24021 5917 24024
rect 5951 24021 5963 24055
rect 5905 24015 5963 24021
rect 8757 24055 8815 24061
rect 8757 24021 8769 24055
rect 8803 24052 8815 24055
rect 9306 24052 9312 24064
rect 8803 24024 9312 24052
rect 8803 24021 8815 24024
rect 8757 24015 8815 24021
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 10594 24012 10600 24064
rect 10652 24052 10658 24064
rect 12544 24061 12572 24228
rect 10689 24055 10747 24061
rect 10689 24052 10701 24055
rect 10652 24024 10701 24052
rect 10652 24012 10658 24024
rect 10689 24021 10701 24024
rect 10735 24021 10747 24055
rect 10689 24015 10747 24021
rect 12529 24055 12587 24061
rect 12529 24021 12541 24055
rect 12575 24052 12587 24055
rect 12710 24052 12716 24064
rect 12575 24024 12716 24052
rect 12575 24021 12587 24024
rect 12529 24015 12587 24021
rect 12710 24012 12716 24024
rect 12768 24012 12774 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 2777 23851 2835 23857
rect 2777 23817 2789 23851
rect 2823 23848 2835 23851
rect 2958 23848 2964 23860
rect 2823 23820 2964 23848
rect 2823 23817 2835 23820
rect 2777 23811 2835 23817
rect 2958 23808 2964 23820
rect 3016 23808 3022 23860
rect 4338 23848 4344 23860
rect 4299 23820 4344 23848
rect 4338 23808 4344 23820
rect 4396 23808 4402 23860
rect 6641 23851 6699 23857
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 6822 23848 6828 23860
rect 6687 23820 6828 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 6822 23808 6828 23820
rect 6880 23848 6886 23860
rect 7377 23851 7435 23857
rect 7377 23848 7389 23851
rect 6880 23820 7389 23848
rect 6880 23808 6886 23820
rect 7377 23817 7389 23820
rect 7423 23848 7435 23851
rect 8202 23848 8208 23860
rect 7423 23820 8208 23848
rect 7423 23817 7435 23820
rect 7377 23811 7435 23817
rect 8202 23808 8208 23820
rect 8260 23848 8266 23860
rect 8941 23851 8999 23857
rect 8941 23848 8953 23851
rect 8260 23820 8953 23848
rect 8260 23808 8266 23820
rect 8941 23817 8953 23820
rect 8987 23848 8999 23851
rect 9582 23848 9588 23860
rect 8987 23820 9588 23848
rect 8987 23817 8999 23820
rect 8941 23811 8999 23817
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 10134 23848 10140 23860
rect 10095 23820 10140 23848
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 11054 23808 11060 23860
rect 11112 23848 11118 23860
rect 11425 23851 11483 23857
rect 11425 23848 11437 23851
rect 11112 23820 11437 23848
rect 11112 23808 11118 23820
rect 11425 23817 11437 23820
rect 11471 23817 11483 23851
rect 12710 23848 12716 23860
rect 12671 23820 12716 23848
rect 11425 23811 11483 23817
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 3326 23780 3332 23792
rect 3287 23752 3332 23780
rect 3326 23740 3332 23752
rect 3384 23740 3390 23792
rect 7282 23789 7288 23792
rect 7266 23783 7288 23789
rect 7266 23749 7278 23783
rect 7340 23780 7346 23792
rect 8481 23783 8539 23789
rect 8481 23780 8493 23783
rect 7340 23752 8493 23780
rect 7266 23743 7288 23749
rect 7282 23740 7288 23743
rect 7340 23740 7346 23752
rect 8481 23749 8493 23752
rect 8527 23780 8539 23783
rect 8754 23780 8760 23792
rect 8527 23752 8760 23780
rect 8527 23749 8539 23752
rect 8481 23743 8539 23749
rect 8754 23740 8760 23752
rect 8812 23789 8818 23792
rect 8812 23783 8861 23789
rect 8812 23749 8815 23783
rect 8849 23749 8861 23783
rect 9306 23780 9312 23792
rect 8812 23743 8861 23749
rect 9048 23752 9312 23780
rect 8812 23740 8818 23743
rect 3970 23712 3976 23724
rect 3931 23684 3976 23712
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 4706 23712 4712 23724
rect 4619 23684 4712 23712
rect 4706 23672 4712 23684
rect 4764 23712 4770 23724
rect 5534 23712 5540 23724
rect 4764 23684 5396 23712
rect 5495 23684 5540 23712
rect 4764 23672 4770 23684
rect 3145 23647 3203 23653
rect 3145 23613 3157 23647
rect 3191 23644 3203 23647
rect 3234 23644 3240 23656
rect 3191 23616 3240 23644
rect 3191 23613 3203 23616
rect 3145 23607 3203 23613
rect 3234 23604 3240 23616
rect 3292 23604 3298 23656
rect 3510 23644 3516 23656
rect 3471 23616 3516 23644
rect 3510 23604 3516 23616
rect 3568 23604 3574 23656
rect 4982 23644 4988 23656
rect 4943 23616 4988 23644
rect 4982 23604 4988 23616
rect 5040 23604 5046 23656
rect 5368 23644 5396 23684
rect 5534 23672 5540 23684
rect 5592 23672 5598 23724
rect 6273 23715 6331 23721
rect 6273 23681 6285 23715
rect 6319 23712 6331 23715
rect 7469 23715 7527 23721
rect 7469 23712 7481 23715
rect 6319 23684 7481 23712
rect 6319 23681 6331 23684
rect 6273 23675 6331 23681
rect 7469 23681 7481 23684
rect 7515 23712 7527 23715
rect 7558 23712 7564 23724
rect 7515 23684 7564 23712
rect 7515 23681 7527 23684
rect 7469 23675 7527 23681
rect 7558 23672 7564 23684
rect 7616 23712 7622 23724
rect 9048 23721 9076 23752
rect 9306 23740 9312 23752
rect 9364 23780 9370 23792
rect 12618 23789 12624 23792
rect 12602 23783 12624 23789
rect 9364 23752 11928 23780
rect 9364 23740 9370 23752
rect 9033 23715 9091 23721
rect 9033 23712 9045 23715
rect 7616 23684 9045 23712
rect 7616 23672 7622 23684
rect 9033 23681 9045 23684
rect 9079 23681 9091 23715
rect 10502 23712 10508 23724
rect 10463 23684 10508 23712
rect 9033 23675 9091 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 11900 23721 11928 23752
rect 12602 23749 12614 23783
rect 12602 23743 12624 23749
rect 12618 23740 12624 23743
rect 12676 23740 12682 23792
rect 11885 23715 11943 23721
rect 11885 23681 11897 23715
rect 11931 23712 11943 23715
rect 12805 23715 12863 23721
rect 12805 23712 12817 23715
rect 11931 23684 12817 23712
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 12805 23681 12817 23684
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 5629 23647 5687 23653
rect 5629 23644 5641 23647
rect 5368 23616 5641 23644
rect 5629 23613 5641 23616
rect 5675 23644 5687 23647
rect 5718 23644 5724 23656
rect 5675 23616 5724 23644
rect 5675 23613 5687 23616
rect 5629 23607 5687 23613
rect 5718 23604 5724 23616
rect 5776 23604 5782 23656
rect 7101 23647 7159 23653
rect 7101 23613 7113 23647
rect 7147 23644 7159 23647
rect 7834 23644 7840 23656
rect 7147 23616 7840 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 3970 23536 3976 23588
rect 4028 23576 4034 23588
rect 5166 23576 5172 23588
rect 4028 23548 5172 23576
rect 4028 23536 4034 23548
rect 5166 23536 5172 23548
rect 5224 23576 5230 23588
rect 7116 23576 7144 23607
rect 7834 23604 7840 23616
rect 7892 23604 7898 23656
rect 8570 23604 8576 23656
rect 8628 23644 8634 23656
rect 8665 23647 8723 23653
rect 8665 23644 8677 23647
rect 8628 23616 8677 23644
rect 8628 23604 8634 23616
rect 8665 23613 8677 23616
rect 8711 23613 8723 23647
rect 8665 23607 8723 23613
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 12032 23616 12173 23644
rect 12032 23604 12038 23616
rect 12161 23613 12173 23616
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 12526 23644 12532 23656
rect 12483 23616 12532 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12526 23604 12532 23616
rect 12584 23604 12590 23656
rect 9398 23576 9404 23588
rect 5224 23548 7144 23576
rect 9359 23548 9404 23576
rect 5224 23536 5230 23548
rect 9398 23536 9404 23548
rect 9456 23536 9462 23588
rect 10502 23536 10508 23588
rect 10560 23576 10566 23588
rect 10597 23579 10655 23585
rect 10597 23576 10609 23579
rect 10560 23548 10609 23576
rect 10560 23536 10566 23548
rect 10597 23545 10609 23548
rect 10643 23545 10655 23579
rect 10597 23539 10655 23545
rect 11149 23579 11207 23585
rect 11149 23545 11161 23579
rect 11195 23576 11207 23579
rect 12342 23576 12348 23588
rect 11195 23548 12348 23576
rect 11195 23545 11207 23548
rect 11149 23539 11207 23545
rect 12342 23536 12348 23548
rect 12400 23536 12406 23588
rect 4890 23508 4896 23520
rect 4851 23480 4896 23508
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 7745 23511 7803 23517
rect 7745 23477 7757 23511
rect 7791 23508 7803 23511
rect 7834 23508 7840 23520
rect 7791 23480 7840 23508
rect 7791 23477 7803 23480
rect 7745 23471 7803 23477
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 9674 23508 9680 23520
rect 9635 23480 9680 23508
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 13078 23508 13084 23520
rect 13039 23480 13084 23508
rect 13078 23468 13084 23480
rect 13136 23468 13142 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 3881 23307 3939 23313
rect 3881 23273 3893 23307
rect 3927 23304 3939 23307
rect 4154 23304 4160 23316
rect 3927 23276 4160 23304
rect 3927 23273 3939 23276
rect 3881 23267 3939 23273
rect 4154 23264 4160 23276
rect 4212 23264 4218 23316
rect 5534 23304 5540 23316
rect 5495 23276 5540 23304
rect 5534 23264 5540 23276
rect 5592 23264 5598 23316
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 6822 23304 6828 23316
rect 5960 23276 6592 23304
rect 6783 23276 6828 23304
rect 5960 23264 5966 23276
rect 2590 23168 2596 23180
rect 2551 23140 2596 23168
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 3970 23168 3976 23180
rect 2832 23140 3976 23168
rect 2832 23128 2838 23140
rect 3970 23128 3976 23140
rect 4028 23128 4034 23180
rect 4132 23171 4190 23177
rect 4132 23137 4144 23171
rect 4178 23168 4190 23171
rect 4522 23168 4528 23180
rect 4178 23140 4528 23168
rect 4178 23137 4190 23140
rect 4132 23131 4190 23137
rect 4522 23128 4528 23140
rect 4580 23128 4586 23180
rect 4893 23171 4951 23177
rect 4893 23137 4905 23171
rect 4939 23168 4951 23171
rect 4982 23168 4988 23180
rect 4939 23140 4988 23168
rect 4939 23137 4951 23140
rect 4893 23131 4951 23137
rect 4982 23128 4988 23140
rect 5040 23168 5046 23180
rect 5537 23171 5595 23177
rect 5537 23168 5549 23171
rect 5040 23140 5549 23168
rect 5040 23128 5046 23140
rect 5537 23137 5549 23140
rect 5583 23168 5595 23171
rect 5902 23168 5908 23180
rect 5583 23140 5908 23168
rect 5583 23137 5595 23140
rect 5537 23131 5595 23137
rect 5902 23128 5908 23140
rect 5960 23128 5966 23180
rect 6086 23168 6092 23180
rect 6047 23140 6092 23168
rect 6086 23128 6092 23140
rect 6144 23128 6150 23180
rect 6270 23168 6276 23180
rect 6231 23140 6276 23168
rect 6270 23128 6276 23140
rect 6328 23128 6334 23180
rect 6564 23168 6592 23276
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 7193 23307 7251 23313
rect 7193 23273 7205 23307
rect 7239 23304 7251 23307
rect 7282 23304 7288 23316
rect 7239 23276 7288 23304
rect 7239 23273 7251 23276
rect 7193 23267 7251 23273
rect 7282 23264 7288 23276
rect 7340 23264 7346 23316
rect 7558 23304 7564 23316
rect 7519 23276 7564 23304
rect 7558 23264 7564 23276
rect 7616 23264 7622 23316
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 9033 23307 9091 23313
rect 9033 23304 9045 23307
rect 8352 23276 9045 23304
rect 8352 23264 8358 23276
rect 9033 23273 9045 23276
rect 9079 23273 9091 23307
rect 9033 23267 9091 23273
rect 12526 23264 12532 23316
rect 12584 23304 12590 23316
rect 12713 23307 12771 23313
rect 12713 23304 12725 23307
rect 12584 23276 12725 23304
rect 12584 23264 12590 23276
rect 12713 23273 12725 23276
rect 12759 23273 12771 23307
rect 12713 23267 12771 23273
rect 10502 23236 10508 23248
rect 10463 23208 10508 23236
rect 10502 23196 10508 23208
rect 10560 23196 10566 23248
rect 11885 23239 11943 23245
rect 11885 23205 11897 23239
rect 11931 23236 11943 23239
rect 11974 23236 11980 23248
rect 11931 23208 11980 23236
rect 11931 23205 11943 23208
rect 11885 23199 11943 23205
rect 11974 23196 11980 23208
rect 12032 23196 12038 23248
rect 6822 23168 6828 23180
rect 6564 23140 6828 23168
rect 6822 23128 6828 23140
rect 6880 23128 6886 23180
rect 7926 23128 7932 23180
rect 7984 23168 7990 23180
rect 8021 23171 8079 23177
rect 8021 23168 8033 23171
rect 7984 23140 8033 23168
rect 7984 23128 7990 23140
rect 8021 23137 8033 23140
rect 8067 23137 8079 23171
rect 8478 23168 8484 23180
rect 8439 23140 8484 23168
rect 8021 23131 8079 23137
rect 8478 23128 8484 23140
rect 8536 23128 8542 23180
rect 12066 23168 12072 23180
rect 12027 23140 12072 23168
rect 12066 23128 12072 23140
rect 12124 23128 12130 23180
rect 8754 23100 8760 23112
rect 8715 23072 8760 23100
rect 8754 23060 8760 23072
rect 8812 23060 8818 23112
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23100 10287 23103
rect 10410 23100 10416 23112
rect 10275 23072 10416 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 10410 23060 10416 23072
rect 10468 23060 10474 23112
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 11146 23100 11152 23112
rect 11103 23072 11152 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 11146 23060 11152 23072
rect 11204 23060 11210 23112
rect 4203 23035 4261 23041
rect 4203 23001 4215 23035
rect 4249 23032 4261 23035
rect 5626 23032 5632 23044
rect 4249 23004 5632 23032
rect 4249 23001 4261 23004
rect 4203 22995 4261 23001
rect 5626 22992 5632 23004
rect 5684 22992 5690 23044
rect 2869 22967 2927 22973
rect 2869 22933 2881 22967
rect 2915 22964 2927 22967
rect 2958 22964 2964 22976
rect 2915 22936 2964 22964
rect 2915 22933 2927 22936
rect 2869 22927 2927 22933
rect 2958 22924 2964 22936
rect 3016 22924 3022 22976
rect 3510 22964 3516 22976
rect 3471 22936 3516 22964
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 11054 22924 11060 22976
rect 11112 22964 11118 22976
rect 12161 22967 12219 22973
rect 12161 22964 12173 22967
rect 11112 22936 12173 22964
rect 11112 22924 11118 22936
rect 12161 22933 12173 22936
rect 12207 22933 12219 22967
rect 12161 22927 12219 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2225 22763 2283 22769
rect 2225 22729 2237 22763
rect 2271 22760 2283 22763
rect 2590 22760 2596 22772
rect 2271 22732 2596 22760
rect 2271 22729 2283 22732
rect 2225 22723 2283 22729
rect 2590 22720 2596 22732
rect 2648 22720 2654 22772
rect 5810 22760 5816 22772
rect 5771 22732 5816 22760
rect 5810 22720 5816 22732
rect 5868 22720 5874 22772
rect 5902 22720 5908 22772
rect 5960 22760 5966 22772
rect 6089 22763 6147 22769
rect 6089 22760 6101 22763
rect 5960 22732 6101 22760
rect 5960 22720 5966 22732
rect 6089 22729 6101 22732
rect 6135 22729 6147 22763
rect 6089 22723 6147 22729
rect 6270 22720 6276 22772
rect 6328 22760 6334 22772
rect 6457 22763 6515 22769
rect 6457 22760 6469 22763
rect 6328 22732 6469 22760
rect 6328 22720 6334 22732
rect 6457 22729 6469 22732
rect 6503 22729 6515 22763
rect 6457 22723 6515 22729
rect 7098 22720 7104 22772
rect 7156 22760 7162 22772
rect 7926 22760 7932 22772
rect 7156 22732 7932 22760
rect 7156 22720 7162 22732
rect 7926 22720 7932 22732
rect 7984 22760 7990 22772
rect 8021 22763 8079 22769
rect 8021 22760 8033 22763
rect 7984 22732 8033 22760
rect 7984 22720 7990 22732
rect 8021 22729 8033 22732
rect 8067 22729 8079 22763
rect 8021 22723 8079 22729
rect 11977 22763 12035 22769
rect 11977 22729 11989 22763
rect 12023 22760 12035 22763
rect 12066 22760 12072 22772
rect 12023 22732 12072 22760
rect 12023 22729 12035 22732
rect 11977 22723 12035 22729
rect 12066 22720 12072 22732
rect 12124 22720 12130 22772
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12575 22763 12633 22769
rect 12575 22760 12587 22763
rect 12492 22732 12587 22760
rect 12492 22720 12498 22732
rect 12575 22729 12587 22732
rect 12621 22729 12633 22763
rect 12575 22723 12633 22729
rect 12894 22720 12900 22772
rect 12952 22760 12958 22772
rect 13587 22763 13645 22769
rect 13587 22760 13599 22763
rect 12952 22732 13599 22760
rect 12952 22720 12958 22732
rect 13587 22729 13599 22732
rect 13633 22729 13645 22763
rect 13587 22723 13645 22729
rect 2501 22695 2559 22701
rect 2501 22661 2513 22695
rect 2547 22661 2559 22695
rect 3970 22692 3976 22704
rect 3931 22664 3976 22692
rect 2501 22655 2559 22661
rect 2516 22624 2544 22655
rect 3970 22652 3976 22664
rect 4028 22652 4034 22704
rect 7282 22692 7288 22704
rect 4724 22664 7288 22692
rect 4724 22624 4752 22664
rect 7282 22652 7288 22664
rect 7340 22692 7346 22704
rect 8389 22695 8447 22701
rect 8389 22692 8401 22695
rect 7340 22664 8401 22692
rect 7340 22652 7346 22664
rect 8389 22661 8401 22664
rect 8435 22692 8447 22695
rect 8478 22692 8484 22704
rect 8435 22664 8484 22692
rect 8435 22661 8447 22664
rect 8389 22655 8447 22661
rect 8478 22652 8484 22664
rect 8536 22652 8542 22704
rect 4890 22624 4896 22636
rect 2516 22596 4752 22624
rect 4851 22596 4896 22624
rect 4890 22584 4896 22596
rect 4948 22584 4954 22636
rect 6086 22584 6092 22636
rect 6144 22624 6150 22636
rect 6730 22624 6736 22636
rect 6144 22596 6736 22624
rect 6144 22584 6150 22596
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 7190 22624 7196 22636
rect 7151 22596 7196 22624
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 9033 22627 9091 22633
rect 9033 22624 9045 22627
rect 8812 22596 9045 22624
rect 8812 22584 8818 22596
rect 9033 22593 9045 22596
rect 9079 22593 9091 22627
rect 9033 22587 9091 22593
rect 10873 22627 10931 22633
rect 10873 22593 10885 22627
rect 10919 22624 10931 22627
rect 10962 22624 10968 22636
rect 10919 22596 10968 22624
rect 10919 22593 10931 22596
rect 10873 22587 10931 22593
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 11146 22624 11152 22636
rect 11107 22596 11152 22624
rect 11146 22584 11152 22596
rect 11204 22584 11210 22636
rect 2317 22559 2375 22565
rect 2317 22525 2329 22559
rect 2363 22525 2375 22559
rect 2317 22519 2375 22525
rect 2332 22488 2360 22519
rect 9674 22516 9680 22568
rect 9732 22556 9738 22568
rect 10321 22559 10379 22565
rect 10321 22556 10333 22559
rect 9732 22528 10333 22556
rect 9732 22516 9738 22528
rect 10321 22525 10333 22528
rect 10367 22556 10379 22559
rect 10502 22556 10508 22568
rect 10367 22528 10508 22556
rect 10367 22525 10379 22528
rect 10321 22519 10379 22525
rect 10502 22516 10508 22528
rect 10560 22516 10566 22568
rect 12158 22516 12164 22568
rect 12216 22556 12222 22568
rect 12472 22559 12530 22565
rect 12472 22556 12484 22559
rect 12216 22528 12484 22556
rect 12216 22516 12222 22528
rect 12472 22525 12484 22528
rect 12518 22556 12530 22559
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12518 22528 12909 22556
rect 12518 22525 12530 22528
rect 12472 22519 12530 22525
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 12897 22519 12955 22525
rect 13170 22516 13176 22568
rect 13228 22556 13234 22568
rect 13484 22559 13542 22565
rect 13484 22556 13496 22559
rect 13228 22528 13496 22556
rect 13228 22516 13234 22528
rect 13484 22525 13496 22528
rect 13530 22556 13542 22559
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 13530 22528 13921 22556
rect 13530 22525 13542 22528
rect 13484 22519 13542 22525
rect 13909 22525 13921 22528
rect 13955 22525 13967 22559
rect 13909 22519 13967 22525
rect 2869 22491 2927 22497
rect 2869 22488 2881 22491
rect 2332 22460 2881 22488
rect 2869 22457 2881 22460
rect 2915 22488 2927 22491
rect 3142 22488 3148 22500
rect 2915 22460 3148 22488
rect 2915 22457 2927 22460
rect 2869 22451 2927 22457
rect 3142 22448 3148 22460
rect 3200 22448 3206 22500
rect 3418 22488 3424 22500
rect 3379 22460 3424 22488
rect 3418 22448 3424 22460
rect 3476 22448 3482 22500
rect 3513 22491 3571 22497
rect 3513 22457 3525 22491
rect 3559 22488 3571 22491
rect 3878 22488 3884 22500
rect 3559 22460 3884 22488
rect 3559 22457 3571 22460
rect 3513 22451 3571 22457
rect 3237 22423 3295 22429
rect 3237 22389 3249 22423
rect 3283 22420 3295 22423
rect 3528 22420 3556 22451
rect 3878 22448 3884 22460
rect 3936 22448 3942 22500
rect 5258 22497 5264 22500
rect 4801 22491 4859 22497
rect 4801 22457 4813 22491
rect 4847 22488 4859 22491
rect 5214 22491 5264 22497
rect 5214 22488 5226 22491
rect 4847 22460 5226 22488
rect 4847 22457 4859 22460
rect 4801 22451 4859 22457
rect 5214 22457 5226 22460
rect 5260 22457 5264 22491
rect 5214 22451 5264 22457
rect 5258 22448 5264 22451
rect 5316 22488 5322 22500
rect 6914 22488 6920 22500
rect 5316 22460 5362 22488
rect 6875 22460 6920 22488
rect 5316 22448 5322 22460
rect 6914 22448 6920 22460
rect 6972 22448 6978 22500
rect 7009 22491 7067 22497
rect 7009 22457 7021 22491
rect 7055 22457 7067 22491
rect 7009 22451 7067 22457
rect 9354 22491 9412 22497
rect 9354 22457 9366 22491
rect 9400 22457 9412 22491
rect 10870 22488 10876 22500
rect 9354 22451 9412 22457
rect 9968 22460 10876 22488
rect 3283 22392 3556 22420
rect 4433 22423 4491 22429
rect 3283 22389 3295 22392
rect 3237 22383 3295 22389
rect 4433 22389 4445 22423
rect 4479 22420 4491 22423
rect 4522 22420 4528 22432
rect 4479 22392 4528 22420
rect 4479 22389 4491 22392
rect 4433 22383 4491 22389
rect 4522 22380 4528 22392
rect 4580 22380 4586 22432
rect 6822 22380 6828 22432
rect 6880 22420 6886 22432
rect 7024 22420 7052 22451
rect 6880 22392 7052 22420
rect 6880 22380 6886 22392
rect 7926 22380 7932 22432
rect 7984 22420 7990 22432
rect 8849 22423 8907 22429
rect 8849 22420 8861 22423
rect 7984 22392 8861 22420
rect 7984 22380 7990 22392
rect 8849 22389 8861 22392
rect 8895 22420 8907 22423
rect 9369 22420 9397 22451
rect 9490 22420 9496 22432
rect 8895 22392 9496 22420
rect 8895 22389 8907 22392
rect 8849 22383 8907 22389
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 9968 22429 9996 22460
rect 10870 22448 10876 22460
rect 10928 22488 10934 22500
rect 10965 22491 11023 22497
rect 10965 22488 10977 22491
rect 10928 22460 10977 22488
rect 10928 22448 10934 22460
rect 10965 22457 10977 22460
rect 11011 22457 11023 22491
rect 10965 22451 11023 22457
rect 9953 22423 10011 22429
rect 9953 22389 9965 22423
rect 9999 22389 10011 22423
rect 9953 22383 10011 22389
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 2685 22219 2743 22225
rect 2685 22185 2697 22219
rect 2731 22216 2743 22219
rect 2774 22216 2780 22228
rect 2731 22188 2780 22216
rect 2731 22185 2743 22188
rect 2685 22179 2743 22185
rect 2774 22176 2780 22188
rect 2832 22176 2838 22228
rect 3099 22219 3157 22225
rect 3099 22185 3111 22219
rect 3145 22216 3157 22219
rect 3418 22216 3424 22228
rect 3145 22188 3424 22216
rect 3145 22185 3157 22188
rect 3099 22179 3157 22185
rect 3418 22176 3424 22188
rect 3476 22176 3482 22228
rect 4525 22219 4583 22225
rect 4525 22185 4537 22219
rect 4571 22216 4583 22219
rect 4890 22216 4896 22228
rect 4571 22188 4896 22216
rect 4571 22185 4583 22188
rect 4525 22179 4583 22185
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 5810 22176 5816 22228
rect 5868 22216 5874 22228
rect 6641 22219 6699 22225
rect 6641 22216 6653 22219
rect 5868 22188 6653 22216
rect 5868 22176 5874 22188
rect 6641 22185 6653 22188
rect 6687 22216 6699 22219
rect 6822 22216 6828 22228
rect 6687 22188 6828 22216
rect 6687 22185 6699 22188
rect 6641 22179 6699 22185
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 7282 22176 7288 22228
rect 7340 22216 7346 22228
rect 7653 22219 7711 22225
rect 7653 22216 7665 22219
rect 7340 22188 7665 22216
rect 7340 22176 7346 22188
rect 7653 22185 7665 22188
rect 7699 22185 7711 22219
rect 7653 22179 7711 22185
rect 8754 22176 8760 22228
rect 8812 22216 8818 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8812 22188 9045 22216
rect 8812 22176 8818 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 9490 22176 9496 22228
rect 9548 22216 9554 22228
rect 9548 22188 9812 22216
rect 9548 22176 9554 22188
rect 5258 22108 5264 22160
rect 5316 22157 5322 22160
rect 5316 22151 5364 22157
rect 5316 22117 5318 22151
rect 5352 22117 5364 22151
rect 5316 22111 5364 22117
rect 5316 22108 5322 22111
rect 5534 22108 5540 22160
rect 5592 22108 5598 22160
rect 6178 22148 6184 22160
rect 5644 22120 6184 22148
rect 3050 22089 3056 22092
rect 3028 22083 3056 22089
rect 3028 22049 3040 22083
rect 3028 22043 3056 22049
rect 3050 22040 3056 22043
rect 3108 22040 3114 22092
rect 5552 22080 5580 22108
rect 5000 22052 5580 22080
rect 5000 22024 5028 22052
rect 2222 21972 2228 22024
rect 2280 22012 2286 22024
rect 3418 22012 3424 22024
rect 2280 21984 3424 22012
rect 2280 21972 2286 21984
rect 3418 21972 3424 21984
rect 3476 21972 3482 22024
rect 4982 22012 4988 22024
rect 4943 21984 4988 22012
rect 4982 21972 4988 21984
rect 5040 21972 5046 22024
rect 5644 22012 5672 22120
rect 6178 22108 6184 22120
rect 6236 22108 6242 22160
rect 6914 22148 6920 22160
rect 6748 22120 6920 22148
rect 6748 22012 6776 22120
rect 6914 22108 6920 22120
rect 6972 22108 6978 22160
rect 7926 22108 7932 22160
rect 7984 22148 7990 22160
rect 8158 22151 8216 22157
rect 8158 22148 8170 22151
rect 7984 22120 8170 22148
rect 7984 22108 7990 22120
rect 8158 22117 8170 22120
rect 8204 22117 8216 22151
rect 8158 22111 8216 22117
rect 9674 22108 9680 22160
rect 9732 22108 9738 22160
rect 9784 22148 9812 22188
rect 10870 22176 10876 22228
rect 10928 22216 10934 22228
rect 10965 22219 11023 22225
rect 10965 22216 10977 22219
rect 10928 22188 10977 22216
rect 10928 22176 10934 22188
rect 10965 22185 10977 22188
rect 11011 22216 11023 22219
rect 11011 22188 13216 22216
rect 11011 22185 11023 22188
rect 10965 22179 11023 22185
rect 9998 22151 10056 22157
rect 9998 22148 10010 22151
rect 9784 22120 10010 22148
rect 9998 22117 10010 22120
rect 10044 22117 10056 22151
rect 11606 22148 11612 22160
rect 11567 22120 11612 22148
rect 9998 22111 10056 22117
rect 11606 22108 11612 22120
rect 11664 22108 11670 22160
rect 11974 22108 11980 22160
rect 12032 22148 12038 22160
rect 13188 22157 13216 22188
rect 13173 22151 13231 22157
rect 12032 22120 12388 22148
rect 12032 22108 12038 22120
rect 6822 22040 6828 22092
rect 6880 22080 6886 22092
rect 6880 22052 6925 22080
rect 6880 22040 6886 22052
rect 8294 22040 8300 22092
rect 8352 22080 8358 22092
rect 8570 22080 8576 22092
rect 8352 22052 8576 22080
rect 8352 22040 8358 22052
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22080 8815 22083
rect 9692 22080 9720 22108
rect 8803 22052 9720 22080
rect 12360 22080 12388 22120
rect 13173 22117 13185 22151
rect 13219 22148 13231 22151
rect 13446 22148 13452 22160
rect 13219 22120 13452 22148
rect 13219 22117 13231 22120
rect 13173 22111 13231 22117
rect 13446 22108 13452 22120
rect 13504 22108 13510 22160
rect 12437 22083 12495 22089
rect 12437 22080 12449 22083
rect 12360 22052 12449 22080
rect 8803 22049 8815 22052
rect 8757 22043 8815 22049
rect 12437 22049 12449 22052
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 5270 21984 5672 22012
rect 6288 21984 6776 22012
rect 7377 22015 7435 22021
rect 4893 21947 4951 21953
rect 4893 21913 4905 21947
rect 4939 21944 4951 21947
rect 5270 21944 5298 21984
rect 4939 21916 5298 21944
rect 4939 21913 4951 21916
rect 4893 21907 4951 21913
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 6288 21953 6316 21984
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7837 22015 7895 22021
rect 7837 22012 7849 22015
rect 7423 21984 7849 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7837 21981 7849 21984
rect 7883 22012 7895 22015
rect 8110 22012 8116 22024
rect 7883 21984 8116 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 9674 22012 9680 22024
rect 9635 21984 9680 22012
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 11517 22015 11575 22021
rect 11517 21981 11529 22015
rect 11563 22012 11575 22015
rect 11974 22012 11980 22024
rect 11563 21984 11980 22012
rect 11563 21981 11575 21984
rect 11517 21975 11575 21981
rect 11974 21972 11980 21984
rect 12032 21972 12038 22024
rect 12158 22012 12164 22024
rect 12119 21984 12164 22012
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 13081 22015 13139 22021
rect 13081 21981 13093 22015
rect 13127 22012 13139 22015
rect 13814 22012 13820 22024
rect 13127 21984 13820 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 6273 21947 6331 21953
rect 6273 21944 6285 21947
rect 5684 21916 6285 21944
rect 5684 21904 5690 21916
rect 6273 21913 6285 21916
rect 6319 21913 6331 21947
rect 6273 21907 6331 21913
rect 7009 21947 7067 21953
rect 7009 21913 7021 21947
rect 7055 21944 7067 21947
rect 7558 21944 7564 21956
rect 7055 21916 7564 21944
rect 7055 21913 7067 21916
rect 7009 21907 7067 21913
rect 7558 21904 7564 21916
rect 7616 21904 7622 21956
rect 10962 21904 10968 21956
rect 11020 21944 11026 21956
rect 11333 21947 11391 21953
rect 11333 21944 11345 21947
rect 11020 21916 11345 21944
rect 11020 21904 11026 21916
rect 11333 21913 11345 21916
rect 11379 21944 11391 21947
rect 11379 21916 12388 21944
rect 11379 21913 11391 21916
rect 11333 21907 11391 21913
rect 12360 21888 12388 21916
rect 12526 21904 12532 21956
rect 12584 21944 12590 21956
rect 13633 21947 13691 21953
rect 13633 21944 13645 21947
rect 12584 21916 13645 21944
rect 12584 21904 12590 21916
rect 13633 21913 13645 21916
rect 13679 21913 13691 21947
rect 13633 21907 13691 21913
rect 4798 21836 4804 21888
rect 4856 21876 4862 21888
rect 5905 21879 5963 21885
rect 5905 21876 5917 21879
rect 4856 21848 5917 21876
rect 4856 21836 4862 21848
rect 5905 21845 5917 21848
rect 5951 21845 5963 21879
rect 5905 21839 5963 21845
rect 10597 21879 10655 21885
rect 10597 21845 10609 21879
rect 10643 21876 10655 21879
rect 11514 21876 11520 21888
rect 10643 21848 11520 21876
rect 10643 21845 10655 21848
rect 10597 21839 10655 21845
rect 11514 21836 11520 21848
rect 11572 21836 11578 21888
rect 12342 21836 12348 21888
rect 12400 21836 12406 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 4157 21675 4215 21681
rect 4157 21641 4169 21675
rect 4203 21672 4215 21675
rect 4982 21672 4988 21684
rect 4203 21644 4988 21672
rect 4203 21641 4215 21644
rect 4157 21635 4215 21641
rect 4982 21632 4988 21644
rect 5040 21632 5046 21684
rect 5258 21632 5264 21684
rect 5316 21672 5322 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5316 21644 5641 21672
rect 5316 21632 5322 21644
rect 5629 21641 5641 21644
rect 5675 21672 5687 21675
rect 7745 21675 7803 21681
rect 7745 21672 7757 21675
rect 5675 21644 7757 21672
rect 5675 21641 5687 21644
rect 5629 21635 5687 21641
rect 7745 21641 7757 21644
rect 7791 21672 7803 21675
rect 7926 21672 7932 21684
rect 7791 21644 7932 21672
rect 7791 21641 7803 21644
rect 7745 21635 7803 21641
rect 7926 21632 7932 21644
rect 7984 21672 7990 21684
rect 8754 21672 8760 21684
rect 7984 21644 8760 21672
rect 7984 21632 7990 21644
rect 8754 21632 8760 21644
rect 8812 21672 8818 21684
rect 9033 21675 9091 21681
rect 9033 21672 9045 21675
rect 8812 21644 9045 21672
rect 8812 21632 8818 21644
rect 9033 21641 9045 21644
rect 9079 21672 9091 21675
rect 9401 21675 9459 21681
rect 9401 21672 9413 21675
rect 9079 21644 9413 21672
rect 9079 21641 9091 21644
rect 9033 21635 9091 21641
rect 9401 21641 9413 21644
rect 9447 21641 9459 21675
rect 9401 21635 9459 21641
rect 10505 21675 10563 21681
rect 10505 21641 10517 21675
rect 10551 21672 10563 21675
rect 11241 21675 11299 21681
rect 11241 21672 11253 21675
rect 10551 21644 11253 21672
rect 10551 21641 10563 21644
rect 10505 21635 10563 21641
rect 11241 21641 11253 21644
rect 11287 21672 11299 21675
rect 11606 21672 11612 21684
rect 11287 21644 11612 21672
rect 11287 21641 11299 21644
rect 11241 21635 11299 21641
rect 3418 21564 3424 21616
rect 3476 21604 3482 21616
rect 3476 21576 6776 21604
rect 3476 21564 3482 21576
rect 3789 21539 3847 21545
rect 3789 21505 3801 21539
rect 3835 21536 3847 21539
rect 4706 21536 4712 21548
rect 3835 21508 4712 21536
rect 3835 21505 3847 21508
rect 3789 21499 3847 21505
rect 4706 21496 4712 21508
rect 4764 21496 4770 21548
rect 4982 21536 4988 21548
rect 4943 21508 4988 21536
rect 4982 21496 4988 21508
rect 5040 21496 5046 21548
rect 6748 21468 6776 21576
rect 6952 21471 7010 21477
rect 6952 21468 6964 21471
rect 6748 21440 6964 21468
rect 6952 21437 6964 21440
rect 6998 21468 7010 21471
rect 7377 21471 7435 21477
rect 7377 21468 7389 21471
rect 6998 21440 7389 21468
rect 6998 21437 7010 21440
rect 6952 21431 7010 21437
rect 7377 21437 7389 21440
rect 7423 21437 7435 21471
rect 7377 21431 7435 21437
rect 7650 21428 7656 21480
rect 7708 21468 7714 21480
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7708 21440 7941 21468
rect 7708 21428 7714 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 8386 21468 8392 21480
rect 8347 21440 8392 21468
rect 7929 21431 7987 21437
rect 8386 21428 8392 21440
rect 8444 21428 8450 21480
rect 4525 21403 4583 21409
rect 4525 21369 4537 21403
rect 4571 21400 4583 21403
rect 4798 21400 4804 21412
rect 4571 21372 4804 21400
rect 4571 21369 4583 21372
rect 4525 21363 4583 21369
rect 4798 21360 4804 21372
rect 4856 21360 4862 21412
rect 8662 21400 8668 21412
rect 8623 21372 8668 21400
rect 8662 21360 8668 21372
rect 8720 21360 8726 21412
rect 9416 21400 9444 21635
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 12161 21675 12219 21681
rect 12161 21672 12173 21675
rect 12032 21644 12173 21672
rect 12032 21632 12038 21644
rect 12161 21641 12173 21644
rect 12207 21641 12219 21675
rect 13446 21672 13452 21684
rect 13407 21644 13452 21672
rect 12161 21635 12219 21641
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 13814 21672 13820 21684
rect 13775 21644 13820 21672
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 9674 21564 9680 21616
rect 9732 21604 9738 21616
rect 10781 21607 10839 21613
rect 10781 21604 10793 21607
rect 9732 21576 10793 21604
rect 9732 21564 9738 21576
rect 10781 21573 10793 21576
rect 10827 21573 10839 21607
rect 10781 21567 10839 21573
rect 11471 21607 11529 21613
rect 11471 21573 11483 21607
rect 11517 21604 11529 21607
rect 13832 21604 13860 21632
rect 11517 21576 13860 21604
rect 11517 21573 11529 21576
rect 11471 21567 11529 21573
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 12805 21539 12863 21545
rect 12805 21536 12817 21539
rect 12216 21508 12817 21536
rect 12216 21496 12222 21508
rect 12805 21505 12817 21508
rect 12851 21505 12863 21539
rect 12805 21499 12863 21505
rect 9582 21468 9588 21480
rect 9543 21440 9588 21468
rect 9582 21428 9588 21440
rect 9640 21428 9646 21480
rect 10778 21428 10784 21480
rect 10836 21468 10842 21480
rect 11330 21468 11336 21480
rect 10836 21440 11336 21468
rect 10836 21428 10842 21440
rect 11330 21428 11336 21440
rect 11388 21477 11394 21480
rect 11388 21471 11437 21477
rect 11388 21437 11391 21471
rect 11425 21468 11437 21471
rect 11793 21471 11851 21477
rect 11793 21468 11805 21471
rect 11425 21440 11805 21468
rect 11425 21437 11437 21440
rect 11388 21431 11437 21437
rect 11793 21437 11805 21440
rect 11839 21437 11851 21471
rect 11793 21431 11851 21437
rect 11388 21428 11394 21431
rect 9950 21409 9956 21412
rect 9906 21403 9956 21409
rect 9906 21400 9918 21403
rect 9416 21372 9918 21400
rect 9906 21369 9918 21372
rect 9952 21369 9956 21403
rect 9906 21363 9956 21369
rect 9950 21360 9956 21363
rect 10008 21400 10014 21412
rect 12526 21400 12532 21412
rect 10008 21372 10054 21400
rect 12487 21372 12532 21400
rect 10008 21360 10014 21372
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 12618 21360 12624 21412
rect 12676 21400 12682 21412
rect 12676 21372 12721 21400
rect 12676 21360 12682 21372
rect 3050 21332 3056 21344
rect 3011 21304 3056 21332
rect 3050 21292 3056 21304
rect 3108 21292 3114 21344
rect 3510 21292 3516 21344
rect 3568 21332 3574 21344
rect 5902 21332 5908 21344
rect 3568 21304 5908 21332
rect 3568 21292 3574 21304
rect 5902 21292 5908 21304
rect 5960 21332 5966 21344
rect 6549 21335 6607 21341
rect 6549 21332 6561 21335
rect 5960 21304 6561 21332
rect 5960 21292 5966 21304
rect 6549 21301 6561 21304
rect 6595 21332 6607 21335
rect 6822 21332 6828 21344
rect 6595 21304 6828 21332
rect 6595 21301 6607 21304
rect 6549 21295 6607 21301
rect 6822 21292 6828 21304
rect 6880 21292 6886 21344
rect 7055 21335 7113 21341
rect 7055 21301 7067 21335
rect 7101 21332 7113 21335
rect 7282 21332 7288 21344
rect 7101 21304 7288 21332
rect 7101 21301 7113 21304
rect 7055 21295 7113 21301
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 7650 21088 7656 21140
rect 7708 21128 7714 21140
rect 7837 21131 7895 21137
rect 7837 21128 7849 21131
rect 7708 21100 7849 21128
rect 7708 21088 7714 21100
rect 7837 21097 7849 21100
rect 7883 21097 7895 21131
rect 8110 21128 8116 21140
rect 8071 21100 8116 21128
rect 7837 21091 7895 21097
rect 8110 21088 8116 21100
rect 8168 21088 8174 21140
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 9033 21131 9091 21137
rect 9033 21128 9045 21131
rect 8720 21100 9045 21128
rect 8720 21088 8726 21100
rect 9033 21097 9045 21100
rect 9079 21097 9091 21131
rect 9033 21091 9091 21097
rect 10597 21131 10655 21137
rect 10597 21097 10609 21131
rect 10643 21128 10655 21131
rect 12529 21131 12587 21137
rect 12529 21128 12541 21131
rect 10643 21100 12541 21128
rect 10643 21097 10655 21100
rect 10597 21091 10655 21097
rect 12529 21097 12541 21100
rect 12575 21128 12587 21131
rect 12618 21128 12624 21140
rect 12575 21100 12624 21128
rect 12575 21097 12587 21100
rect 12529 21091 12587 21097
rect 12618 21088 12624 21100
rect 12676 21088 12682 21140
rect 13170 21137 13176 21140
rect 13127 21131 13176 21137
rect 13127 21097 13139 21131
rect 13173 21097 13176 21131
rect 13127 21091 13176 21097
rect 13170 21088 13176 21091
rect 13228 21088 13234 21140
rect 7190 21060 7196 21072
rect 7151 21032 7196 21060
rect 7190 21020 7196 21032
rect 7248 21020 7254 21072
rect 7374 21020 7380 21072
rect 7432 21060 7438 21072
rect 7432 21032 8064 21060
rect 7432 21020 7438 21032
rect 4798 20992 4804 21004
rect 4759 20964 4804 20992
rect 4798 20952 4804 20964
rect 4856 20952 4862 21004
rect 6086 20952 6092 21004
rect 6144 20992 6150 21004
rect 6362 20992 6368 21004
rect 6144 20964 6368 20992
rect 6144 20952 6150 20964
rect 6362 20952 6368 20964
rect 6420 20992 6426 21004
rect 8036 21001 8064 21032
rect 9950 21020 9956 21072
rect 10008 21069 10014 21072
rect 10008 21063 10056 21069
rect 10008 21029 10010 21063
rect 10044 21029 10056 21063
rect 10008 21023 10056 21029
rect 10008 21020 10014 21023
rect 11514 21020 11520 21072
rect 11572 21060 11578 21072
rect 11609 21063 11667 21069
rect 11609 21060 11621 21063
rect 11572 21032 11621 21060
rect 11572 21020 11578 21032
rect 11609 21029 11621 21032
rect 11655 21029 11667 21063
rect 11609 21023 11667 21029
rect 6457 20995 6515 21001
rect 6457 20992 6469 20995
rect 6420 20964 6469 20992
rect 6420 20952 6426 20964
rect 6457 20961 6469 20964
rect 6503 20961 6515 20995
rect 6457 20955 6515 20961
rect 7009 20995 7067 21001
rect 7009 20961 7021 20995
rect 7055 20961 7067 20995
rect 7009 20955 7067 20961
rect 8021 20995 8079 21001
rect 8021 20961 8033 20995
rect 8067 20992 8079 20995
rect 8202 20992 8208 21004
rect 8067 20964 8208 20992
rect 8067 20961 8079 20964
rect 8021 20955 8079 20961
rect 4430 20924 4436 20936
rect 4391 20896 4436 20924
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 6546 20884 6552 20936
rect 6604 20924 6610 20936
rect 7024 20924 7052 20955
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 13078 21001 13084 21004
rect 8481 20995 8539 21001
rect 8481 20961 8493 20995
rect 8527 20961 8539 20995
rect 8481 20955 8539 20961
rect 13056 20995 13084 21001
rect 13056 20961 13068 20995
rect 13056 20955 13084 20961
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 6604 20896 7573 20924
rect 6604 20884 6610 20896
rect 7561 20893 7573 20896
rect 7607 20924 7619 20927
rect 8386 20924 8392 20936
rect 7607 20896 8392 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 8386 20884 8392 20896
rect 8444 20924 8450 20936
rect 8496 20924 8524 20955
rect 13078 20952 13084 20955
rect 13136 20952 13142 21004
rect 9674 20924 9680 20936
rect 8444 20896 8524 20924
rect 9635 20896 9680 20924
rect 8444 20884 8450 20896
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11204 20896 11529 20924
rect 11204 20884 11210 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 12158 20924 12164 20936
rect 12119 20896 12164 20924
rect 11517 20887 11575 20893
rect 12158 20884 12164 20896
rect 12216 20924 12222 20936
rect 12216 20896 12480 20924
rect 12216 20884 12222 20896
rect 12452 20856 12480 20896
rect 12526 20884 12532 20936
rect 12584 20924 12590 20936
rect 12805 20927 12863 20933
rect 12805 20924 12817 20927
rect 12584 20896 12817 20924
rect 12584 20884 12590 20896
rect 12805 20893 12817 20896
rect 12851 20893 12863 20927
rect 12805 20887 12863 20893
rect 13078 20856 13084 20868
rect 12452 20828 13084 20856
rect 13078 20816 13084 20828
rect 13136 20816 13142 20868
rect 9493 20791 9551 20797
rect 9493 20757 9505 20791
rect 9539 20788 9551 20791
rect 9582 20788 9588 20800
rect 9539 20760 9588 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 10962 20788 10968 20800
rect 10923 20760 10968 20788
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 4249 20587 4307 20593
rect 4249 20553 4261 20587
rect 4295 20584 4307 20587
rect 4430 20584 4436 20596
rect 4295 20556 4436 20584
rect 4295 20553 4307 20556
rect 4249 20547 4307 20553
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4798 20544 4804 20596
rect 4856 20584 4862 20596
rect 5353 20587 5411 20593
rect 5353 20584 5365 20587
rect 4856 20556 5365 20584
rect 4856 20544 4862 20556
rect 5353 20553 5365 20556
rect 5399 20553 5411 20587
rect 6546 20584 6552 20596
rect 6507 20556 6552 20584
rect 5353 20547 5411 20553
rect 6546 20544 6552 20556
rect 6604 20584 6610 20596
rect 7193 20587 7251 20593
rect 7193 20584 7205 20587
rect 6604 20556 7205 20584
rect 6604 20544 6610 20556
rect 7193 20553 7205 20556
rect 7239 20553 7251 20587
rect 7193 20547 7251 20553
rect 4982 20516 4988 20528
rect 4943 20488 4988 20516
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 7208 20448 7236 20547
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8389 20587 8447 20593
rect 8389 20584 8401 20587
rect 8352 20556 8401 20584
rect 8352 20544 8358 20556
rect 8389 20553 8401 20556
rect 8435 20553 8447 20587
rect 8754 20584 8760 20596
rect 8715 20556 8760 20584
rect 8389 20547 8447 20553
rect 8754 20544 8760 20556
rect 8812 20584 8818 20596
rect 9306 20584 9312 20596
rect 8812 20556 9312 20584
rect 8812 20544 8818 20556
rect 9306 20544 9312 20556
rect 9364 20584 9370 20596
rect 10137 20587 10195 20593
rect 10137 20584 10149 20587
rect 9364 20556 10149 20584
rect 9364 20544 9370 20556
rect 10137 20553 10149 20556
rect 10183 20553 10195 20587
rect 10137 20547 10195 20553
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11701 20587 11759 20593
rect 11701 20584 11713 20587
rect 11572 20556 11713 20584
rect 11572 20544 11578 20556
rect 11701 20553 11713 20556
rect 11747 20553 11759 20587
rect 11701 20547 11759 20553
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 12575 20587 12633 20593
rect 12575 20584 12587 20587
rect 12492 20556 12587 20584
rect 12492 20544 12498 20556
rect 12575 20553 12587 20556
rect 12621 20553 12633 20587
rect 12575 20547 12633 20553
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 13136 20556 13277 20584
rect 13136 20544 13142 20556
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13265 20547 13323 20553
rect 10962 20516 10968 20528
rect 10796 20488 10968 20516
rect 7208 20420 7880 20448
rect 7852 20389 7880 20420
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 10796 20457 10824 20488
rect 10962 20476 10968 20488
rect 11020 20516 11026 20528
rect 13587 20519 13645 20525
rect 13587 20516 13599 20519
rect 11020 20488 13599 20516
rect 11020 20476 11026 20488
rect 13587 20485 13599 20488
rect 13633 20485 13645 20519
rect 13587 20479 13645 20485
rect 8941 20451 8999 20457
rect 8941 20448 8953 20451
rect 8720 20420 8953 20448
rect 8720 20408 8726 20420
rect 8941 20417 8953 20420
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20417 10839 20451
rect 11146 20448 11152 20460
rect 11107 20420 11152 20448
rect 10781 20411 10839 20417
rect 11146 20408 11152 20420
rect 11204 20448 11210 20460
rect 12069 20451 12127 20457
rect 12069 20448 12081 20451
rect 11204 20420 12081 20448
rect 11204 20408 11210 20420
rect 12069 20417 12081 20420
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 5813 20383 5871 20389
rect 5813 20349 5825 20383
rect 5859 20380 5871 20383
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 5859 20352 7665 20380
rect 5859 20349 5871 20352
rect 5813 20343 5871 20349
rect 7653 20349 7665 20352
rect 7699 20349 7711 20383
rect 7653 20343 7711 20349
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 9674 20380 9680 20392
rect 8159 20352 9680 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 3329 20315 3387 20321
rect 3329 20281 3341 20315
rect 3375 20312 3387 20315
rect 3881 20315 3939 20321
rect 3881 20312 3893 20315
rect 3375 20284 3893 20312
rect 3375 20281 3387 20284
rect 3329 20275 3387 20281
rect 3881 20281 3893 20284
rect 3927 20312 3939 20315
rect 4433 20315 4491 20321
rect 4433 20312 4445 20315
rect 3927 20284 4445 20312
rect 3927 20281 3939 20284
rect 3881 20275 3939 20281
rect 4433 20281 4445 20284
rect 4479 20281 4491 20315
rect 4433 20275 4491 20281
rect 4522 20272 4528 20324
rect 4580 20312 4586 20324
rect 4580 20284 4625 20312
rect 4580 20272 4586 20284
rect 5534 20272 5540 20324
rect 5592 20312 5598 20324
rect 6089 20315 6147 20321
rect 6089 20312 6101 20315
rect 5592 20284 6101 20312
rect 5592 20272 5598 20284
rect 6089 20281 6101 20284
rect 6135 20312 6147 20315
rect 6362 20312 6368 20324
rect 6135 20284 6368 20312
rect 6135 20281 6147 20284
rect 6089 20275 6147 20281
rect 6362 20272 6368 20284
rect 6420 20272 6426 20324
rect 7668 20312 7696 20343
rect 9674 20340 9680 20352
rect 9732 20340 9738 20392
rect 12526 20389 12532 20392
rect 12488 20383 12532 20389
rect 12488 20349 12500 20383
rect 12584 20380 12590 20392
rect 12897 20383 12955 20389
rect 12897 20380 12909 20383
rect 12584 20352 12909 20380
rect 12488 20343 12532 20349
rect 12526 20340 12532 20343
rect 12584 20340 12590 20352
rect 12897 20349 12909 20352
rect 12943 20349 12955 20383
rect 12897 20343 12955 20349
rect 13446 20340 13452 20392
rect 13504 20389 13510 20392
rect 13504 20383 13542 20389
rect 13530 20380 13542 20383
rect 13906 20380 13912 20392
rect 13530 20352 13912 20380
rect 13530 20349 13542 20352
rect 13504 20343 13542 20349
rect 13504 20340 13510 20343
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 7742 20312 7748 20324
rect 7655 20284 7748 20312
rect 7742 20272 7748 20284
rect 7800 20312 7806 20324
rect 8202 20312 8208 20324
rect 7800 20284 8208 20312
rect 7800 20272 7806 20284
rect 8202 20272 8208 20284
rect 8260 20272 8266 20324
rect 9306 20321 9312 20324
rect 9303 20312 9312 20321
rect 9267 20284 9312 20312
rect 9303 20275 9312 20284
rect 9306 20272 9312 20275
rect 9364 20272 9370 20324
rect 10597 20315 10655 20321
rect 10597 20312 10609 20315
rect 9876 20284 10609 20312
rect 9876 20253 9904 20284
rect 10597 20281 10609 20284
rect 10643 20312 10655 20315
rect 10873 20315 10931 20321
rect 10873 20312 10885 20315
rect 10643 20284 10885 20312
rect 10643 20281 10655 20284
rect 10597 20275 10655 20281
rect 10873 20281 10885 20284
rect 10919 20312 10931 20315
rect 10962 20312 10968 20324
rect 10919 20284 10968 20312
rect 10919 20281 10931 20284
rect 10873 20275 10931 20281
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 9861 20247 9919 20253
rect 9861 20213 9873 20247
rect 9907 20213 9919 20247
rect 9861 20207 9919 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 3099 20043 3157 20049
rect 3099 20040 3111 20043
rect 2924 20012 3111 20040
rect 2924 20000 2930 20012
rect 3099 20009 3111 20012
rect 3145 20009 3157 20043
rect 3099 20003 3157 20009
rect 6178 20000 6184 20052
rect 6236 20040 6242 20052
rect 6822 20040 6828 20052
rect 6236 20012 6828 20040
rect 6236 20000 6242 20012
rect 6822 20000 6828 20012
rect 6880 20040 6886 20052
rect 6917 20043 6975 20049
rect 6917 20040 6929 20043
rect 6880 20012 6929 20040
rect 6880 20000 6886 20012
rect 6917 20009 6929 20012
rect 6963 20040 6975 20043
rect 7193 20043 7251 20049
rect 7193 20040 7205 20043
rect 6963 20012 7205 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7193 20009 7205 20012
rect 7239 20009 7251 20043
rect 7193 20003 7251 20009
rect 9493 20043 9551 20049
rect 9493 20009 9505 20043
rect 9539 20040 9551 20043
rect 9674 20040 9680 20052
rect 9539 20012 9680 20040
rect 9539 20009 9551 20012
rect 9493 20003 9551 20009
rect 4982 19972 4988 19984
rect 3988 19944 4988 19972
rect 3028 19907 3086 19913
rect 3028 19873 3040 19907
rect 3074 19904 3086 19907
rect 3142 19904 3148 19916
rect 3074 19876 3148 19904
rect 3074 19873 3086 19876
rect 3028 19867 3086 19873
rect 3142 19864 3148 19876
rect 3200 19904 3206 19916
rect 3988 19904 4016 19944
rect 4982 19932 4988 19944
rect 5040 19932 5046 19984
rect 4890 19904 4896 19916
rect 3200 19876 4016 19904
rect 4851 19876 4896 19904
rect 3200 19864 3206 19876
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 6457 19907 6515 19913
rect 6457 19873 6469 19907
rect 6503 19873 6515 19907
rect 7208 19904 7236 20003
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10962 20000 10968 20052
rect 11020 20000 11026 20052
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 11974 20040 11980 20052
rect 11931 20012 11980 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 10226 19932 10232 19984
rect 10284 19972 10290 19984
rect 10413 19975 10471 19981
rect 10413 19972 10425 19975
rect 10284 19944 10425 19972
rect 10284 19932 10290 19944
rect 10413 19941 10425 19944
rect 10459 19941 10471 19975
rect 10413 19935 10471 19941
rect 10505 19975 10563 19981
rect 10505 19941 10517 19975
rect 10551 19972 10563 19975
rect 10980 19972 11008 20000
rect 10551 19944 11008 19972
rect 10551 19941 10563 19944
rect 10505 19935 10563 19941
rect 11422 19932 11428 19984
rect 11480 19972 11486 19984
rect 12066 19972 12072 19984
rect 11480 19944 12072 19972
rect 11480 19932 11486 19944
rect 12066 19932 12072 19944
rect 12124 19932 12130 19984
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 7208 19876 7389 19904
rect 6457 19867 6515 19873
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7650 19904 7656 19916
rect 7611 19876 7656 19904
rect 7377 19867 7435 19873
rect 4982 19836 4988 19848
rect 4943 19808 4988 19836
rect 4982 19796 4988 19808
rect 5040 19796 5046 19848
rect 6270 19796 6276 19848
rect 6328 19836 6334 19848
rect 6472 19836 6500 19867
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 8386 19864 8392 19916
rect 8444 19904 8450 19916
rect 9953 19907 10011 19913
rect 9953 19904 9965 19907
rect 8444 19876 9965 19904
rect 8444 19864 8450 19876
rect 9953 19873 9965 19876
rect 9999 19904 10011 19907
rect 10042 19904 10048 19916
rect 9999 19876 10048 19904
rect 9999 19873 10011 19876
rect 9953 19867 10011 19873
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 7006 19836 7012 19848
rect 6328 19808 7012 19836
rect 6328 19796 6334 19808
rect 7006 19796 7012 19808
rect 7064 19836 7070 19848
rect 7469 19839 7527 19845
rect 7469 19836 7481 19839
rect 7064 19808 7481 19836
rect 7064 19796 7070 19808
rect 7469 19805 7481 19808
rect 7515 19805 7527 19839
rect 7834 19836 7840 19848
rect 7795 19808 7840 19836
rect 7469 19799 7527 19805
rect 7484 19768 7512 19799
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 10870 19836 10876 19848
rect 10831 19808 10876 19836
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 8389 19771 8447 19777
rect 8389 19768 8401 19771
rect 7484 19740 8401 19768
rect 8389 19737 8401 19740
rect 8435 19768 8447 19771
rect 8478 19768 8484 19780
rect 8435 19740 8484 19768
rect 8435 19737 8447 19740
rect 8389 19731 8447 19737
rect 8478 19728 8484 19740
rect 8536 19728 8542 19780
rect 5258 19700 5264 19712
rect 5219 19672 5264 19700
rect 5258 19660 5264 19672
rect 5316 19700 5322 19712
rect 6086 19700 6092 19712
rect 5316 19672 6092 19700
rect 5316 19660 5322 19672
rect 6086 19660 6092 19672
rect 6144 19660 6150 19712
rect 8754 19700 8760 19712
rect 8715 19672 8760 19700
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 3053 19499 3111 19505
rect 3053 19465 3065 19499
rect 3099 19496 3111 19499
rect 3142 19496 3148 19508
rect 3099 19468 3148 19496
rect 3099 19465 3111 19468
rect 3053 19459 3111 19465
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 6270 19496 6276 19508
rect 6231 19468 6276 19496
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 10962 19496 10968 19508
rect 10923 19468 10968 19496
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 5258 19428 5264 19440
rect 5219 19400 5264 19428
rect 5258 19388 5264 19400
rect 5316 19388 5322 19440
rect 8478 19428 8484 19440
rect 8439 19400 8484 19428
rect 8478 19388 8484 19400
rect 8536 19388 8542 19440
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19360 4123 19363
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4111 19332 4721 19360
rect 4111 19329 4123 19332
rect 4065 19323 4123 19329
rect 4709 19329 4721 19332
rect 4755 19360 4767 19363
rect 4890 19360 4896 19372
rect 4755 19332 4896 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 4890 19320 4896 19332
rect 4948 19360 4954 19372
rect 4948 19332 5488 19360
rect 4948 19320 4954 19332
rect 3697 19295 3755 19301
rect 3697 19261 3709 19295
rect 3743 19292 3755 19295
rect 4154 19292 4160 19304
rect 3743 19264 4160 19292
rect 3743 19261 3755 19264
rect 3697 19255 3755 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5169 19295 5227 19301
rect 5169 19292 5181 19295
rect 5123 19264 5181 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5169 19261 5181 19264
rect 5215 19292 5227 19295
rect 5258 19292 5264 19304
rect 5215 19264 5264 19292
rect 5215 19261 5227 19264
rect 5169 19255 5227 19261
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 5460 19301 5488 19332
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 6917 19363 6975 19369
rect 6917 19360 6929 19363
rect 6144 19332 6929 19360
rect 6144 19320 6150 19332
rect 6917 19329 6929 19332
rect 6963 19329 6975 19363
rect 6917 19323 6975 19329
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7926 19360 7932 19372
rect 7524 19332 7932 19360
rect 7524 19320 7530 19332
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 5445 19295 5503 19301
rect 5445 19292 5457 19295
rect 5355 19264 5457 19292
rect 5445 19261 5457 19264
rect 5491 19261 5503 19295
rect 5445 19255 5503 19261
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19261 6883 19295
rect 7101 19295 7159 19301
rect 7101 19292 7113 19295
rect 6825 19255 6883 19261
rect 6932 19264 7113 19292
rect 5460 19168 5488 19255
rect 6840 19168 6868 19255
rect 6932 19236 6960 19264
rect 7101 19261 7113 19264
rect 7147 19292 7159 19295
rect 7650 19292 7656 19304
rect 7147 19264 7656 19292
rect 7147 19261 7159 19264
rect 7101 19255 7159 19261
rect 7650 19252 7656 19264
rect 7708 19292 7714 19304
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 7708 19264 7849 19292
rect 7708 19252 7714 19264
rect 7837 19261 7849 19264
rect 7883 19261 7895 19295
rect 7837 19255 7895 19261
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8343 19264 8401 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 8665 19295 8723 19301
rect 8665 19261 8677 19295
rect 8711 19292 8723 19295
rect 8754 19292 8760 19304
rect 8711 19264 8760 19292
rect 8711 19261 8723 19264
rect 8665 19255 8723 19261
rect 6914 19184 6920 19236
rect 6972 19184 6978 19236
rect 7558 19224 7564 19236
rect 7519 19196 7564 19224
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 7926 19184 7932 19236
rect 7984 19224 7990 19236
rect 8312 19224 8340 19255
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 9824 19264 9965 19292
rect 9824 19252 9830 19264
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 10042 19252 10048 19304
rect 10100 19292 10106 19304
rect 10413 19295 10471 19301
rect 10413 19292 10425 19295
rect 10100 19264 10425 19292
rect 10100 19252 10106 19264
rect 10413 19261 10425 19264
rect 10459 19261 10471 19295
rect 10413 19255 10471 19261
rect 7984 19196 8340 19224
rect 7984 19184 7990 19196
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 9640 19196 10088 19224
rect 9640 19184 9646 19196
rect 4338 19156 4344 19168
rect 4299 19128 4344 19156
rect 4338 19116 4344 19128
rect 4396 19116 4402 19168
rect 5442 19116 5448 19168
rect 5500 19116 5506 19168
rect 5626 19156 5632 19168
rect 5587 19128 5632 19156
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 6178 19116 6184 19168
rect 6236 19156 6242 19168
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6236 19128 6561 19156
rect 6236 19116 6242 19128
rect 6549 19125 6561 19128
rect 6595 19156 6607 19159
rect 6638 19156 6644 19168
rect 6595 19128 6644 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 6638 19116 6644 19128
rect 6696 19116 6702 19168
rect 6822 19116 6828 19168
rect 6880 19116 6886 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 8849 19159 8907 19165
rect 8849 19156 8861 19159
rect 8352 19128 8861 19156
rect 8352 19116 8358 19128
rect 8849 19125 8861 19128
rect 8895 19125 8907 19159
rect 9766 19156 9772 19168
rect 9727 19128 9772 19156
rect 8849 19119 8907 19125
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10060 19165 10088 19196
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19125 10103 19159
rect 10045 19119 10103 19125
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 4154 18912 4160 18964
rect 4212 18952 4218 18964
rect 5169 18955 5227 18961
rect 5169 18952 5181 18955
rect 4212 18924 5181 18952
rect 4212 18912 4218 18924
rect 5169 18921 5181 18924
rect 5215 18921 5227 18955
rect 6086 18952 6092 18964
rect 6047 18924 6092 18952
rect 5169 18915 5227 18921
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7377 18955 7435 18961
rect 7377 18952 7389 18955
rect 7064 18924 7389 18952
rect 7064 18912 7070 18924
rect 7377 18921 7389 18924
rect 7423 18921 7435 18955
rect 7377 18915 7435 18921
rect 10226 18912 10232 18964
rect 10284 18952 10290 18964
rect 10321 18955 10379 18961
rect 10321 18952 10333 18955
rect 10284 18924 10333 18952
rect 10284 18912 10290 18924
rect 10321 18921 10333 18924
rect 10367 18921 10379 18955
rect 10321 18915 10379 18921
rect 4617 18887 4675 18893
rect 4617 18853 4629 18887
rect 4663 18884 4675 18887
rect 6822 18884 6828 18896
rect 4663 18856 6828 18884
rect 4663 18853 4675 18856
rect 4617 18847 4675 18853
rect 4724 18825 4752 18856
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 8754 18844 8760 18896
rect 8812 18844 8818 18896
rect 4709 18819 4767 18825
rect 4709 18785 4721 18819
rect 4755 18816 4767 18819
rect 4982 18816 4988 18828
rect 4755 18788 4789 18816
rect 4943 18788 4988 18816
rect 4755 18785 4767 18788
rect 4709 18779 4767 18785
rect 4982 18776 4988 18788
rect 5040 18776 5046 18828
rect 5258 18776 5264 18828
rect 5316 18816 5322 18828
rect 5810 18816 5816 18828
rect 5316 18788 5816 18816
rect 5316 18776 5322 18788
rect 5810 18776 5816 18788
rect 5868 18816 5874 18828
rect 6270 18816 6276 18828
rect 5868 18788 6276 18816
rect 5868 18776 5874 18788
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18816 6607 18819
rect 6914 18816 6920 18828
rect 6595 18788 6920 18816
rect 6595 18785 6607 18788
rect 6549 18779 6607 18785
rect 5442 18708 5448 18760
rect 5500 18748 5506 18760
rect 6178 18748 6184 18760
rect 5500 18720 6184 18748
rect 5500 18708 5506 18720
rect 6178 18708 6184 18720
rect 6236 18748 6242 18760
rect 6564 18748 6592 18779
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 8202 18816 8208 18828
rect 8163 18788 8208 18816
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 8772 18816 8800 18844
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 8619 18788 8708 18816
rect 8772 18788 9689 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 6236 18720 6592 18748
rect 6236 18708 6242 18720
rect 6638 18708 6644 18760
rect 6696 18748 6702 18760
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6696 18720 6745 18748
rect 6696 18708 6702 18720
rect 6733 18717 6745 18720
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 4798 18680 4804 18692
rect 4711 18652 4804 18680
rect 4798 18640 4804 18652
rect 4856 18680 4862 18692
rect 6365 18683 6423 18689
rect 6365 18680 6377 18683
rect 4856 18652 6377 18680
rect 4856 18640 4862 18652
rect 6365 18649 6377 18652
rect 6411 18680 6423 18683
rect 6822 18680 6828 18692
rect 6411 18652 6828 18680
rect 6411 18649 6423 18652
rect 6365 18643 6423 18649
rect 6822 18640 6828 18652
rect 6880 18680 6886 18692
rect 7006 18680 7012 18692
rect 6880 18652 7012 18680
rect 6880 18640 6886 18652
rect 7006 18640 7012 18652
rect 7064 18640 7070 18692
rect 7929 18683 7987 18689
rect 7929 18649 7941 18683
rect 7975 18680 7987 18683
rect 8386 18680 8392 18692
rect 7975 18652 8392 18680
rect 7975 18649 7987 18652
rect 7929 18643 7987 18649
rect 8386 18640 8392 18652
rect 8444 18680 8450 18692
rect 8680 18680 8708 18788
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 10686 18816 10692 18828
rect 10647 18788 10692 18816
rect 9677 18779 9735 18785
rect 10686 18776 10692 18788
rect 10744 18776 10750 18828
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18748 8815 18751
rect 9582 18748 9588 18760
rect 8803 18720 9588 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 11514 18708 11520 18760
rect 11572 18748 11578 18760
rect 11701 18751 11759 18757
rect 11701 18748 11713 18751
rect 11572 18720 11713 18748
rect 11572 18708 11578 18720
rect 11701 18717 11713 18720
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 9861 18683 9919 18689
rect 9861 18680 9873 18683
rect 8444 18652 9873 18680
rect 8444 18640 8450 18652
rect 9861 18649 9873 18652
rect 9907 18649 9919 18683
rect 9861 18643 9919 18649
rect 5810 18612 5816 18624
rect 5771 18584 5816 18612
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 10870 18612 10876 18624
rect 10831 18584 10876 18612
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 2866 18408 2872 18420
rect 2827 18380 2872 18408
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3881 18411 3939 18417
rect 3881 18377 3893 18411
rect 3927 18408 3939 18411
rect 4982 18408 4988 18420
rect 3927 18380 4988 18408
rect 3927 18377 3939 18380
rect 3881 18371 3939 18377
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 6328 18380 6377 18408
rect 6328 18368 6334 18380
rect 6365 18377 6377 18380
rect 6411 18408 6423 18411
rect 7926 18408 7932 18420
rect 6411 18380 7932 18408
rect 6411 18377 6423 18380
rect 6365 18371 6423 18377
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 8754 18368 8760 18420
rect 8812 18408 8818 18420
rect 8849 18411 8907 18417
rect 8849 18408 8861 18411
rect 8812 18380 8861 18408
rect 8812 18368 8818 18380
rect 8849 18377 8861 18380
rect 8895 18377 8907 18411
rect 9306 18408 9312 18420
rect 9267 18380 9312 18408
rect 8849 18371 8907 18377
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 10686 18408 10692 18420
rect 10647 18380 10692 18408
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 3145 18343 3203 18349
rect 3145 18309 3157 18343
rect 3191 18340 3203 18343
rect 4062 18340 4068 18352
rect 3191 18312 4068 18340
rect 3191 18309 3203 18312
rect 3145 18303 3203 18309
rect 4062 18300 4068 18312
rect 4120 18300 4126 18352
rect 4798 18340 4804 18352
rect 4759 18312 4804 18340
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 5810 18300 5816 18352
rect 5868 18340 5874 18352
rect 7009 18343 7067 18349
rect 7009 18340 7021 18343
rect 5868 18312 7021 18340
rect 5868 18300 5874 18312
rect 7009 18309 7021 18312
rect 7055 18340 7067 18343
rect 7055 18312 7788 18340
rect 7055 18309 7067 18312
rect 7009 18303 7067 18309
rect 5828 18272 5856 18300
rect 5276 18244 5856 18272
rect 2866 18164 2872 18216
rect 2924 18204 2930 18216
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2924 18176 2973 18204
rect 2924 18164 2930 18176
rect 2961 18173 2973 18176
rect 3007 18173 3019 18207
rect 2961 18167 3019 18173
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3970 18204 3976 18216
rect 3559 18176 3976 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 5276 18213 5304 18244
rect 5261 18207 5319 18213
rect 5261 18173 5273 18207
rect 5307 18173 5319 18207
rect 5442 18204 5448 18216
rect 5403 18176 5448 18204
rect 5261 18167 5319 18173
rect 5442 18164 5448 18176
rect 5500 18164 5506 18216
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 7190 18204 7196 18216
rect 6871 18176 7196 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 7760 18213 7788 18312
rect 9324 18272 9352 18368
rect 9324 18244 9536 18272
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18204 7803 18207
rect 8018 18204 8024 18216
rect 7791 18176 8024 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 8018 18164 8024 18176
rect 8076 18164 8082 18216
rect 8386 18204 8392 18216
rect 8347 18176 8392 18204
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 9398 18204 9404 18216
rect 8619 18176 9404 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 5350 18136 5356 18148
rect 4172 18108 5356 18136
rect 4172 18077 4200 18108
rect 5350 18096 5356 18108
rect 5408 18096 5414 18148
rect 7374 18136 7380 18148
rect 7287 18108 7380 18136
rect 7374 18096 7380 18108
rect 7432 18136 7438 18148
rect 8404 18136 8432 18164
rect 7432 18108 8432 18136
rect 9508 18136 9536 18244
rect 10321 18207 10379 18213
rect 10321 18173 10333 18207
rect 10367 18204 10379 18207
rect 11054 18204 11060 18216
rect 10367 18176 11060 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 11146 18164 11152 18216
rect 11204 18204 11210 18216
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 11204 18176 11621 18204
rect 11204 18164 11210 18176
rect 11609 18173 11621 18176
rect 11655 18173 11667 18207
rect 11609 18167 11667 18173
rect 9763 18139 9821 18145
rect 9763 18136 9775 18139
rect 9508 18108 9775 18136
rect 7432 18096 7438 18108
rect 9763 18105 9775 18108
rect 9809 18136 9821 18139
rect 10042 18136 10048 18148
rect 9809 18108 10048 18136
rect 9809 18105 9821 18108
rect 9763 18099 9821 18105
rect 10042 18096 10048 18108
rect 10100 18096 10106 18148
rect 4157 18071 4215 18077
rect 4157 18037 4169 18071
rect 4203 18037 4215 18071
rect 5074 18068 5080 18080
rect 5035 18040 5080 18068
rect 4157 18031 4215 18037
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 11333 18071 11391 18077
rect 11333 18068 11345 18071
rect 11204 18040 11345 18068
rect 11204 18028 11210 18040
rect 11333 18037 11345 18040
rect 11379 18037 11391 18071
rect 11333 18031 11391 18037
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 6273 17867 6331 17873
rect 6273 17864 6285 17867
rect 6236 17836 6285 17864
rect 6236 17824 6242 17836
rect 6273 17833 6285 17836
rect 6319 17833 6331 17867
rect 6273 17827 6331 17833
rect 6733 17867 6791 17873
rect 6733 17833 6745 17867
rect 6779 17864 6791 17867
rect 6822 17864 6828 17876
rect 6779 17836 6828 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 8202 17864 8208 17876
rect 7484 17836 8208 17864
rect 5258 17805 5264 17808
rect 5255 17796 5264 17805
rect 5219 17768 5264 17796
rect 5255 17759 5264 17768
rect 5258 17756 5264 17759
rect 5316 17756 5322 17808
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 3142 17728 3148 17740
rect 3007 17700 3148 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 3142 17688 3148 17700
rect 3200 17688 3206 17740
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 5074 17728 5080 17740
rect 4939 17700 5080 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 5074 17688 5080 17700
rect 5132 17688 5138 17740
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 7484 17737 7512 17836
rect 8202 17824 8208 17836
rect 8260 17864 8266 17876
rect 8570 17864 8576 17876
rect 8260 17836 8576 17864
rect 8260 17824 8266 17836
rect 8570 17824 8576 17836
rect 8628 17824 8634 17876
rect 9398 17864 9404 17876
rect 9359 17836 9404 17864
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11422 17864 11428 17876
rect 11112 17836 11428 17864
rect 11112 17824 11118 17836
rect 11422 17824 11428 17836
rect 11480 17864 11486 17876
rect 11480 17836 11652 17864
rect 11480 17824 11486 17836
rect 10042 17805 10048 17808
rect 10039 17796 10048 17805
rect 10003 17768 10048 17796
rect 10039 17759 10048 17768
rect 10042 17756 10048 17759
rect 10100 17756 10106 17808
rect 11514 17796 11520 17808
rect 11475 17768 11520 17796
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 11624 17805 11652 17836
rect 11609 17799 11667 17805
rect 11609 17765 11621 17799
rect 11655 17765 11667 17799
rect 11609 17759 11667 17765
rect 7469 17731 7527 17737
rect 7469 17728 7481 17731
rect 7340 17700 7481 17728
rect 7340 17688 7346 17700
rect 7469 17697 7481 17700
rect 7515 17697 7527 17731
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7469 17691 7527 17697
rect 7576 17700 7941 17728
rect 7006 17620 7012 17672
rect 7064 17660 7070 17672
rect 7576 17660 7604 17700
rect 7929 17697 7941 17700
rect 7975 17728 7987 17731
rect 8110 17728 8116 17740
rect 7975 17700 8116 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 9674 17728 9680 17740
rect 9635 17700 9680 17728
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 8018 17660 8024 17672
rect 7064 17632 7604 17660
rect 7979 17632 8024 17660
rect 7064 17620 7070 17632
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17660 12219 17663
rect 12802 17660 12808 17672
rect 12207 17632 12808 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 3145 17527 3203 17533
rect 3145 17493 3157 17527
rect 3191 17524 3203 17527
rect 4801 17527 4859 17533
rect 4801 17524 4813 17527
rect 3191 17496 4813 17524
rect 3191 17493 3203 17496
rect 3145 17487 3203 17493
rect 4801 17493 4813 17496
rect 4847 17524 4859 17527
rect 4890 17524 4896 17536
rect 4847 17496 4896 17524
rect 4847 17493 4859 17496
rect 4801 17487 4859 17493
rect 4890 17484 4896 17496
rect 4948 17524 4954 17536
rect 5442 17524 5448 17536
rect 4948 17496 5448 17524
rect 4948 17484 4954 17496
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 5718 17484 5724 17536
rect 5776 17524 5782 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5776 17496 5825 17524
rect 5776 17484 5782 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 5813 17487 5871 17493
rect 7101 17527 7159 17533
rect 7101 17493 7113 17527
rect 7147 17524 7159 17527
rect 7190 17524 7196 17536
rect 7147 17496 7196 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 10597 17527 10655 17533
rect 10597 17493 10609 17527
rect 10643 17524 10655 17527
rect 12158 17524 12164 17536
rect 10643 17496 12164 17524
rect 10643 17493 10655 17496
rect 10597 17487 10655 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 3053 17323 3111 17329
rect 3053 17289 3065 17323
rect 3099 17320 3111 17323
rect 3142 17320 3148 17332
rect 3099 17292 3148 17320
rect 3099 17289 3111 17292
rect 3053 17283 3111 17289
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 4246 17320 4252 17332
rect 4207 17292 4252 17320
rect 4246 17280 4252 17292
rect 4304 17280 4310 17332
rect 4617 17323 4675 17329
rect 4617 17289 4629 17323
rect 4663 17320 4675 17323
rect 5074 17320 5080 17332
rect 4663 17292 5080 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 5408 17292 6561 17320
rect 5408 17280 5414 17292
rect 6549 17289 6561 17292
rect 6595 17320 6607 17323
rect 7006 17320 7012 17332
rect 6595 17292 7012 17320
rect 6595 17289 6607 17292
rect 6549 17283 6607 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 8941 17323 8999 17329
rect 8941 17289 8953 17323
rect 8987 17320 8999 17323
rect 10042 17320 10048 17332
rect 8987 17292 10048 17320
rect 8987 17289 8999 17292
rect 8941 17283 8999 17289
rect 4893 17255 4951 17261
rect 4893 17221 4905 17255
rect 4939 17252 4951 17255
rect 5810 17252 5816 17264
rect 4939 17224 5816 17252
rect 4939 17221 4951 17224
rect 4893 17215 4951 17221
rect 5810 17212 5816 17224
rect 5868 17212 5874 17264
rect 7101 17255 7159 17261
rect 7101 17221 7113 17255
rect 7147 17252 7159 17255
rect 7282 17252 7288 17264
rect 7147 17224 7288 17252
rect 7147 17221 7159 17224
rect 7101 17215 7159 17221
rect 7282 17212 7288 17224
rect 7340 17212 7346 17264
rect 4062 17144 4068 17196
rect 4120 17184 4126 17196
rect 5258 17184 5264 17196
rect 4120 17156 4752 17184
rect 5171 17156 5264 17184
rect 4120 17144 4126 17156
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 4246 17116 4252 17128
rect 3743 17088 4252 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 4246 17076 4252 17088
rect 4304 17076 4310 17128
rect 4724 17125 4752 17156
rect 5258 17144 5264 17156
rect 5316 17184 5322 17196
rect 8202 17184 8208 17196
rect 5316 17156 8208 17184
rect 5316 17144 5322 17156
rect 8202 17144 8208 17156
rect 8260 17184 8266 17196
rect 8956 17184 8984 17283
rect 8260 17156 8984 17184
rect 8260 17144 8266 17156
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17116 4767 17119
rect 4755 17088 5580 17116
rect 4755 17085 4767 17088
rect 4709 17079 4767 17085
rect 5552 17057 5580 17088
rect 5626 17076 5632 17128
rect 5684 17116 5690 17128
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 5684 17088 5733 17116
rect 5684 17076 5690 17088
rect 5721 17085 5733 17088
rect 5767 17116 5779 17119
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 5767 17088 6193 17116
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 6181 17085 6193 17088
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 7374 17076 7380 17128
rect 7432 17116 7438 17128
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 7432 17088 7573 17116
rect 7432 17076 7438 17088
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7984 17088 8033 17116
rect 7984 17076 7990 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 9122 17116 9128 17128
rect 8343 17088 9128 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 5537 17051 5595 17057
rect 5537 17017 5549 17051
rect 5583 17048 5595 17051
rect 5994 17048 6000 17060
rect 5583 17020 6000 17048
rect 5583 17017 5595 17020
rect 5537 17011 5595 17017
rect 5994 17008 6000 17020
rect 6052 17008 6058 17060
rect 9508 17057 9536 17292
rect 10042 17280 10048 17292
rect 10100 17320 10106 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 10100 17292 10333 17320
rect 10100 17280 10106 17292
rect 10321 17289 10333 17292
rect 10367 17289 10379 17323
rect 11330 17320 11336 17332
rect 11291 17292 11336 17320
rect 10321 17283 10379 17289
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 11572 17292 11713 17320
rect 11572 17280 11578 17292
rect 11701 17289 11713 17292
rect 11747 17289 11759 17323
rect 12158 17320 12164 17332
rect 12119 17292 12164 17320
rect 11701 17283 11759 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12526 17184 12532 17196
rect 12487 17156 12532 17184
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12802 17184 12808 17196
rect 12763 17156 12808 17184
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 10940 17119 10998 17125
rect 10940 17116 10952 17119
rect 9916 17088 10952 17116
rect 9916 17076 9922 17088
rect 10940 17085 10952 17088
rect 10986 17116 10998 17119
rect 11330 17116 11336 17128
rect 10986 17088 11336 17116
rect 10986 17085 10998 17088
rect 10940 17079 10998 17085
rect 11330 17076 11336 17088
rect 11388 17076 11394 17128
rect 9487 17051 9545 17057
rect 9487 17017 9499 17051
rect 9533 17017 9545 17051
rect 9487 17011 9545 17017
rect 12158 17008 12164 17060
rect 12216 17048 12222 17060
rect 12621 17051 12679 17057
rect 12621 17048 12633 17051
rect 12216 17020 12633 17048
rect 12216 17008 12222 17020
rect 12621 17017 12633 17020
rect 12667 17017 12679 17051
rect 12621 17011 12679 17017
rect 3881 16983 3939 16989
rect 3881 16949 3893 16983
rect 3927 16980 3939 16983
rect 3970 16980 3976 16992
rect 3927 16952 3976 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 5902 16980 5908 16992
rect 5863 16952 5908 16980
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 10042 16980 10048 16992
rect 10003 16952 10048 16980
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 11054 16989 11060 16992
rect 11011 16983 11060 16989
rect 11011 16949 11023 16983
rect 11057 16949 11060 16983
rect 11011 16943 11060 16949
rect 11054 16940 11060 16943
rect 11112 16940 11118 16992
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 3145 16779 3203 16785
rect 3145 16745 3157 16779
rect 3191 16776 3203 16779
rect 4062 16776 4068 16788
rect 3191 16748 4068 16776
rect 3191 16745 3203 16748
rect 3145 16739 3203 16745
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 5810 16776 5816 16788
rect 5771 16748 5816 16776
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 6549 16779 6607 16785
rect 6549 16745 6561 16779
rect 6595 16776 6607 16779
rect 6822 16776 6828 16788
rect 6595 16748 6828 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 9122 16776 9128 16788
rect 9083 16748 9128 16776
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9732 16748 9873 16776
rect 9732 16736 9738 16748
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10100 16748 11376 16776
rect 10100 16736 10106 16748
rect 5350 16708 5356 16720
rect 5000 16680 5356 16708
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 5000 16649 5028 16680
rect 5350 16668 5356 16680
rect 5408 16708 5414 16720
rect 5828 16708 5856 16736
rect 5408 16680 5856 16708
rect 5408 16668 5414 16680
rect 5902 16668 5908 16720
rect 5960 16708 5966 16720
rect 7561 16711 7619 16717
rect 7561 16708 7573 16711
rect 5960 16680 7573 16708
rect 5960 16668 5966 16680
rect 7561 16677 7573 16680
rect 7607 16708 7619 16711
rect 7926 16708 7932 16720
rect 7607 16680 7932 16708
rect 7607 16677 7619 16680
rect 7561 16671 7619 16677
rect 7926 16668 7932 16680
rect 7984 16668 7990 16720
rect 8202 16717 8208 16720
rect 8199 16708 8208 16717
rect 8163 16680 8208 16708
rect 8199 16671 8208 16680
rect 8260 16708 8266 16720
rect 8570 16708 8576 16720
rect 8260 16680 8576 16708
rect 8202 16668 8208 16671
rect 8260 16668 8266 16680
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 10686 16708 10692 16720
rect 10647 16680 10692 16708
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 11348 16708 11376 16748
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11480 16748 11529 16776
rect 11480 16736 11486 16748
rect 11517 16745 11529 16748
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 12158 16708 12164 16720
rect 11348 16680 12164 16708
rect 12158 16668 12164 16680
rect 12216 16708 12222 16720
rect 12253 16711 12311 16717
rect 12253 16708 12265 16711
rect 12216 16680 12265 16708
rect 12216 16668 12222 16680
rect 12253 16677 12265 16680
rect 12299 16677 12311 16711
rect 12802 16708 12808 16720
rect 12763 16680 12808 16708
rect 12253 16671 12311 16677
rect 12802 16668 12808 16680
rect 12860 16668 12866 16720
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2924 16612 2973 16640
rect 2924 16600 2930 16612
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 4985 16603 5043 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5261 16603 5319 16609
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 5276 16572 5304 16603
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 6546 16640 6552 16652
rect 6507 16612 6552 16640
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16640 6883 16643
rect 7374 16640 7380 16652
rect 6871 16612 7380 16640
rect 6871 16609 6883 16612
rect 6825 16603 6883 16609
rect 6840 16572 6868 16603
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8018 16640 8024 16652
rect 7883 16612 8024 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8018 16600 8024 16612
rect 8076 16640 8082 16652
rect 8294 16640 8300 16652
rect 8076 16612 8300 16640
rect 8076 16600 8082 16612
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 8757 16643 8815 16649
rect 8757 16609 8769 16643
rect 8803 16640 8815 16643
rect 9582 16640 9588 16652
rect 8803 16612 9588 16640
rect 8803 16609 8815 16612
rect 8757 16603 8815 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10594 16572 10600 16584
rect 4856 16544 6868 16572
rect 10555 16544 10600 16572
rect 4856 16532 4862 16544
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12618 16572 12624 16584
rect 12207 16544 12624 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 11146 16504 11152 16516
rect 11107 16476 11152 16504
rect 11146 16464 11152 16476
rect 11204 16504 11210 16516
rect 12176 16504 12204 16535
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 11204 16476 12204 16504
rect 11204 16464 11210 16476
rect 4617 16439 4675 16445
rect 4617 16405 4629 16439
rect 4663 16436 4675 16439
rect 4890 16436 4896 16448
rect 4663 16408 4896 16436
rect 4663 16405 4675 16408
rect 4617 16399 4675 16405
rect 4890 16396 4896 16408
rect 4948 16436 4954 16448
rect 5626 16436 5632 16448
rect 4948 16408 5632 16436
rect 4948 16396 4954 16408
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 2866 16192 2872 16244
rect 2924 16232 2930 16244
rect 2961 16235 3019 16241
rect 2961 16232 2973 16235
rect 2924 16204 2973 16232
rect 2924 16192 2930 16204
rect 2961 16201 2973 16204
rect 3007 16201 3019 16235
rect 3970 16232 3976 16244
rect 3931 16204 3976 16232
rect 2961 16195 3019 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4798 16232 4804 16244
rect 4759 16204 4804 16232
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 6365 16235 6423 16241
rect 6365 16201 6377 16235
rect 6411 16232 6423 16235
rect 7374 16232 7380 16244
rect 6411 16204 7380 16232
rect 6411 16201 6423 16204
rect 6365 16195 6423 16201
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 8570 16232 8576 16244
rect 8531 16204 8576 16232
rect 8570 16192 8576 16204
rect 8628 16232 8634 16244
rect 8754 16232 8760 16244
rect 8628 16204 8760 16232
rect 8628 16192 8634 16204
rect 8754 16192 8760 16204
rect 8812 16232 8818 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 8812 16204 8953 16232
rect 8812 16192 8818 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 7392 16096 7420 16192
rect 8956 16164 8984 16195
rect 10594 16192 10600 16244
rect 10652 16232 10658 16244
rect 11011 16235 11069 16241
rect 11011 16232 11023 16235
rect 10652 16204 11023 16232
rect 10652 16192 10658 16204
rect 11011 16201 11023 16204
rect 11057 16232 11069 16235
rect 11701 16235 11759 16241
rect 11701 16232 11713 16235
rect 11057 16204 11713 16232
rect 11057 16201 11069 16204
rect 11011 16195 11069 16201
rect 11701 16201 11713 16204
rect 11747 16201 11759 16235
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 11701 16195 11759 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12618 16192 12624 16244
rect 12676 16232 12682 16244
rect 12897 16235 12955 16241
rect 12897 16232 12909 16235
rect 12676 16204 12909 16232
rect 12676 16192 12682 16204
rect 12897 16201 12909 16204
rect 12943 16201 12955 16235
rect 12897 16195 12955 16201
rect 8956 16136 9260 16164
rect 7392 16068 8064 16096
rect 3970 15988 3976 16040
rect 4028 16028 4034 16040
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 4028 16000 4077 16028
rect 4028 15988 4034 16000
rect 4065 15997 4077 16000
rect 4111 15997 4123 16031
rect 5350 16028 5356 16040
rect 5311 16000 5356 16028
rect 4065 15991 4123 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5626 16028 5632 16040
rect 5587 16000 5632 16028
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 8036 16037 8064 16068
rect 8846 16056 8852 16108
rect 8904 16096 8910 16108
rect 9125 16099 9183 16105
rect 9125 16096 9137 16099
rect 8904 16068 9137 16096
rect 8904 16056 8910 16068
rect 9125 16065 9137 16068
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 5810 15960 5816 15972
rect 5771 15932 5816 15960
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 6546 15920 6552 15972
rect 6604 15960 6610 15972
rect 7098 15960 7104 15972
rect 6604 15932 7104 15960
rect 6604 15920 6610 15932
rect 7098 15920 7104 15932
rect 7156 15960 7162 15972
rect 7742 15960 7748 15972
rect 7156 15932 7748 15960
rect 7156 15920 7162 15932
rect 7742 15920 7748 15932
rect 7800 15920 7806 15972
rect 8297 15963 8355 15969
rect 8297 15929 8309 15963
rect 8343 15960 8355 15963
rect 8386 15960 8392 15972
rect 8343 15932 8392 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 8386 15920 8392 15932
rect 8444 15920 8450 15972
rect 9232 15960 9260 16136
rect 12575 16099 12633 16105
rect 12575 16065 12587 16099
rect 12621 16096 12633 16099
rect 12710 16096 12716 16108
rect 12621 16068 12716 16096
rect 12621 16065 12633 16068
rect 12575 16059 12633 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 10940 16031 10998 16037
rect 10940 15997 10952 16031
rect 10986 16028 10998 16031
rect 12488 16031 12546 16037
rect 10986 15997 11008 16028
rect 10940 15991 11008 15997
rect 12488 15997 12500 16031
rect 12534 16028 12546 16031
rect 12802 16028 12808 16040
rect 12534 16000 12808 16028
rect 12534 15997 12546 16000
rect 12488 15991 12546 15997
rect 9446 15963 9504 15969
rect 9446 15960 9458 15963
rect 9232 15932 9458 15960
rect 9446 15929 9458 15932
rect 9492 15960 9504 15963
rect 9950 15960 9956 15972
rect 9492 15932 9956 15960
rect 9492 15929 9504 15932
rect 9446 15923 9504 15929
rect 9950 15920 9956 15932
rect 10008 15920 10014 15972
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 6564 15892 6592 15920
rect 4295 15864 6592 15892
rect 10045 15895 10103 15901
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10594 15892 10600 15904
rect 10091 15864 10600 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 10980 15892 11008 15991
rect 12802 15988 12808 16000
rect 12860 16028 12866 16040
rect 13265 16031 13323 16037
rect 13265 16028 13277 16031
rect 12860 16000 13277 16028
rect 12860 15988 12866 16000
rect 13265 15997 13277 16000
rect 13311 15997 13323 16031
rect 13265 15991 13323 15997
rect 11333 15895 11391 15901
rect 11333 15892 11345 15895
rect 10928 15864 11345 15892
rect 10928 15852 10934 15864
rect 11333 15861 11345 15864
rect 11379 15861 11391 15895
rect 11333 15855 11391 15861
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 5350 15688 5356 15700
rect 4847 15660 5356 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 6822 15688 6828 15700
rect 6735 15660 6828 15688
rect 6822 15648 6828 15660
rect 6880 15688 6886 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6880 15660 7021 15688
rect 6880 15648 6886 15660
rect 7009 15657 7021 15660
rect 7055 15657 7067 15691
rect 7009 15651 7067 15657
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7892 15660 7941 15688
rect 7892 15648 7898 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 8294 15688 8300 15700
rect 8255 15660 8300 15688
rect 7929 15651 7987 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8662 15688 8668 15700
rect 8623 15660 8668 15688
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 8904 15660 9137 15688
rect 8904 15648 8910 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 10652 15660 11652 15688
rect 10652 15648 10658 15660
rect 5258 15580 5264 15632
rect 5316 15620 5322 15632
rect 5442 15620 5448 15632
rect 5316 15592 5448 15620
rect 5316 15580 5322 15592
rect 5442 15580 5448 15592
rect 5500 15629 5506 15632
rect 5500 15623 5549 15629
rect 5500 15589 5503 15623
rect 5537 15589 5549 15623
rect 5500 15583 5549 15589
rect 5500 15580 5506 15583
rect 5626 15580 5632 15632
rect 5684 15620 5690 15632
rect 5684 15592 7420 15620
rect 5684 15580 5690 15592
rect 7098 15552 7104 15564
rect 7059 15524 7104 15552
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 7392 15561 7420 15592
rect 9950 15580 9956 15632
rect 10008 15629 10014 15632
rect 10008 15623 10056 15629
rect 10008 15589 10010 15623
rect 10044 15589 10056 15623
rect 10008 15583 10056 15589
rect 10008 15580 10014 15583
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 11514 15620 11520 15632
rect 11112 15592 11520 15620
rect 11112 15580 11118 15592
rect 11514 15580 11520 15592
rect 11572 15580 11578 15632
rect 11624 15629 11652 15660
rect 11609 15623 11667 15629
rect 11609 15589 11621 15623
rect 11655 15620 11667 15623
rect 11698 15620 11704 15632
rect 11655 15592 11704 15620
rect 11655 15589 11667 15592
rect 11609 15583 11667 15589
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 7377 15555 7435 15561
rect 7377 15521 7389 15555
rect 7423 15552 7435 15555
rect 8018 15552 8024 15564
rect 7423 15524 8024 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8478 15552 8484 15564
rect 8439 15524 8484 15552
rect 8478 15512 8484 15524
rect 8536 15512 8542 15564
rect 9677 15555 9735 15561
rect 9677 15521 9689 15555
rect 9723 15552 9735 15555
rect 9766 15552 9772 15564
rect 9723 15524 9772 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 12986 15552 12992 15564
rect 13044 15561 13050 15564
rect 13044 15555 13082 15561
rect 12308 15524 12992 15552
rect 12308 15512 12314 15524
rect 12986 15512 12992 15524
rect 13070 15521 13082 15555
rect 13044 15515 13082 15521
rect 13044 15512 13050 15515
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5810 15484 5816 15496
rect 5215 15456 5816 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15484 12219 15487
rect 12342 15484 12348 15496
rect 12207 15456 12348 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 6086 15348 6092 15360
rect 6047 15320 6092 15348
rect 6086 15308 6092 15320
rect 6144 15308 6150 15360
rect 10594 15348 10600 15360
rect 10555 15320 10600 15348
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 12802 15308 12808 15360
rect 12860 15348 12866 15360
rect 13127 15351 13185 15357
rect 13127 15348 13139 15351
rect 12860 15320 13139 15348
rect 12860 15308 12866 15320
rect 13127 15317 13139 15320
rect 13173 15317 13185 15351
rect 13127 15311 13185 15317
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5500 15116 6009 15144
rect 5500 15104 5506 15116
rect 5997 15113 6009 15116
rect 6043 15144 6055 15147
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 6043 15116 6561 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 8018 15144 8024 15156
rect 7979 15116 8024 15144
rect 6549 15107 6607 15113
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4212 14912 4905 14940
rect 4212 14900 4218 14912
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5258 14940 5264 14952
rect 4939 14912 5264 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 5626 14940 5632 14952
rect 5491 14912 5632 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 5460 14872 5488 14903
rect 5626 14900 5632 14912
rect 5684 14900 5690 14952
rect 4540 14844 5488 14872
rect 6564 14872 6592 15107
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 8478 15144 8484 15156
rect 8439 15116 8484 15144
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 8754 15144 8760 15156
rect 8715 15116 8760 15144
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10008 15116 10149 15144
rect 10008 15104 10014 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10594 15144 10600 15156
rect 10555 15116 10600 15144
rect 10137 15107 10195 15113
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 11698 15144 11704 15156
rect 11659 15116 11704 15144
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 13538 15104 13544 15156
rect 13596 15144 13602 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13596 15116 13921 15144
rect 13596 15104 13602 15116
rect 6822 15008 6828 15020
rect 6783 14980 6828 15008
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 8938 15008 8944 15020
rect 8444 14980 8944 15008
rect 8444 14968 8450 14980
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 10962 15008 10968 15020
rect 10827 14980 10968 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 10962 14968 10968 14980
rect 11020 15008 11026 15020
rect 13587 15011 13645 15017
rect 13587 15008 13599 15011
rect 11020 14980 13599 15008
rect 11020 14968 11026 14980
rect 13587 14977 13599 14980
rect 13633 14977 13645 15011
rect 13587 14971 13645 14977
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12488 14943 12546 14949
rect 12488 14940 12500 14943
rect 12299 14912 12500 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12488 14909 12500 14912
rect 12534 14940 12546 14943
rect 12710 14940 12716 14952
rect 12534 14912 12716 14940
rect 12534 14909 12546 14912
rect 12488 14903 12546 14909
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 13500 14943 13558 14949
rect 13500 14940 13512 14943
rect 13320 14912 13512 14940
rect 13320 14900 13326 14912
rect 13500 14909 13512 14912
rect 13546 14940 13558 14943
rect 13740 14940 13768 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 13909 15107 13967 15113
rect 13546 14912 13768 14940
rect 13546 14909 13558 14912
rect 13500 14903 13558 14909
rect 7146 14875 7204 14881
rect 7146 14872 7158 14875
rect 6564 14844 7158 14872
rect 4540 14816 4568 14844
rect 7146 14841 7158 14844
rect 7192 14841 7204 14875
rect 7146 14835 7204 14841
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 9262 14875 9320 14881
rect 9262 14872 9274 14875
rect 8812 14844 9274 14872
rect 8812 14832 8818 14844
rect 9262 14841 9274 14844
rect 9308 14841 9320 14875
rect 9262 14835 9320 14841
rect 10594 14832 10600 14884
rect 10652 14872 10658 14884
rect 10873 14875 10931 14881
rect 10873 14872 10885 14875
rect 10652 14844 10885 14872
rect 10652 14832 10658 14844
rect 10873 14841 10885 14844
rect 10919 14841 10931 14875
rect 10873 14835 10931 14841
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11425 14875 11483 14881
rect 11425 14872 11437 14875
rect 11112 14844 11437 14872
rect 11112 14832 11118 14844
rect 11425 14841 11437 14844
rect 11471 14841 11483 14875
rect 11425 14835 11483 14841
rect 4522 14804 4528 14816
rect 4483 14776 4528 14804
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 5258 14804 5264 14816
rect 5219 14776 5264 14804
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 6822 14804 6828 14816
rect 6696 14776 6828 14804
rect 6696 14764 6702 14776
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 9858 14804 9864 14816
rect 9819 14776 9864 14804
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12575 14807 12633 14813
rect 12575 14804 12587 14807
rect 12032 14776 12587 14804
rect 12032 14764 12038 14776
rect 12575 14773 12587 14776
rect 12621 14773 12633 14807
rect 12986 14804 12992 14816
rect 12947 14776 12992 14804
rect 12575 14767 12633 14773
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 5316 14572 5457 14600
rect 5316 14560 5322 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5445 14563 5503 14569
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 7156 14572 7389 14600
rect 7156 14560 7162 14572
rect 7377 14569 7389 14572
rect 7423 14569 7435 14603
rect 7377 14563 7435 14569
rect 7837 14603 7895 14609
rect 7837 14569 7849 14603
rect 7883 14600 7895 14603
rect 8478 14600 8484 14612
rect 7883 14572 8484 14600
rect 7883 14569 7895 14572
rect 7837 14563 7895 14569
rect 6549 14535 6607 14541
rect 6549 14501 6561 14535
rect 6595 14532 6607 14535
rect 6638 14532 6644 14544
rect 6595 14504 6644 14532
rect 6595 14501 6607 14504
rect 6549 14495 6607 14501
rect 6638 14492 6644 14504
rect 6696 14532 6702 14544
rect 7742 14532 7748 14544
rect 6696 14504 7748 14532
rect 6696 14492 6702 14504
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 5074 14473 5080 14476
rect 5052 14467 5080 14473
rect 5052 14433 5064 14467
rect 5052 14427 5080 14433
rect 5074 14424 5080 14427
rect 5132 14424 5138 14476
rect 8110 14464 8116 14476
rect 8071 14436 8116 14464
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8404 14473 8432 14572
rect 8478 14560 8484 14572
rect 8536 14600 8542 14612
rect 8662 14600 8668 14612
rect 8536 14572 8668 14600
rect 8536 14560 8542 14572
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 8938 14600 8944 14612
rect 8899 14572 8944 14600
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9824 14572 9965 14600
rect 9824 14560 9830 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 11514 14600 11520 14612
rect 11475 14572 11520 14600
rect 9953 14563 10011 14569
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 10505 14535 10563 14541
rect 10505 14532 10517 14535
rect 9916 14504 10517 14532
rect 9916 14492 9922 14504
rect 10505 14501 10517 14504
rect 10551 14532 10563 14535
rect 11146 14532 11152 14544
rect 10551 14504 11152 14532
rect 10551 14501 10563 14504
rect 10505 14495 10563 14501
rect 11146 14492 11152 14504
rect 11204 14532 11210 14544
rect 12069 14535 12127 14541
rect 12069 14532 12081 14535
rect 11204 14504 12081 14532
rect 11204 14492 11210 14504
rect 12069 14501 12081 14504
rect 12115 14501 12127 14535
rect 12069 14495 12127 14501
rect 12434 14492 12440 14544
rect 12492 14532 12498 14544
rect 12621 14535 12679 14541
rect 12621 14532 12633 14535
rect 12492 14504 12633 14532
rect 12492 14492 12498 14504
rect 12621 14501 12633 14504
rect 12667 14501 12679 14535
rect 12621 14495 12679 14501
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11112 14436 11157 14464
rect 11112 14424 11118 14436
rect 6454 14396 6460 14408
rect 6415 14368 6460 14396
rect 6454 14356 6460 14368
rect 6512 14356 6518 14408
rect 7098 14396 7104 14408
rect 7059 14368 7104 14396
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8481 14399 8539 14405
rect 8481 14396 8493 14399
rect 8352 14368 8493 14396
rect 8352 14356 8358 14368
rect 8481 14365 8493 14368
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 11606 14396 11612 14408
rect 10459 14368 11612 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14396 12035 14399
rect 12802 14396 12808 14408
rect 12023 14368 12808 14396
rect 12023 14365 12035 14368
rect 11977 14359 12035 14365
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 5123 14263 5181 14269
rect 5123 14260 5135 14263
rect 4304 14232 5135 14260
rect 4304 14220 4310 14232
rect 5123 14229 5135 14232
rect 5169 14229 5181 14263
rect 5123 14223 5181 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 3007 14059 3065 14065
rect 3007 14025 3019 14059
rect 3053 14056 3065 14059
rect 4062 14056 4068 14068
rect 3053 14028 4068 14056
rect 3053 14025 3065 14028
rect 3007 14019 3065 14025
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4430 14056 4436 14068
rect 4391 14028 4436 14056
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 5074 14056 5080 14068
rect 4847 14028 5080 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 3418 13988 3424 14000
rect 3379 13960 3424 13988
rect 3418 13948 3424 13960
rect 3476 13948 3482 14000
rect 4448 13988 4476 14016
rect 3931 13960 4476 13988
rect 2936 13855 2994 13861
rect 2936 13821 2948 13855
rect 2982 13852 2994 13855
rect 3436 13852 3464 13948
rect 3931 13861 3959 13960
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4816 13920 4844 14019
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 6273 14059 6331 14065
rect 6273 14025 6285 14059
rect 6319 14056 6331 14059
rect 6638 14056 6644 14068
rect 6319 14028 6644 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 6638 14016 6644 14028
rect 6696 14056 6702 14068
rect 7006 14056 7012 14068
rect 6696 14028 7012 14056
rect 6696 14016 6702 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8110 14056 8116 14068
rect 8067 14028 8116 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 10045 14059 10103 14065
rect 10045 14025 10057 14059
rect 10091 14056 10103 14059
rect 10318 14056 10324 14068
rect 10091 14028 10324 14056
rect 10091 14025 10103 14028
rect 10045 14019 10103 14025
rect 10318 14016 10324 14028
rect 10376 14056 10382 14068
rect 10594 14056 10600 14068
rect 10376 14028 10600 14056
rect 10376 14016 10382 14028
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11606 14056 11612 14068
rect 11519 14028 11612 14056
rect 11606 14016 11612 14028
rect 11664 14056 11670 14068
rect 11974 14056 11980 14068
rect 11664 14028 11980 14056
rect 11664 14016 11670 14028
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12713 14059 12771 14065
rect 12713 14025 12725 14059
rect 12759 14056 12771 14059
rect 12802 14056 12808 14068
rect 12759 14028 12808 14056
rect 12759 14025 12771 14028
rect 12713 14019 12771 14025
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 11164 13988 11192 14016
rect 11885 13991 11943 13997
rect 11885 13988 11897 13991
rect 11164 13960 11897 13988
rect 11885 13957 11897 13960
rect 11931 13957 11943 13991
rect 11885 13951 11943 13957
rect 4212 13892 4844 13920
rect 4893 13923 4951 13929
rect 4212 13880 4218 13892
rect 4893 13889 4905 13923
rect 4939 13920 4951 13923
rect 5258 13920 5264 13932
rect 4939 13892 5264 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 6972 13892 9413 13920
rect 6972 13880 6978 13892
rect 4062 13861 4068 13864
rect 2982 13824 3464 13852
rect 3916 13855 3974 13861
rect 2982 13821 2994 13824
rect 2936 13815 2994 13821
rect 3916 13821 3928 13855
rect 3962 13821 3974 13855
rect 3916 13815 3974 13821
rect 4019 13855 4068 13861
rect 4019 13821 4031 13855
rect 4065 13821 4068 13855
rect 4019 13815 4068 13821
rect 4062 13812 4068 13815
rect 4120 13812 4126 13864
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 5813 13855 5871 13861
rect 5813 13852 5825 13855
rect 5592 13824 5825 13852
rect 5592 13812 5598 13824
rect 5813 13821 5825 13824
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 7616 13824 7661 13852
rect 7616 13812 7622 13824
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8168 13824 8401 13852
rect 8168 13812 8174 13824
rect 8389 13821 8401 13824
rect 8435 13852 8447 13855
rect 8754 13852 8760 13864
rect 8435 13824 8760 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 8864 13861 8892 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 10873 13923 10931 13929
rect 10873 13889 10885 13923
rect 10919 13920 10931 13923
rect 12434 13920 12440 13932
rect 10919 13892 12440 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 5258 13793 5264 13796
rect 5255 13747 5264 13793
rect 5316 13784 5322 13796
rect 6914 13784 6920 13796
rect 5316 13756 5355 13784
rect 6875 13756 6920 13784
rect 5258 13744 5264 13747
rect 5316 13744 5322 13756
rect 6914 13744 6920 13756
rect 6972 13744 6978 13796
rect 7006 13744 7012 13796
rect 7064 13784 7070 13796
rect 10226 13784 10232 13796
rect 7064 13756 7109 13784
rect 10187 13756 10232 13784
rect 7064 13744 7070 13756
rect 10226 13744 10232 13756
rect 10284 13744 10290 13796
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10376 13756 10421 13784
rect 10376 13744 10382 13756
rect 8662 13716 8668 13728
rect 8623 13688 8668 13716
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 5258 13472 5264 13484
rect 5316 13512 5322 13524
rect 5316 13484 6224 13512
rect 5316 13472 5322 13484
rect 4246 13444 4252 13456
rect 4207 13416 4252 13444
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 4338 13404 4344 13456
rect 4396 13444 4402 13456
rect 5442 13444 5448 13456
rect 4396 13416 5448 13444
rect 4396 13404 4402 13416
rect 5442 13404 5448 13416
rect 5500 13404 5506 13456
rect 5813 13447 5871 13453
rect 5813 13444 5825 13447
rect 5644 13416 5825 13444
rect 4982 13336 4988 13388
rect 5040 13376 5046 13388
rect 5644 13376 5672 13416
rect 5813 13413 5825 13416
rect 5859 13413 5871 13447
rect 5813 13407 5871 13413
rect 5905 13447 5963 13453
rect 5905 13413 5917 13447
rect 5951 13444 5963 13447
rect 6086 13444 6092 13456
rect 5951 13416 6092 13444
rect 5951 13413 5963 13416
rect 5905 13407 5963 13413
rect 6086 13404 6092 13416
rect 6144 13404 6150 13456
rect 6196 13444 6224 13484
rect 6638 13472 6644 13524
rect 6696 13512 6702 13524
rect 6733 13515 6791 13521
rect 6733 13512 6745 13515
rect 6696 13484 6745 13512
rect 6696 13472 6702 13484
rect 6733 13481 6745 13484
rect 6779 13481 6791 13515
rect 6733 13475 6791 13481
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7101 13515 7159 13521
rect 7101 13512 7113 13515
rect 6972 13484 7113 13512
rect 6972 13472 6978 13484
rect 7101 13481 7113 13484
rect 7147 13481 7159 13515
rect 7101 13475 7159 13481
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 8849 13515 8907 13521
rect 8849 13512 8861 13515
rect 8812 13484 8861 13512
rect 8812 13472 8818 13484
rect 8849 13481 8861 13484
rect 8895 13481 8907 13515
rect 8849 13475 8907 13481
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10284 13484 10701 13512
rect 10284 13472 10290 13484
rect 10689 13481 10701 13484
rect 10735 13512 10747 13515
rect 11379 13515 11437 13521
rect 11379 13512 11391 13515
rect 10735 13484 11391 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 11379 13481 11391 13484
rect 11425 13481 11437 13515
rect 11379 13475 11437 13481
rect 7650 13444 7656 13456
rect 6196 13416 7656 13444
rect 7650 13404 7656 13416
rect 7708 13444 7714 13456
rect 7974 13447 8032 13453
rect 7974 13444 7986 13447
rect 7708 13416 7986 13444
rect 7708 13404 7714 13416
rect 7974 13413 7986 13416
rect 8020 13413 8032 13447
rect 9858 13444 9864 13456
rect 9819 13416 9864 13444
rect 7974 13407 8032 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 5040 13348 5672 13376
rect 5040 13336 5046 13348
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11276 13379 11334 13385
rect 11276 13376 11288 13379
rect 11204 13348 11288 13376
rect 11204 13336 11210 13348
rect 11276 13345 11288 13348
rect 11322 13345 11334 13379
rect 11276 13339 11334 13345
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 5626 13308 5632 13320
rect 4939 13280 5632 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 5868 13280 6469 13308
rect 5868 13268 5874 13280
rect 6457 13277 6469 13280
rect 6503 13308 6515 13311
rect 7558 13308 7564 13320
rect 6503 13280 7564 13308
rect 6503 13277 6515 13280
rect 6457 13271 6515 13277
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 8662 13308 8668 13320
rect 7699 13280 8668 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 9766 13308 9772 13320
rect 9727 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 10502 13308 10508 13320
rect 10459 13280 10508 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 8570 13172 8576 13184
rect 8531 13144 8576 13172
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 3697 12971 3755 12977
rect 3697 12937 3709 12971
rect 3743 12968 3755 12971
rect 4246 12968 4252 12980
rect 3743 12940 4252 12968
rect 3743 12937 3755 12940
rect 3697 12931 3755 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 6144 12940 6193 12968
rect 6144 12928 6150 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 7650 12968 7656 12980
rect 7611 12940 7656 12968
rect 6181 12931 6239 12937
rect 7650 12928 7656 12940
rect 7708 12928 7714 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 8941 12971 8999 12977
rect 8941 12968 8953 12971
rect 8720 12940 8953 12968
rect 8720 12928 8726 12940
rect 8941 12937 8953 12940
rect 8987 12937 8999 12971
rect 8941 12931 8999 12937
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 9824 12940 10885 12968
rect 9824 12928 9830 12940
rect 10873 12937 10885 12940
rect 10919 12968 10931 12971
rect 11054 12968 11060 12980
rect 10919 12940 11060 12968
rect 10919 12937 10931 12940
rect 10873 12931 10931 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11204 12940 11897 12968
rect 11204 12928 11210 12940
rect 11885 12937 11897 12940
rect 11931 12968 11943 12971
rect 12526 12968 12532 12980
rect 11931 12940 12532 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 4065 12903 4123 12909
rect 4065 12869 4077 12903
rect 4111 12900 4123 12903
rect 4338 12900 4344 12912
rect 4111 12872 4344 12900
rect 4111 12869 4123 12872
rect 4065 12863 4123 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 5810 12900 5816 12912
rect 5771 12872 5816 12900
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 5040 12804 6561 12832
rect 5040 12792 5046 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12832 7343 12835
rect 7745 12835 7803 12841
rect 7745 12832 7757 12835
rect 7331 12804 7757 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 7745 12801 7757 12804
rect 7791 12832 7803 12835
rect 8202 12832 8208 12844
rect 7791 12804 8208 12832
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 9858 12832 9864 12844
rect 8680 12804 9864 12832
rect 4208 12767 4266 12773
rect 4208 12733 4220 12767
rect 4254 12764 4266 12767
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4254 12736 4629 12764
rect 4254 12733 4266 12736
rect 4208 12727 4266 12733
rect 4617 12733 4629 12736
rect 4663 12764 4675 12767
rect 5074 12764 5080 12776
rect 4663 12736 5080 12764
rect 4663 12733 4675 12736
rect 4617 12727 4675 12733
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 4295 12699 4353 12705
rect 4295 12665 4307 12699
rect 4341 12696 4353 12699
rect 5258 12696 5264 12708
rect 4341 12668 5264 12696
rect 4341 12665 4353 12668
rect 4295 12659 4353 12665
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 5353 12699 5411 12705
rect 5353 12665 5365 12699
rect 5399 12696 5411 12699
rect 5442 12696 5448 12708
rect 5399 12668 5448 12696
rect 5399 12665 5411 12668
rect 5353 12659 5411 12665
rect 5077 12631 5135 12637
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 5368 12628 5396 12659
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 7650 12656 7656 12708
rect 7708 12696 7714 12708
rect 8066 12699 8124 12705
rect 8066 12696 8078 12699
rect 7708 12668 8078 12696
rect 7708 12656 7714 12668
rect 8066 12665 8078 12668
rect 8112 12665 8124 12699
rect 8066 12659 8124 12665
rect 5123 12600 5396 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 6178 12628 6184 12640
rect 5960 12600 6184 12628
rect 5960 12588 5966 12600
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 8680 12637 8708 12804
rect 9858 12792 9864 12804
rect 9916 12832 9922 12844
rect 10505 12835 10563 12841
rect 10505 12832 10517 12835
rect 9916 12804 10517 12832
rect 9916 12792 9922 12804
rect 10505 12801 10517 12804
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 11146 12773 11152 12776
rect 11124 12767 11152 12773
rect 11124 12733 11136 12767
rect 11204 12764 11210 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 11204 12736 11529 12764
rect 11124 12727 11152 12733
rect 11146 12724 11152 12727
rect 11204 12724 11210 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 9309 12699 9367 12705
rect 9309 12696 9321 12699
rect 8812 12668 9321 12696
rect 8812 12656 8818 12668
rect 9309 12665 9321 12668
rect 9355 12665 9367 12699
rect 9582 12696 9588 12708
rect 9543 12668 9588 12696
rect 9309 12659 9367 12665
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 8260 12600 8677 12628
rect 8260 12588 8266 12600
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 9324 12628 9352 12659
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12665 9735 12699
rect 10226 12696 10232 12708
rect 10187 12668 10232 12696
rect 9677 12659 9735 12665
rect 9692 12628 9720 12659
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 9324 12600 9720 12628
rect 11195 12631 11253 12637
rect 8665 12591 8723 12597
rect 11195 12597 11207 12631
rect 11241 12628 11253 12631
rect 11330 12628 11336 12640
rect 11241 12600 11336 12628
rect 11241 12597 11253 12600
rect 11195 12591 11253 12597
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 4982 12384 4988 12436
rect 5040 12433 5046 12436
rect 5040 12427 5089 12433
rect 5040 12393 5043 12427
rect 5077 12393 5089 12427
rect 5040 12387 5089 12393
rect 5040 12384 5046 12387
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5353 12427 5411 12433
rect 5353 12424 5365 12427
rect 5316 12396 5365 12424
rect 5316 12384 5322 12396
rect 5353 12393 5365 12396
rect 5399 12393 5411 12427
rect 5353 12387 5411 12393
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 7098 12424 7104 12436
rect 5684 12396 7104 12424
rect 5684 12384 5690 12396
rect 6089 12359 6147 12365
rect 6089 12325 6101 12359
rect 6135 12356 6147 12359
rect 6178 12356 6184 12368
rect 6135 12328 6184 12356
rect 6135 12325 6147 12328
rect 6089 12319 6147 12325
rect 6178 12316 6184 12328
rect 6236 12316 6242 12368
rect 6656 12365 6684 12396
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 7708 12396 7849 12424
rect 7708 12384 7714 12396
rect 7837 12393 7849 12396
rect 7883 12424 7895 12427
rect 7926 12424 7932 12436
rect 7883 12396 7932 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 7926 12384 7932 12396
rect 7984 12424 7990 12436
rect 9950 12424 9956 12436
rect 7984 12396 9956 12424
rect 7984 12384 7990 12396
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 10560 12396 12020 12424
rect 10560 12384 10566 12396
rect 6641 12359 6699 12365
rect 6641 12325 6653 12359
rect 6687 12356 6699 12359
rect 6687 12328 6721 12356
rect 6687 12325 6699 12328
rect 6641 12319 6699 12325
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 8110 12356 8116 12368
rect 7340 12328 8116 12356
rect 7340 12316 7346 12328
rect 8110 12316 8116 12328
rect 8168 12356 8174 12368
rect 8205 12359 8263 12365
rect 8205 12356 8217 12359
rect 8168 12328 8217 12356
rect 8168 12316 8174 12328
rect 8205 12325 8217 12328
rect 8251 12325 8263 12359
rect 8205 12319 8263 12325
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 9490 12356 9496 12368
rect 8628 12328 9496 12356
rect 8628 12316 8634 12328
rect 9490 12316 9496 12328
rect 9548 12356 9554 12368
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 9548 12328 9873 12356
rect 9548 12316 9554 12328
rect 9861 12325 9873 12328
rect 9907 12356 9919 12359
rect 11422 12356 11428 12368
rect 9907 12328 11428 12356
rect 9907 12325 9919 12328
rect 9861 12319 9919 12325
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 11992 12365 12020 12396
rect 11977 12359 12035 12365
rect 11977 12325 11989 12359
rect 12023 12325 12035 12359
rect 11977 12319 12035 12325
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 4928 12291 4986 12297
rect 4928 12288 4940 12291
rect 4764 12260 4940 12288
rect 4764 12248 4770 12260
rect 4928 12257 4940 12260
rect 4974 12257 4986 12291
rect 4928 12251 4986 12257
rect 12802 12248 12808 12300
rect 12860 12297 12866 12300
rect 12860 12291 12898 12297
rect 12886 12257 12898 12291
rect 12860 12251 12898 12257
rect 12860 12248 12866 12251
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5684 12192 6009 12220
rect 5684 12180 5690 12192
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 8113 12223 8171 12229
rect 8113 12220 8125 12223
rect 7892 12192 8125 12220
rect 7892 12180 7898 12192
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9456 12192 9781 12220
rect 9456 12180 9462 12192
rect 9769 12189 9781 12192
rect 9815 12220 9827 12223
rect 11330 12220 11336 12232
rect 9815 12192 10548 12220
rect 11291 12192 11336 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 8018 12152 8024 12164
rect 7708 12124 8024 12152
rect 7708 12112 7714 12124
rect 8018 12112 8024 12124
rect 8076 12112 8082 12164
rect 8665 12155 8723 12161
rect 8665 12121 8677 12155
rect 8711 12152 8723 12155
rect 10226 12152 10232 12164
rect 8711 12124 10232 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 10226 12112 10232 12124
rect 10284 12152 10290 12164
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 10284 12124 10333 12152
rect 10284 12112 10290 12124
rect 10321 12121 10333 12124
rect 10367 12121 10379 12155
rect 10520 12152 10548 12192
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 12943 12223 13001 12229
rect 12943 12220 12955 12223
rect 11440 12192 12955 12220
rect 11440 12152 11468 12192
rect 12943 12189 12955 12192
rect 12989 12189 13001 12223
rect 12943 12183 13001 12189
rect 10520 12124 11468 12152
rect 10321 12115 10379 12121
rect 9493 12087 9551 12093
rect 9493 12053 9505 12087
rect 9539 12084 9551 12087
rect 9582 12084 9588 12096
rect 9539 12056 9588 12084
rect 9539 12053 9551 12056
rect 9493 12047 9551 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 4893 11883 4951 11889
rect 4893 11849 4905 11883
rect 4939 11880 4951 11883
rect 5350 11880 5356 11892
rect 4939 11852 5356 11880
rect 4939 11849 4951 11852
rect 4893 11843 4951 11849
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 5810 11880 5816 11892
rect 5675 11852 5816 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 5166 11812 5172 11824
rect 4764 11784 5172 11812
rect 4764 11772 4770 11784
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 5644 11676 5672 11843
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6236 11852 6561 11880
rect 6236 11840 6242 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 6549 11843 6607 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 8665 11883 8723 11889
rect 8665 11849 8677 11883
rect 8711 11880 8723 11883
rect 8754 11880 8760 11892
rect 8711 11852 8760 11880
rect 8711 11849 8723 11852
rect 8665 11843 8723 11849
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 9490 11880 9496 11892
rect 9451 11852 9496 11880
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 11149 11883 11207 11889
rect 11149 11849 11161 11883
rect 11195 11880 11207 11883
rect 11330 11880 11336 11892
rect 11195 11852 11336 11880
rect 11195 11849 11207 11852
rect 11149 11843 11207 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 11480 11852 12081 11880
rect 11480 11840 11486 11852
rect 12069 11849 12081 11852
rect 12115 11849 12127 11883
rect 12069 11843 12127 11849
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 13265 11883 13323 11889
rect 13265 11880 13277 11883
rect 12860 11852 13277 11880
rect 12860 11840 12866 11852
rect 13265 11849 13277 11852
rect 13311 11849 13323 11883
rect 13265 11843 13323 11849
rect 7653 11815 7711 11821
rect 7653 11781 7665 11815
rect 7699 11812 7711 11815
rect 7926 11812 7932 11824
rect 7699 11784 7932 11812
rect 7699 11781 7711 11784
rect 7653 11775 7711 11781
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9180 11716 9781 11744
rect 9180 11704 9186 11716
rect 9769 11713 9781 11716
rect 9815 11744 9827 11747
rect 10502 11744 10508 11756
rect 9815 11716 10508 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11379 11747 11437 11753
rect 11379 11744 11391 11747
rect 11112 11716 11391 11744
rect 11112 11704 11118 11716
rect 11379 11713 11391 11716
rect 11425 11713 11437 11747
rect 11379 11707 11437 11713
rect 4755 11648 5672 11676
rect 5788 11679 5846 11685
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 5788 11645 5800 11679
rect 5834 11676 5846 11679
rect 6086 11676 6092 11688
rect 5834 11648 6092 11676
rect 5834 11645 5846 11648
rect 5788 11639 5846 11645
rect 6086 11636 6092 11648
rect 6144 11676 6150 11688
rect 6181 11679 6239 11685
rect 6181 11676 6193 11679
rect 6144 11648 6193 11676
rect 6144 11636 6150 11648
rect 6181 11645 6193 11648
rect 6227 11645 6239 11679
rect 7742 11676 7748 11688
rect 7703 11648 7748 11676
rect 6181 11639 6239 11645
rect 7742 11636 7748 11648
rect 7800 11676 7806 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 7800 11648 8953 11676
rect 7800 11636 7806 11648
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 11238 11636 11244 11688
rect 11296 11685 11302 11688
rect 11296 11679 11334 11685
rect 11322 11676 11334 11679
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11322 11648 11713 11676
rect 11322 11645 11334 11648
rect 11296 11639 11334 11645
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 12504 11679 12562 11685
rect 12504 11645 12516 11679
rect 12550 11676 12562 11679
rect 12618 11676 12624 11688
rect 12550 11648 12624 11676
rect 12550 11645 12562 11648
rect 12504 11639 12562 11645
rect 11296 11636 11302 11639
rect 12618 11636 12624 11648
rect 12676 11676 12682 11688
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12676 11648 12909 11676
rect 12676 11636 12682 11648
rect 12897 11645 12909 11648
rect 12943 11676 12955 11679
rect 12986 11676 12992 11688
rect 12943 11648 12992 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 12986 11636 12992 11648
rect 13044 11636 13050 11688
rect 7926 11568 7932 11620
rect 7984 11608 7990 11620
rect 8066 11611 8124 11617
rect 8066 11608 8078 11611
rect 7984 11580 8078 11608
rect 7984 11568 7990 11580
rect 8066 11577 8078 11580
rect 8112 11577 8124 11611
rect 8066 11571 8124 11577
rect 9861 11611 9919 11617
rect 9861 11577 9873 11611
rect 9907 11577 9919 11611
rect 10410 11608 10416 11620
rect 10371 11580 10416 11608
rect 9861 11571 9919 11577
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 5859 11543 5917 11549
rect 5859 11540 5871 11543
rect 5684 11512 5871 11540
rect 5684 11500 5690 11512
rect 5859 11509 5871 11512
rect 5905 11509 5917 11543
rect 5859 11503 5917 11509
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9876 11540 9904 11571
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 9732 11512 10701 11540
rect 9732 11500 9738 11512
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 10689 11503 10747 11509
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 11238 11540 11244 11552
rect 10836 11512 11244 11540
rect 10836 11500 10842 11512
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12575 11543 12633 11549
rect 12575 11540 12587 11543
rect 12492 11512 12587 11540
rect 12492 11500 12498 11512
rect 12575 11509 12587 11512
rect 12621 11509 12633 11543
rect 12575 11503 12633 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 5718 11336 5724 11348
rect 5679 11308 5724 11336
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 6236 11308 6684 11336
rect 6236 11296 6242 11308
rect 4724 11240 6592 11268
rect 4062 11160 4068 11212
rect 4120 11200 4126 11212
rect 4724 11209 4752 11240
rect 6564 11212 6592 11240
rect 4709 11203 4767 11209
rect 4709 11200 4721 11203
rect 4120 11172 4721 11200
rect 4120 11160 4126 11172
rect 4709 11169 4721 11172
rect 4755 11169 4767 11203
rect 4709 11163 4767 11169
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 4856 11172 5273 11200
rect 4856 11160 4862 11172
rect 5261 11169 5273 11172
rect 5307 11200 5319 11203
rect 5810 11200 5816 11212
rect 5307 11172 5816 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6546 11200 6552 11212
rect 6507 11172 6552 11200
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 6656 11200 6684 11308
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 7156 11308 7297 11336
rect 7156 11296 7162 11308
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 9122 11336 9128 11348
rect 9083 11308 9128 11336
rect 7285 11299 7343 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9398 11336 9404 11348
rect 9359 11308 9404 11336
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 11379 11339 11437 11345
rect 11379 11305 11391 11339
rect 11425 11336 11437 11339
rect 12066 11336 12072 11348
rect 11425 11308 12072 11336
rect 11425 11305 11437 11308
rect 11379 11299 11437 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 7009 11271 7067 11277
rect 7009 11237 7021 11271
rect 7055 11268 7067 11271
rect 7742 11268 7748 11280
rect 7055 11240 7748 11268
rect 7055 11237 7067 11240
rect 7009 11231 7067 11237
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 8158 11271 8216 11277
rect 8158 11268 8170 11271
rect 7984 11240 8170 11268
rect 7984 11228 7990 11240
rect 8158 11237 8170 11240
rect 8204 11237 8216 11271
rect 8158 11231 8216 11237
rect 9490 11228 9496 11280
rect 9548 11268 9554 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 9548 11240 9873 11268
rect 9548 11228 9554 11240
rect 9861 11237 9873 11240
rect 9907 11237 9919 11271
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 9861 11231 9919 11237
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 6730 11200 6736 11212
rect 6656 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11200 6794 11212
rect 10428 11200 10456 11228
rect 11276 11203 11334 11209
rect 11276 11200 11288 11203
rect 6788 11172 6881 11200
rect 10428 11172 11288 11200
rect 6788 11160 6794 11172
rect 11276 11169 11288 11172
rect 11322 11169 11334 11203
rect 11276 11163 11334 11169
rect 12320 11203 12378 11209
rect 12320 11169 12332 11203
rect 12366 11200 12378 11203
rect 12526 11200 12532 11212
rect 12366 11172 12532 11200
rect 12366 11169 12378 11172
rect 12320 11163 12378 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 5491 11104 7849 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 7837 11101 7849 11104
rect 7883 11132 7895 11135
rect 8294 11132 8300 11144
rect 7883 11104 8300 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 10226 11132 10232 11144
rect 9815 11104 10232 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10226 11092 10232 11104
rect 10284 11132 10290 11144
rect 10962 11132 10968 11144
rect 10284 11104 10968 11132
rect 10284 11092 10290 11104
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 5350 11024 5356 11076
rect 5408 11064 5414 11076
rect 5810 11064 5816 11076
rect 5408 11036 5816 11064
rect 5408 11024 5414 11036
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 7742 11064 7748 11076
rect 7703 11036 7748 11064
rect 7742 11024 7748 11036
rect 7800 11024 7806 11076
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 6089 10999 6147 11005
rect 6089 10996 6101 10999
rect 5684 10968 6101 10996
rect 5684 10956 5690 10968
rect 6089 10965 6101 10968
rect 6135 10965 6147 10999
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 6089 10959 6147 10965
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 12391 10999 12449 11005
rect 12391 10996 12403 10999
rect 11112 10968 12403 10996
rect 11112 10956 11118 10968
rect 12391 10965 12403 10968
rect 12437 10965 12449 10999
rect 12391 10959 12449 10965
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 4062 10792 4068 10804
rect 4023 10764 4068 10792
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10792 6423 10795
rect 6546 10792 6552 10804
rect 6411 10764 6552 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7926 10792 7932 10804
rect 7887 10764 7932 10792
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 9490 10792 9496 10804
rect 8812 10764 9496 10792
rect 8812 10752 8818 10764
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11425 10795 11483 10801
rect 11425 10792 11437 10795
rect 11204 10764 11437 10792
rect 11204 10752 11210 10764
rect 11425 10761 11437 10764
rect 11471 10761 11483 10795
rect 11425 10755 11483 10761
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 12584 10764 12633 10792
rect 12584 10752 12590 10764
rect 12621 10761 12633 10764
rect 12667 10792 12679 10795
rect 13170 10792 13176 10804
rect 12667 10764 13176 10792
rect 12667 10761 12679 10764
rect 12621 10755 12679 10761
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 9125 10727 9183 10733
rect 5552 10696 7236 10724
rect 5552 10668 5580 10696
rect 5534 10656 5540 10668
rect 5495 10628 5540 10656
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7098 10656 7104 10668
rect 6963 10628 7104 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7208 10665 7236 10696
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9306 10724 9312 10736
rect 9171 10696 9312 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 8018 10656 8024 10668
rect 7239 10628 8024 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 8754 10656 8760 10668
rect 8619 10628 8760 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8754 10616 8760 10628
rect 8812 10656 8818 10668
rect 9398 10656 9404 10668
rect 8812 10628 9404 10656
rect 8812 10616 8818 10628
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 10410 10656 10416 10668
rect 10371 10628 10416 10656
rect 10410 10616 10416 10628
rect 10468 10656 10474 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 10468 10628 11805 10656
rect 10468 10616 10474 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 4157 10523 4215 10529
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 5258 10520 5264 10532
rect 4203 10492 5264 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5353 10523 5411 10529
rect 5353 10489 5365 10523
rect 5399 10520 5411 10523
rect 5442 10520 5448 10532
rect 5399 10492 5448 10520
rect 5399 10489 5411 10492
rect 5353 10483 5411 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7064 10492 7109 10520
rect 7064 10480 7070 10492
rect 8662 10480 8668 10532
rect 8720 10520 8726 10532
rect 9953 10523 10011 10529
rect 8720 10492 8765 10520
rect 8720 10480 8726 10492
rect 9953 10489 9965 10523
rect 9999 10520 10011 10523
rect 10134 10520 10140 10532
rect 9999 10492 10140 10520
rect 9999 10489 10011 10492
rect 9953 10483 10011 10489
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 10229 10523 10287 10529
rect 10229 10489 10241 10523
rect 10275 10489 10287 10523
rect 10229 10483 10287 10489
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8680 10452 8708 10480
rect 8435 10424 8708 10452
rect 10244 10452 10272 10483
rect 10594 10452 10600 10464
rect 10244 10424 10600 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 10594 10412 10600 10424
rect 10652 10452 10658 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 10652 10424 11069 10452
rect 10652 10412 10658 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 11057 10415 11115 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 5258 10248 5264 10260
rect 5219 10220 5264 10248
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 6730 10248 6736 10260
rect 6691 10220 6736 10248
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 8294 10248 8300 10260
rect 8255 10220 8300 10248
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 8754 10248 8760 10260
rect 8715 10220 8760 10248
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 10594 10248 10600 10260
rect 10555 10220 10600 10248
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 5899 10183 5957 10189
rect 5899 10149 5911 10183
rect 5945 10180 5957 10183
rect 6270 10180 6276 10192
rect 5945 10152 6276 10180
rect 5945 10149 5957 10152
rect 5899 10143 5957 10149
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 7466 10180 7472 10192
rect 7427 10152 7472 10180
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 8018 10180 8024 10192
rect 7979 10152 8024 10180
rect 8018 10140 8024 10152
rect 8076 10140 8082 10192
rect 10042 10189 10048 10192
rect 10039 10180 10048 10189
rect 10003 10152 10048 10180
rect 10039 10143 10048 10152
rect 10042 10140 10048 10143
rect 10100 10140 10106 10192
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 10192 10152 11437 10180
rect 10192 10140 10198 10152
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 11425 10143 11483 10149
rect 4522 10112 4528 10124
rect 4483 10084 4528 10112
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 7006 10112 7012 10124
rect 6503 10084 7012 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 7006 10072 7012 10084
rect 7064 10112 7070 10124
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 7064 10084 7113 10112
rect 7064 10072 7070 10084
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 10060 10112 10088 10140
rect 10410 10112 10416 10124
rect 10060 10084 10416 10112
rect 7101 10075 7159 10081
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 5534 10044 5540 10056
rect 5495 10016 5540 10044
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 7558 10044 7564 10056
rect 7423 10016 7564 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 7558 10004 7564 10016
rect 7616 10044 7622 10056
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 7616 10016 9045 10044
rect 7616 10004 7622 10016
rect 9033 10013 9045 10016
rect 9079 10013 9091 10047
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9033 10007 9091 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 4522 9704 4528 9716
rect 4483 9676 4528 9704
rect 4522 9664 4528 9676
rect 4580 9664 4586 9716
rect 6270 9704 6276 9716
rect 6183 9676 6276 9704
rect 6270 9664 6276 9676
rect 6328 9704 6334 9716
rect 7926 9704 7932 9716
rect 6328 9676 7932 9704
rect 6328 9664 6334 9676
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 10036 9704 10042 9716
rect 9815 9676 10042 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10036 9664 10042 9676
rect 10094 9704 10100 9716
rect 10410 9704 10416 9716
rect 10094 9676 10416 9704
rect 10094 9664 10100 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 5905 9639 5963 9645
rect 5905 9605 5917 9639
rect 5951 9636 5963 9639
rect 7466 9636 7472 9648
rect 5951 9608 7472 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 7466 9596 7472 9608
rect 7524 9636 7530 9648
rect 7837 9639 7895 9645
rect 7837 9636 7849 9639
rect 7524 9608 7849 9636
rect 7524 9596 7530 9608
rect 7837 9605 7849 9608
rect 7883 9605 7895 9639
rect 7837 9599 7895 9605
rect 7116 9540 8616 9568
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 4203 9472 4997 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4985 9469 4997 9472
rect 5031 9500 5043 9503
rect 5442 9500 5448 9512
rect 5031 9472 5448 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7116 9509 7144 9540
rect 8588 9512 8616 9540
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 9732 9540 10701 9568
rect 9732 9528 9738 9540
rect 10689 9537 10701 9540
rect 10735 9568 10747 9571
rect 11333 9571 11391 9577
rect 11333 9568 11345 9571
rect 10735 9540 11345 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 11333 9537 11345 9540
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 7064 9472 7113 9500
rect 7064 9460 7070 9472
rect 7101 9469 7113 9472
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 7285 9463 7343 9469
rect 4893 9435 4951 9441
rect 4893 9401 4905 9435
rect 4939 9432 4951 9435
rect 5347 9435 5405 9441
rect 5347 9432 5359 9435
rect 4939 9404 5359 9432
rect 4939 9401 4951 9404
rect 4893 9395 4951 9401
rect 5347 9401 5359 9404
rect 5393 9432 5405 9435
rect 6270 9432 6276 9444
rect 5393 9404 6276 9432
rect 5393 9401 5405 9404
rect 5347 9395 5405 9401
rect 6270 9392 6276 9404
rect 6328 9392 6334 9444
rect 7300 9432 7328 9463
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8846 9500 8852 9512
rect 8807 9472 8852 9500
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 10229 9503 10287 9509
rect 10229 9500 10241 9503
rect 9916 9472 10241 9500
rect 9916 9460 9922 9472
rect 10229 9469 10241 9472
rect 10275 9469 10287 9503
rect 10410 9500 10416 9512
rect 10371 9472 10416 9500
rect 10229 9463 10287 9469
rect 6564 9404 7328 9432
rect 8297 9435 8355 9441
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6564 9373 6592 9404
rect 8297 9401 8309 9435
rect 8343 9432 8355 9435
rect 8864 9432 8892 9460
rect 8343 9404 8892 9432
rect 9125 9435 9183 9441
rect 8343 9401 8355 9404
rect 8297 9395 8355 9401
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 9582 9432 9588 9444
rect 9171 9404 9588 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 9582 9392 9588 9404
rect 9640 9392 9646 9444
rect 10244 9432 10272 9463
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10244 9404 10977 9432
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6236 9336 6561 9364
rect 6236 9324 6242 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6914 9364 6920 9376
rect 6875 9336 6920 9364
rect 6549 9327 6607 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 5169 9163 5227 9169
rect 5169 9160 5181 9163
rect 4764 9132 5181 9160
rect 4764 9120 4770 9132
rect 5169 9129 5181 9132
rect 5215 9129 5227 9163
rect 5442 9160 5448 9172
rect 5403 9132 5448 9160
rect 5169 9123 5227 9129
rect 5184 9092 5212 9123
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 5592 9132 6469 9160
rect 5592 9120 5598 9132
rect 6457 9129 6469 9132
rect 6503 9160 6515 9163
rect 6914 9160 6920 9172
rect 6503 9132 6920 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8570 9160 8576 9172
rect 8527 9132 8576 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 8754 9160 8760 9172
rect 8715 9132 8760 9160
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9766 9120 9772 9172
rect 9824 9169 9830 9172
rect 9824 9163 9873 9169
rect 9824 9129 9827 9163
rect 9861 9129 9873 9163
rect 9824 9123 9873 9129
rect 9824 9120 9830 9123
rect 5626 9092 5632 9104
rect 5184 9064 5632 9092
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 7463 9095 7521 9101
rect 7463 9061 7475 9095
rect 7509 9092 7521 9095
rect 7742 9092 7748 9104
rect 7509 9064 7748 9092
rect 7509 9061 7521 9064
rect 7463 9055 7521 9061
rect 7742 9052 7748 9064
rect 7800 9092 7806 9104
rect 7926 9092 7932 9104
rect 7800 9064 7932 9092
rect 7800 9052 7806 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 8772 9092 8800 9120
rect 10410 9092 10416 9104
rect 8772 9064 10416 9092
rect 10410 9052 10416 9064
rect 10468 9092 10474 9104
rect 10505 9095 10563 9101
rect 10505 9092 10517 9095
rect 10468 9064 10517 9092
rect 10468 9052 10474 9064
rect 10505 9061 10517 9064
rect 10551 9061 10563 9095
rect 10505 9055 10563 9061
rect 4338 8984 4344 9036
rect 4396 9033 4402 9036
rect 4396 9027 4434 9033
rect 4422 9024 4434 9027
rect 5258 9024 5264 9036
rect 4422 8996 5264 9024
rect 4422 8993 4434 8996
rect 4396 8987 4434 8993
rect 4396 8984 4402 8987
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 5718 9024 5724 9036
rect 5583 8996 5724 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 6178 9024 6184 9036
rect 5859 8996 6184 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 5828 8956 5856 8987
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7006 9024 7012 9036
rect 6963 8996 7012 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 9744 9027 9802 9033
rect 9744 8993 9756 9027
rect 9790 9024 9802 9027
rect 9950 9024 9956 9036
rect 9790 8996 9956 9024
rect 9790 8993 9802 8996
rect 9744 8987 9802 8993
rect 9950 8984 9956 8996
rect 10008 9024 10014 9036
rect 10134 9024 10140 9036
rect 10008 8996 10140 9024
rect 10008 8984 10014 8996
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10686 9024 10692 9036
rect 10647 8996 10692 9024
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 7098 8956 7104 8968
rect 4580 8928 5856 8956
rect 7059 8928 7104 8956
rect 4580 8916 4586 8928
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 10226 8888 10232 8900
rect 10139 8860 10232 8888
rect 10226 8848 10232 8860
rect 10284 8888 10290 8900
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 10284 8860 10885 8888
rect 10284 8848 10290 8860
rect 10873 8857 10885 8860
rect 10919 8857 10931 8891
rect 10873 8851 10931 8857
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 4479 8823 4537 8829
rect 4479 8820 4491 8823
rect 4120 8792 4491 8820
rect 4120 8780 4126 8792
rect 4479 8789 4491 8792
rect 4525 8789 4537 8823
rect 8018 8820 8024 8832
rect 7979 8792 8024 8820
rect 4479 8783 4537 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4338 8616 4344 8628
rect 4299 8588 4344 8616
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 4488 8588 4629 8616
rect 4488 8576 4494 8588
rect 4617 8585 4629 8588
rect 4663 8585 4675 8619
rect 4617 8579 4675 8585
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 4985 8619 5043 8625
rect 4985 8616 4997 8619
rect 4856 8588 4997 8616
rect 4856 8576 4862 8588
rect 4985 8585 4997 8588
rect 5031 8585 5043 8619
rect 4985 8579 5043 8585
rect 5000 8412 5028 8579
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 5868 8588 6193 8616
rect 5868 8576 5874 8588
rect 6181 8585 6193 8588
rect 6227 8616 6239 8619
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 6227 8588 9229 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 9217 8585 9229 8588
rect 9263 8616 9275 8619
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9263 8588 9505 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10744 8588 10793 8616
rect 10744 8576 10750 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 7742 8548 7748 8560
rect 7703 8520 7748 8548
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 5951 8452 7021 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7009 8449 7021 8452
rect 7055 8480 7067 8483
rect 7098 8480 7104 8492
rect 7055 8452 7104 8480
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7984 8452 8125 8480
rect 7984 8440 7990 8452
rect 8113 8449 8125 8452
rect 8159 8480 8171 8483
rect 8846 8480 8852 8492
rect 8159 8452 8852 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5000 8384 5181 8412
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 5626 8412 5632 8424
rect 5587 8384 5632 8412
rect 5169 8375 5227 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 5994 8412 6000 8424
rect 5868 8384 6000 8412
rect 5868 8372 5874 8384
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8412 8539 8415
rect 8662 8412 8668 8424
rect 8527 8384 8668 8412
rect 8527 8381 8539 8384
rect 8481 8375 8539 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8772 8421 8800 8452
rect 8846 8440 8852 8452
rect 8904 8480 8910 8492
rect 8904 8452 10272 8480
rect 8904 8440 8910 8452
rect 10244 8424 10272 8452
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9769 8415 9827 8421
rect 9769 8412 9781 8415
rect 9539 8384 9781 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9769 8381 9781 8384
rect 9815 8381 9827 8415
rect 10226 8412 10232 8424
rect 10187 8384 10232 8412
rect 9769 8375 9827 8381
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 7193 8347 7251 8353
rect 7193 8313 7205 8347
rect 7239 8344 7251 8347
rect 8110 8344 8116 8356
rect 7239 8316 8116 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 8941 8347 8999 8353
rect 8941 8344 8953 8347
rect 8904 8316 8953 8344
rect 8904 8304 8910 8316
rect 8941 8313 8953 8316
rect 8987 8313 8999 8347
rect 8941 8307 8999 8313
rect 9677 8347 9735 8353
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 9950 8344 9956 8356
rect 9723 8316 9956 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 9950 8304 9956 8316
rect 10008 8344 10014 8356
rect 12250 8344 12256 8356
rect 10008 8316 12256 8344
rect 10008 8304 10014 8316
rect 12250 8304 12256 8316
rect 12308 8304 12314 8356
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 6549 8007 6607 8013
rect 6549 8004 6561 8007
rect 6236 7976 6561 8004
rect 6236 7964 6242 7976
rect 6549 7973 6561 7976
rect 6595 7973 6607 8007
rect 8110 8004 8116 8016
rect 8071 7976 8116 8004
rect 6549 7967 6607 7973
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 10042 8013 10048 8016
rect 10039 8004 10048 8013
rect 10003 7976 10048 8004
rect 10039 7967 10048 7976
rect 10042 7964 10048 7967
rect 10100 7964 10106 8016
rect 5074 7936 5080 7948
rect 5035 7908 5080 7936
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5626 7936 5632 7948
rect 5399 7908 5632 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 6086 7868 6092 7880
rect 5583 7840 6092 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6196 7840 6469 7868
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 6196 7741 6224 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 7098 7868 7104 7880
rect 7059 7840 7104 7868
rect 6457 7831 6515 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7892 7840 8033 7868
rect 7892 7828 7898 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7868 8723 7871
rect 8754 7868 8760 7880
rect 8711 7840 8760 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11112 7840 11437 7868
rect 11112 7828 11118 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 5592 7704 6193 7732
rect 5592 7692 5598 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 10594 7732 10600 7744
rect 10555 7704 10600 7732
rect 6181 7695 6239 7701
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5626 7528 5632 7540
rect 4939 7500 5632 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 7745 7531 7803 7537
rect 7745 7497 7757 7531
rect 7791 7528 7803 7531
rect 8110 7528 8116 7540
rect 7791 7500 8116 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 10781 7531 10839 7537
rect 10781 7528 10793 7531
rect 9732 7500 10793 7528
rect 9732 7488 9738 7500
rect 10781 7497 10793 7500
rect 10827 7497 10839 7531
rect 10781 7491 10839 7497
rect 4525 7463 4583 7469
rect 4525 7429 4537 7463
rect 4571 7460 4583 7463
rect 5074 7460 5080 7472
rect 4571 7432 5080 7460
rect 4571 7429 4583 7432
rect 4525 7423 4583 7429
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 9125 7463 9183 7469
rect 9125 7429 9137 7463
rect 9171 7460 9183 7463
rect 10042 7460 10048 7472
rect 9171 7432 10048 7460
rect 9171 7429 9183 7432
rect 9125 7423 9183 7429
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6144 7364 6837 7392
rect 6144 7352 6150 7364
rect 6825 7361 6837 7364
rect 6871 7392 6883 7395
rect 7006 7392 7012 7404
rect 6871 7364 7012 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 8846 7352 8852 7404
rect 8904 7392 8910 7404
rect 9214 7392 9220 7404
rect 8904 7364 9220 7392
rect 8904 7352 8910 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 5442 7324 5448 7336
rect 5403 7296 5448 7324
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5626 7324 5632 7336
rect 5587 7296 5632 7324
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 6914 7256 6920 7268
rect 5951 7228 6920 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7187 7259 7245 7265
rect 7187 7225 7199 7259
rect 7233 7256 7245 7259
rect 7742 7256 7748 7268
rect 7233 7228 7748 7256
rect 7233 7225 7245 7228
rect 7187 7219 7245 7225
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 6641 7191 6699 7197
rect 6641 7157 6653 7191
rect 6687 7188 6699 7191
rect 7202 7188 7230 7219
rect 7742 7216 7748 7228
rect 7800 7216 7806 7268
rect 9600 7265 9628 7432
rect 10042 7420 10048 7432
rect 10100 7460 10106 7472
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 10100 7432 10425 7460
rect 10100 7420 10106 7432
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 10413 7423 10471 7429
rect 11103 7463 11161 7469
rect 11103 7429 11115 7463
rect 11149 7460 11161 7463
rect 11698 7460 11704 7472
rect 11149 7432 11704 7460
rect 11149 7429 11161 7432
rect 11103 7423 11161 7429
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 11032 7327 11090 7333
rect 11032 7293 11044 7327
rect 11078 7324 11090 7327
rect 11146 7324 11152 7336
rect 11078 7296 11152 7324
rect 11078 7293 11090 7296
rect 11032 7287 11090 7293
rect 11146 7284 11152 7296
rect 11204 7324 11210 7336
rect 11425 7327 11483 7333
rect 11425 7324 11437 7327
rect 11204 7296 11437 7324
rect 11204 7284 11210 7296
rect 11425 7293 11437 7296
rect 11471 7293 11483 7327
rect 11425 7287 11483 7293
rect 9579 7259 9637 7265
rect 9579 7225 9591 7259
rect 9625 7225 9637 7259
rect 9579 7219 9637 7225
rect 6687 7160 7230 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 7834 7188 7840 7200
rect 7340 7160 7840 7188
rect 7340 7148 7346 7160
rect 7834 7148 7840 7160
rect 7892 7188 7898 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 7892 7160 8401 7188
rect 7892 7148 7898 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 10134 7188 10140 7200
rect 10095 7160 10140 7188
rect 8389 7151 8447 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 5353 6987 5411 6993
rect 5353 6953 5365 6987
rect 5399 6984 5411 6987
rect 5626 6984 5632 6996
rect 5399 6956 5632 6984
rect 5399 6953 5411 6956
rect 5353 6947 5411 6953
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 7742 6944 7748 6996
rect 7800 6944 7806 6996
rect 9214 6984 9220 6996
rect 9175 6956 9220 6984
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 10134 6944 10140 6996
rect 10192 6984 10198 6996
rect 10410 6984 10416 6996
rect 10192 6956 10416 6984
rect 10192 6944 10198 6956
rect 10410 6944 10416 6956
rect 10468 6984 10474 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10468 6956 10885 6984
rect 10468 6944 10474 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 5442 6876 5448 6928
rect 5500 6916 5506 6928
rect 6175 6919 6233 6925
rect 5500 6888 5672 6916
rect 5500 6876 5506 6888
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4836 6851 4894 6857
rect 4836 6848 4848 6851
rect 4672 6820 4848 6848
rect 4672 6808 4678 6820
rect 4836 6817 4848 6820
rect 4882 6817 4894 6851
rect 4836 6811 4894 6817
rect 4939 6851 4997 6857
rect 4939 6817 4951 6851
rect 4985 6848 4997 6851
rect 5534 6848 5540 6860
rect 4985 6820 5540 6848
rect 4985 6817 4997 6820
rect 4939 6811 4997 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5644 6848 5672 6888
rect 6175 6885 6187 6919
rect 6221 6916 6233 6919
rect 6546 6916 6552 6928
rect 6221 6888 6552 6916
rect 6221 6885 6233 6888
rect 6175 6879 6233 6885
rect 6546 6876 6552 6888
rect 6604 6916 6610 6928
rect 7760 6916 7788 6944
rect 10042 6925 10048 6928
rect 8066 6919 8124 6925
rect 8066 6916 8078 6919
rect 6604 6888 8078 6916
rect 6604 6876 6610 6888
rect 8066 6885 8078 6888
rect 8112 6885 8124 6919
rect 10039 6916 10048 6925
rect 10003 6888 10048 6916
rect 8066 6879 8124 6885
rect 10039 6879 10048 6888
rect 10042 6876 10048 6879
rect 10100 6876 10106 6928
rect 11609 6919 11667 6925
rect 11609 6916 11621 6919
rect 11348 6888 11621 6916
rect 11348 6860 11376 6888
rect 11609 6885 11621 6888
rect 11655 6885 11667 6919
rect 11609 6879 11667 6885
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 5644 6820 5733 6848
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 6972 6820 7573 6848
rect 6972 6808 6978 6820
rect 7561 6817 7573 6820
rect 7607 6848 7619 6851
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7607 6820 7757 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9858 6848 9864 6860
rect 9723 6820 9864 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 11330 6848 11336 6860
rect 10643 6820 11336 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5684 6752 5825 6780
rect 5684 6740 5690 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 7006 6780 7012 6792
rect 6967 6752 7012 6780
rect 5813 6743 5871 6749
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 11514 6780 11520 6792
rect 11475 6752 11520 6780
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6236 6616 6745 6644
rect 6236 6604 6242 6616
rect 6733 6613 6745 6616
rect 6779 6644 6791 6647
rect 7006 6644 7012 6656
rect 6779 6616 7012 6644
rect 6779 6613 6791 6616
rect 6733 6607 6791 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 8665 6647 8723 6653
rect 8665 6613 8677 6647
rect 8711 6644 8723 6647
rect 8754 6644 8760 6656
rect 8711 6616 8760 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4614 6440 4620 6452
rect 4396 6412 4620 6440
rect 4396 6400 4402 6412
rect 4614 6400 4620 6412
rect 4672 6440 4678 6452
rect 4801 6443 4859 6449
rect 4801 6440 4813 6443
rect 4672 6412 4813 6440
rect 4672 6400 4678 6412
rect 4801 6409 4813 6412
rect 4847 6409 4859 6443
rect 6546 6440 6552 6452
rect 6507 6412 6552 6440
rect 4801 6403 4859 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7800 6412 7849 6440
rect 7800 6400 7806 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8389 6443 8447 6449
rect 8389 6440 8401 6443
rect 8352 6412 8401 6440
rect 8352 6400 8358 6412
rect 8389 6409 8401 6412
rect 8435 6409 8447 6443
rect 8389 6403 8447 6409
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 10042 6440 10048 6452
rect 9815 6412 10048 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 7190 6304 7196 6316
rect 7151 6276 7196 6304
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 8404 6304 8432 6403
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 11425 6443 11483 6449
rect 11425 6440 11437 6443
rect 11388 6412 11437 6440
rect 11388 6400 11394 6412
rect 11425 6409 11437 6412
rect 11471 6409 11483 6443
rect 11425 6403 11483 6409
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11572 6412 11805 6440
rect 11572 6400 11578 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8404 6276 8677 6304
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8938 6304 8944 6316
rect 8899 6276 8944 6304
rect 8665 6267 8723 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 10183 6276 10333 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10321 6273 10333 6276
rect 10367 6304 10379 6307
rect 10962 6304 10968 6316
rect 10367 6276 10968 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 3050 6196 3056 6248
rect 3108 6236 3114 6248
rect 5534 6236 5540 6248
rect 3108 6208 5540 6236
rect 3108 6196 3114 6208
rect 5534 6196 5540 6208
rect 5592 6236 5598 6248
rect 5756 6239 5814 6245
rect 5756 6236 5768 6239
rect 5592 6208 5768 6236
rect 5592 6196 5598 6208
rect 5756 6205 5768 6208
rect 5802 6236 5814 6239
rect 6181 6239 6239 6245
rect 6181 6236 6193 6239
rect 5802 6208 6193 6236
rect 5802 6205 5814 6208
rect 5756 6199 5814 6205
rect 6181 6205 6193 6208
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 5859 6171 5917 6177
rect 5859 6137 5871 6171
rect 5905 6168 5917 6171
rect 6914 6168 6920 6180
rect 5905 6140 6920 6168
rect 5905 6137 5917 6140
rect 5859 6131 5917 6137
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7064 6140 7109 6168
rect 7064 6128 7070 6140
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 8812 6140 8857 6168
rect 8812 6128 8818 6140
rect 10410 6128 10416 6180
rect 10468 6168 10474 6180
rect 10962 6168 10968 6180
rect 10468 6140 10513 6168
rect 10923 6140 10968 6168
rect 10468 6128 10474 6140
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 5626 6100 5632 6112
rect 5587 6072 5632 6100
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 5684 5868 6101 5896
rect 5684 5856 5690 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 6972 5868 7389 5896
rect 6972 5856 6978 5868
rect 7377 5865 7389 5868
rect 7423 5865 7435 5899
rect 8754 5896 8760 5908
rect 8715 5868 8760 5896
rect 7377 5859 7435 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9858 5896 9864 5908
rect 9819 5868 9864 5896
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 5718 5788 5724 5840
rect 5776 5828 5782 5840
rect 7006 5828 7012 5840
rect 5776 5800 6500 5828
rect 6967 5800 7012 5828
rect 5776 5788 5782 5800
rect 6472 5769 6500 5800
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 7098 5788 7104 5840
rect 7156 5828 7162 5840
rect 7745 5831 7803 5837
rect 7745 5828 7757 5831
rect 7156 5800 7757 5828
rect 7156 5788 7162 5800
rect 7745 5797 7757 5800
rect 7791 5797 7803 5831
rect 7745 5791 7803 5797
rect 7837 5831 7895 5837
rect 7837 5797 7849 5831
rect 7883 5828 7895 5831
rect 8018 5828 8024 5840
rect 7883 5800 8024 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 8938 5828 8944 5840
rect 8435 5800 8944 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 10229 5831 10287 5837
rect 10229 5797 10241 5831
rect 10275 5828 10287 5831
rect 10594 5828 10600 5840
rect 10275 5800 10600 5828
rect 10275 5797 10287 5800
rect 10229 5791 10287 5797
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5729 6331 5763
rect 6273 5723 6331 5729
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6546 5760 6552 5772
rect 6503 5732 6552 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 6288 5692 6316 5723
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 10962 5760 10968 5772
rect 10827 5732 10968 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 10962 5720 10968 5732
rect 11020 5760 11026 5772
rect 11676 5763 11734 5769
rect 11676 5760 11688 5763
rect 11020 5732 11688 5760
rect 11020 5720 11026 5732
rect 11676 5729 11688 5732
rect 11722 5760 11734 5763
rect 11974 5760 11980 5772
rect 11722 5732 11980 5760
rect 11722 5729 11734 5732
rect 11676 5723 11734 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 6822 5692 6828 5704
rect 5684 5664 6828 5692
rect 5684 5652 5690 5664
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11514 5556 11520 5568
rect 11020 5528 11520 5556
rect 11020 5516 11026 5528
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 11747 5559 11805 5565
rect 11747 5525 11759 5559
rect 11793 5556 11805 5559
rect 12066 5556 12072 5568
rect 11793 5528 12072 5556
rect 11793 5525 11805 5528
rect 11747 5519 11805 5525
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 5626 5352 5632 5364
rect 5587 5324 5632 5352
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6270 5352 6276 5364
rect 6231 5324 6276 5352
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 6546 5352 6552 5364
rect 6507 5324 6552 5352
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7193 5355 7251 5361
rect 7193 5321 7205 5355
rect 7239 5352 7251 5355
rect 8018 5352 8024 5364
rect 7239 5324 8024 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5352 10379 5355
rect 10594 5352 10600 5364
rect 10367 5324 10600 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 11974 5352 11980 5364
rect 11747 5324 11980 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12894 5352 12900 5364
rect 12855 5324 12900 5352
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 7561 5287 7619 5293
rect 7561 5253 7573 5287
rect 7607 5284 7619 5287
rect 7926 5284 7932 5296
rect 7607 5256 7932 5284
rect 7607 5253 7619 5256
rect 7561 5247 7619 5253
rect 7926 5244 7932 5256
rect 7984 5284 7990 5296
rect 8570 5284 8576 5296
rect 7984 5256 8576 5284
rect 7984 5244 7990 5256
rect 8570 5244 8576 5256
rect 8628 5284 8634 5296
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8628 5256 9045 5284
rect 8628 5244 8634 5256
rect 9033 5253 9045 5256
rect 9079 5253 9091 5287
rect 11238 5284 11244 5296
rect 9033 5247 9091 5253
rect 10831 5256 11244 5284
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6638 5216 6644 5228
rect 5684 5188 6644 5216
rect 5684 5176 5690 5188
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 7156 5188 8677 5216
rect 7156 5176 7162 5188
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 9048 5216 9076 5247
rect 9766 5216 9772 5228
rect 9048 5188 9352 5216
rect 9727 5188 9772 5216
rect 8665 5179 8723 5185
rect 5788 5151 5846 5157
rect 5788 5117 5800 5151
rect 5834 5148 5846 5151
rect 6270 5148 6276 5160
rect 5834 5120 6276 5148
rect 5834 5117 5846 5120
rect 5788 5111 5846 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6822 5108 6828 5160
rect 6880 5148 6886 5160
rect 7650 5148 7656 5160
rect 6880 5120 7656 5148
rect 6880 5108 6886 5120
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7984 5120 8125 5148
rect 7984 5108 7990 5120
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 9214 5148 9220 5160
rect 8536 5120 9220 5148
rect 8536 5108 8542 5120
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9324 5148 9352 5188
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 10192 5188 10609 5216
rect 10192 5176 10198 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10831 5157 10859 5256
rect 11238 5244 11244 5256
rect 11296 5284 11302 5296
rect 13446 5284 13452 5296
rect 11296 5256 13452 5284
rect 11296 5244 11302 5256
rect 13446 5244 13452 5256
rect 13504 5244 13510 5296
rect 9677 5151 9735 5157
rect 9677 5148 9689 5151
rect 9324 5120 9689 5148
rect 9677 5117 9689 5120
rect 9723 5117 9735 5151
rect 9677 5111 9735 5117
rect 10827 5151 10885 5157
rect 10827 5117 10839 5151
rect 10873 5117 10885 5151
rect 10827 5111 10885 5117
rect 11238 5108 11244 5160
rect 11296 5148 11302 5160
rect 12504 5151 12562 5157
rect 12504 5148 12516 5151
rect 11296 5120 12516 5148
rect 11296 5108 11302 5120
rect 12504 5117 12516 5120
rect 12550 5148 12562 5151
rect 12894 5148 12900 5160
rect 12550 5120 12900 5148
rect 12550 5117 12562 5120
rect 12504 5111 12562 5117
rect 12894 5108 12900 5120
rect 12952 5108 12958 5160
rect 8386 5080 8392 5092
rect 8347 5052 8392 5080
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 5859 5015 5917 5021
rect 5859 4981 5871 5015
rect 5905 5012 5917 5015
rect 6086 5012 6092 5024
rect 5905 4984 6092 5012
rect 5905 4981 5917 4984
rect 5859 4975 5917 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 9950 4972 9956 5024
rect 10008 5012 10014 5024
rect 10919 5015 10977 5021
rect 10919 5012 10931 5015
rect 10008 4984 10931 5012
rect 10008 4972 10014 4984
rect 10919 4981 10931 4984
rect 10965 4981 10977 5015
rect 10919 4975 10977 4981
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12575 5015 12633 5021
rect 12575 5012 12587 5015
rect 12492 4984 12587 5012
rect 12492 4972 12498 4984
rect 12575 4981 12587 4984
rect 12621 4981 12633 5015
rect 12575 4975 12633 4981
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 5258 4808 5264 4820
rect 5219 4780 5264 4808
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 7650 4808 7656 4820
rect 7611 4780 7656 4808
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 9214 4808 9220 4820
rect 9175 4780 9220 4808
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 6641 4743 6699 4749
rect 6641 4740 6653 4743
rect 6236 4712 6653 4740
rect 6236 4700 6242 4712
rect 6641 4709 6653 4712
rect 6687 4709 6699 4743
rect 6641 4703 6699 4709
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 9861 4743 9919 4749
rect 6972 4712 8064 4740
rect 6972 4700 6978 4712
rect 5496 4675 5554 4681
rect 5496 4641 5508 4675
rect 5542 4672 5554 4675
rect 5644 4672 5672 4700
rect 8036 4684 8064 4712
rect 9861 4709 9873 4743
rect 9907 4740 9919 4743
rect 10042 4740 10048 4752
rect 9907 4712 10048 4740
rect 9907 4709 9919 4712
rect 9861 4703 9919 4709
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 8018 4672 8024 4684
rect 5542 4644 5672 4672
rect 7931 4644 8024 4672
rect 5542 4641 5554 4644
rect 5496 4635 5554 4641
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 11238 4672 11244 4684
rect 11199 4644 11244 4672
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12308 4644 12357 4672
rect 12308 4632 12314 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 13354 4632 13360 4684
rect 13412 4672 13418 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13412 4644 13461 4672
rect 13412 4632 13418 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 5583 4607 5641 4613
rect 5583 4573 5595 4607
rect 5629 4604 5641 4607
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5629 4576 6009 4604
rect 5629 4573 5641 4576
rect 5583 4567 5641 4573
rect 5997 4573 6009 4576
rect 6043 4604 6055 4607
rect 6549 4607 6607 4613
rect 6549 4604 6561 4607
rect 6043 4576 6561 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6549 4573 6561 4576
rect 6595 4573 6607 4607
rect 8754 4604 8760 4616
rect 8715 4576 8760 4604
rect 6549 4567 6607 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4573 9827 4607
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 9769 4567 9827 4573
rect 7098 4536 7104 4548
rect 7059 4508 7104 4536
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 6273 4471 6331 4477
rect 6273 4468 6285 4471
rect 6236 4440 6285 4468
rect 6236 4428 6242 4440
rect 6273 4437 6285 4440
rect 6319 4437 6331 4471
rect 9784 4468 9812 4567
rect 10134 4564 10140 4576
rect 10192 4604 10198 4616
rect 10502 4604 10508 4616
rect 10192 4576 10508 4604
rect 10192 4564 10198 4576
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 12529 4539 12587 4545
rect 12529 4505 12541 4539
rect 12575 4536 12587 4539
rect 13814 4536 13820 4548
rect 12575 4508 13820 4536
rect 12575 4505 12587 4508
rect 12529 4499 12587 4505
rect 13814 4496 13820 4508
rect 13872 4496 13878 4548
rect 10778 4468 10784 4480
rect 9784 4440 10784 4468
rect 6273 4431 6331 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11425 4471 11483 4477
rect 11425 4437 11437 4471
rect 11471 4468 11483 4471
rect 12158 4468 12164 4480
rect 11471 4440 12164 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 14642 4468 14648 4480
rect 13679 4440 14648 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 7926 4264 7932 4276
rect 7887 4236 7932 4264
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 11238 4264 11244 4276
rect 11199 4236 11244 4264
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 12250 4264 12256 4276
rect 12211 4236 12256 4264
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 13354 4264 13360 4276
rect 13315 4236 13360 4264
rect 13354 4224 13360 4236
rect 13412 4224 13418 4276
rect 10796 4168 11100 4196
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 4948 4100 5089 4128
rect 4948 4088 4954 4100
rect 5077 4097 5089 4100
rect 5123 4128 5135 4131
rect 5718 4128 5724 4140
rect 5123 4100 5724 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 4062 4060 4068 4072
rect 2924 4032 4068 4060
rect 2924 4020 2930 4032
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 4208 4063 4266 4069
rect 4208 4029 4220 4063
rect 4254 4029 4266 4063
rect 5258 4060 5264 4072
rect 5219 4032 5264 4060
rect 4208 4023 4266 4029
rect 4223 3924 4251 4023
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5644 4069 5672 4100
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 7190 4128 7196 4140
rect 6696 4100 7196 4128
rect 6696 4088 6702 4100
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 7800 4100 8217 4128
rect 7800 4088 7806 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 9674 4128 9680 4140
rect 9635 4100 9680 4128
rect 8205 4091 8263 4097
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 5675 4032 5709 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 4295 3995 4353 4001
rect 4295 3961 4307 3995
rect 4341 3992 4353 3995
rect 5074 3992 5080 4004
rect 4341 3964 5080 3992
rect 4341 3961 4353 3964
rect 4295 3955 4353 3961
rect 5074 3952 5080 3964
rect 5132 3952 5138 4004
rect 5902 3992 5908 4004
rect 5863 3964 5908 3992
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 6914 3992 6920 4004
rect 6875 3964 6920 3992
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3961 7067 3995
rect 8220 3992 8248 4091
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 10226 4128 10232 4140
rect 10187 4100 10232 4128
rect 10226 4088 10232 4100
rect 10284 4128 10290 4140
rect 10796 4128 10824 4168
rect 10284 4100 10824 4128
rect 10873 4131 10931 4137
rect 10284 4088 10290 4100
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 10962 4128 10968 4140
rect 10919 4100 10968 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11072 4128 11100 4168
rect 11609 4131 11667 4137
rect 11609 4128 11621 4131
rect 11072 4100 11621 4128
rect 11609 4097 11621 4100
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 8386 4060 8392 4072
rect 8347 4032 8392 4060
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12526 4060 12532 4072
rect 12483 4032 12532 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 12526 4020 12532 4032
rect 12584 4060 12590 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12584 4032 13001 4060
rect 12584 4020 12590 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13538 4020 13544 4072
rect 13596 4069 13602 4072
rect 13596 4063 13634 4069
rect 13622 4060 13634 4063
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13622 4032 14013 4060
rect 13622 4029 13634 4032
rect 13596 4023 13634 4029
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 13596 4020 13602 4023
rect 8710 3995 8768 4001
rect 8710 3992 8722 3995
rect 8220 3964 8722 3992
rect 7009 3955 7067 3961
rect 8710 3961 8722 3964
rect 8756 3961 8768 3995
rect 10321 3995 10379 4001
rect 8710 3955 8768 3961
rect 9508 3964 10180 3992
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 4223 3896 4721 3924
rect 4709 3893 4721 3896
rect 4755 3924 4767 3927
rect 5534 3924 5540 3936
rect 4755 3896 5540 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 6086 3924 6092 3936
rect 5684 3896 6092 3924
rect 5684 3884 5690 3896
rect 6086 3884 6092 3896
rect 6144 3924 6150 3936
rect 6181 3927 6239 3933
rect 6181 3924 6193 3927
rect 6144 3896 6193 3924
rect 6144 3884 6150 3896
rect 6181 3893 6193 3896
rect 6227 3893 6239 3927
rect 6181 3887 6239 3893
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 6730 3924 6736 3936
rect 6687 3896 6736 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 6730 3884 6736 3896
rect 6788 3924 6794 3936
rect 7024 3924 7052 3955
rect 9508 3936 9536 3964
rect 7742 3924 7748 3936
rect 6788 3896 7748 3924
rect 6788 3884 6794 3896
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 9309 3927 9367 3933
rect 9309 3893 9321 3927
rect 9355 3924 9367 3927
rect 9490 3924 9496 3936
rect 9355 3896 9496 3924
rect 9355 3893 9367 3896
rect 9309 3887 9367 3893
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10152 3924 10180 3964
rect 10321 3961 10333 3995
rect 10367 3961 10379 3995
rect 10321 3955 10379 3961
rect 10336 3924 10364 3955
rect 10686 3924 10692 3936
rect 10152 3896 10692 3924
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 12894 3924 12900 3936
rect 12667 3896 12900 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13679 3927 13737 3933
rect 13679 3924 13691 3927
rect 13136 3896 13691 3924
rect 13136 3884 13142 3896
rect 13679 3893 13691 3896
rect 13725 3893 13737 3927
rect 13679 3887 13737 3893
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 8812 3692 9413 3720
rect 8812 3680 8818 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9401 3683 9459 3689
rect 10410 3680 10416 3732
rect 10468 3720 10474 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 10468 3692 11161 3720
rect 10468 3680 10474 3692
rect 11149 3689 11161 3692
rect 11195 3720 11207 3723
rect 12342 3720 12348 3732
rect 11195 3692 12348 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 6270 3661 6276 3664
rect 6267 3652 6276 3661
rect 6183 3624 6276 3652
rect 6267 3615 6276 3624
rect 6328 3652 6334 3664
rect 7650 3652 7656 3664
rect 6328 3624 7656 3652
rect 6270 3612 6276 3615
rect 6328 3612 6334 3624
rect 7650 3612 7656 3624
rect 7708 3652 7714 3664
rect 8018 3652 8024 3664
rect 7708 3624 8024 3652
rect 7708 3612 7714 3624
rect 8018 3612 8024 3624
rect 8076 3652 8082 3664
rect 8158 3655 8216 3661
rect 8158 3652 8170 3655
rect 8076 3624 8170 3652
rect 8076 3612 8082 3624
rect 8158 3621 8170 3624
rect 8204 3621 8216 3655
rect 8158 3615 8216 3621
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 9033 3655 9091 3661
rect 9033 3652 9045 3655
rect 8444 3624 9045 3652
rect 8444 3612 8450 3624
rect 9033 3621 9045 3624
rect 9079 3621 9091 3655
rect 9858 3652 9864 3664
rect 9771 3624 9864 3652
rect 9033 3615 9091 3621
rect 9858 3612 9864 3624
rect 9916 3652 9922 3664
rect 11422 3652 11428 3664
rect 9916 3624 11428 3652
rect 9916 3612 9922 3624
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 4614 3584 4620 3596
rect 4575 3556 4620 3584
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4890 3584 4896 3596
rect 4851 3556 4896 3584
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3584 5135 3587
rect 6822 3584 6828 3596
rect 5123 3556 6828 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 6822 3544 6828 3556
rect 6880 3584 6886 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6880 3556 7113 3584
rect 6880 3544 6886 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7834 3584 7840 3596
rect 7795 3556 7840 3584
rect 7101 3547 7159 3553
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 13446 3584 13452 3596
rect 13407 3556 13452 3584
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 5902 3516 5908 3528
rect 5863 3488 5908 3516
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 9950 3516 9956 3528
rect 9815 3488 9956 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 9950 3476 9956 3488
rect 10008 3516 10014 3528
rect 11054 3516 11060 3528
rect 10008 3488 11060 3516
rect 10008 3476 10014 3488
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11790 3516 11796 3528
rect 11379 3488 11796 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11790 3476 11796 3488
rect 11848 3516 11854 3528
rect 13078 3516 13084 3528
rect 11848 3488 13084 3516
rect 11848 3476 11854 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 6178 3448 6184 3460
rect 5368 3420 6184 3448
rect 5368 3392 5396 3420
rect 6178 3408 6184 3420
rect 6236 3448 6242 3460
rect 6825 3451 6883 3457
rect 6825 3448 6837 3451
rect 6236 3420 6837 3448
rect 6236 3408 6242 3420
rect 6825 3417 6837 3420
rect 6871 3417 6883 3451
rect 6825 3411 6883 3417
rect 8757 3451 8815 3457
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 10042 3448 10048 3460
rect 8803 3420 10048 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 10321 3451 10379 3457
rect 10321 3417 10333 3451
rect 10367 3448 10379 3451
rect 10962 3448 10968 3460
rect 10367 3420 10968 3448
rect 10367 3417 10379 3420
rect 10321 3411 10379 3417
rect 10962 3408 10968 3420
rect 11020 3408 11026 3460
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3417 11943 3451
rect 11885 3411 11943 3417
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 5718 3380 5724 3392
rect 5679 3352 5724 3380
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 7466 3380 7472 3392
rect 7427 3352 7472 3380
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 11900 3380 11928 3411
rect 13630 3380 13636 3392
rect 10560 3352 11928 3380
rect 13591 3352 13636 3380
rect 10560 3340 10566 3352
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 4295 3179 4353 3185
rect 4295 3145 4307 3179
rect 4341 3176 4353 3179
rect 5442 3176 5448 3188
rect 4341 3148 5448 3176
rect 4341 3145 4353 3148
rect 4295 3139 4353 3145
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3176 6334 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6328 3148 6561 3176
rect 6328 3136 6334 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 7742 3176 7748 3188
rect 7703 3148 7748 3176
rect 6549 3139 6607 3145
rect 4065 3111 4123 3117
rect 4065 3077 4077 3111
rect 4111 3108 4123 3111
rect 4614 3108 4620 3120
rect 4111 3080 4620 3108
rect 4111 3077 4123 3080
rect 4065 3071 4123 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 4890 3068 4896 3120
rect 4948 3108 4954 3120
rect 4985 3111 5043 3117
rect 4985 3108 4997 3111
rect 4948 3080 4997 3108
rect 4948 3068 4954 3080
rect 4985 3077 4997 3080
rect 5031 3077 5043 3111
rect 6564 3108 6592 3139
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 8018 3176 8024 3188
rect 7979 3148 8024 3176
rect 8018 3136 8024 3148
rect 8076 3176 8082 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 8076 3148 8401 3176
rect 8076 3136 8082 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 9493 3179 9551 3185
rect 9493 3145 9505 3179
rect 9539 3176 9551 3179
rect 9858 3176 9864 3188
rect 9539 3148 9864 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 6564 3080 7189 3108
rect 4985 3071 5043 3077
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 4488 3012 5273 3040
rect 4488 3000 4494 3012
rect 5261 3009 5273 3012
rect 5307 3040 5319 3043
rect 5718 3040 5724 3052
rect 5307 3012 5724 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 6638 3040 6644 3052
rect 5951 3012 6644 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 3212 2975 3270 2981
rect 3212 2941 3224 2975
rect 3258 2972 3270 2975
rect 3694 2972 3700 2984
rect 3258 2944 3700 2972
rect 3258 2941 3270 2944
rect 3212 2935 3270 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 4208 2975 4266 2981
rect 4208 2941 4220 2975
rect 4254 2972 4266 2975
rect 7161 2972 7189 3080
rect 4254 2941 4267 2972
rect 7161 2944 7230 2972
rect 4208 2935 4267 2941
rect 382 2864 388 2916
rect 440 2904 446 2916
rect 4239 2904 4267 2935
rect 4617 2907 4675 2913
rect 4617 2904 4629 2907
rect 440 2876 4629 2904
rect 440 2864 446 2876
rect 4617 2873 4629 2876
rect 4663 2873 4675 2907
rect 5350 2904 5356 2916
rect 5311 2876 5356 2904
rect 4617 2867 4675 2873
rect 3283 2839 3341 2845
rect 3283 2805 3295 2839
rect 3329 2836 3341 2839
rect 3510 2836 3516 2848
rect 3329 2808 3516 2836
rect 3329 2805 3341 2808
rect 3283 2799 3341 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 4632 2836 4660 2867
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 7202 2913 7230 2944
rect 7187 2907 7245 2913
rect 7187 2873 7199 2907
rect 7233 2873 7245 2907
rect 8404 2904 8432 3139
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 12989 3179 13047 3185
rect 12989 3176 13001 3179
rect 12768 3148 13001 3176
rect 12768 3136 12774 3148
rect 12989 3145 13001 3148
rect 13035 3145 13047 3179
rect 12989 3139 13047 3145
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 13679 3179 13737 3185
rect 13679 3176 13691 3179
rect 13320 3148 13691 3176
rect 13320 3136 13326 3148
rect 13679 3145 13691 3148
rect 13725 3145 13737 3179
rect 13679 3139 13737 3145
rect 10962 3108 10968 3120
rect 10923 3080 10968 3108
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 11388 3080 12633 3108
rect 11388 3068 11394 3080
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 13446 3108 13452 3120
rect 13407 3080 13452 3108
rect 12621 3071 12679 3077
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8754 3040 8760 3052
rect 8619 3012 8760 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 10410 3040 10416 3052
rect 10371 3012 10416 3040
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12710 2972 12716 2984
rect 12483 2944 12716 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 13538 2932 13544 2984
rect 13596 2981 13602 2984
rect 13596 2975 13634 2981
rect 13622 2972 13634 2975
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13622 2944 14013 2972
rect 13622 2941 13634 2944
rect 13596 2935 13634 2941
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 13596 2932 13602 2935
rect 8894 2907 8952 2913
rect 8894 2904 8906 2907
rect 8404 2876 8906 2904
rect 7187 2867 7245 2873
rect 8894 2873 8906 2876
rect 8940 2873 8952 2907
rect 8894 2867 8952 2873
rect 10042 2864 10048 2916
rect 10100 2904 10106 2916
rect 10229 2907 10287 2913
rect 10229 2904 10241 2907
rect 10100 2876 10241 2904
rect 10100 2864 10106 2876
rect 10229 2873 10241 2876
rect 10275 2904 10287 2907
rect 10505 2907 10563 2913
rect 10505 2904 10517 2907
rect 10275 2876 10517 2904
rect 10275 2873 10287 2876
rect 10229 2867 10287 2873
rect 10505 2873 10517 2876
rect 10551 2873 10563 2907
rect 10505 2867 10563 2873
rect 7282 2836 7288 2848
rect 4632 2808 7288 2836
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 4430 2641 4436 2644
rect 4387 2635 4436 2641
rect 4387 2601 4399 2635
rect 4433 2601 4436 2635
rect 4387 2595 4436 2601
rect 4430 2592 4436 2595
rect 4488 2592 4494 2644
rect 5902 2592 5908 2644
rect 5960 2632 5966 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 5960 2604 6285 2632
rect 5960 2592 5966 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 6730 2632 6736 2644
rect 6691 2604 6736 2632
rect 6273 2595 6331 2601
rect 6730 2592 6736 2604
rect 6788 2632 6794 2644
rect 6788 2604 7052 2632
rect 6788 2592 6794 2604
rect 5258 2564 5264 2576
rect 4724 2536 5264 2564
rect 4246 2456 4252 2508
rect 4304 2505 4310 2508
rect 4724 2505 4752 2536
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 5994 2564 6000 2576
rect 5955 2536 6000 2564
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 7024 2564 7052 2604
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7156 2604 7788 2632
rect 7156 2592 7162 2604
rect 7760 2573 7788 2604
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7892 2604 8033 2632
rect 7892 2592 7898 2604
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 8021 2595 8079 2601
rect 9490 2592 9496 2604
rect 9548 2632 9554 2644
rect 9548 2604 9996 2632
rect 9548 2592 9554 2604
rect 9968 2573 9996 2604
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 11112 2604 11161 2632
rect 11112 2592 11118 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 13170 2632 13176 2644
rect 13131 2604 13176 2632
rect 11149 2595 11207 2601
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 7193 2567 7251 2573
rect 7193 2564 7205 2567
rect 7024 2536 7205 2564
rect 7193 2533 7205 2536
rect 7239 2533 7251 2567
rect 7193 2527 7251 2533
rect 7745 2567 7803 2573
rect 7745 2533 7757 2567
rect 7791 2533 7803 2567
rect 7745 2527 7803 2533
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2533 10011 2567
rect 10502 2564 10508 2576
rect 10463 2536 10508 2564
rect 9953 2527 10011 2533
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 4304 2499 4342 2505
rect 4330 2496 4342 2499
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 4330 2468 4721 2496
rect 4330 2465 4342 2468
rect 4304 2459 4342 2465
rect 4709 2465 4721 2468
rect 4755 2465 4767 2499
rect 4709 2459 4767 2465
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5902 2496 5908 2508
rect 5215 2468 5908 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 4304 2456 4310 2459
rect 5902 2456 5908 2468
rect 5960 2456 5966 2508
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8628 2468 9137 2496
rect 8628 2456 8634 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 11238 2456 11244 2508
rect 11296 2496 11302 2508
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 11296 2468 11345 2496
rect 11296 2456 11302 2468
rect 11333 2465 11345 2468
rect 11379 2496 11391 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11379 2468 11897 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13188 2496 13216 2592
rect 12667 2468 13216 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 7098 2428 7104 2440
rect 7011 2400 7104 2428
rect 7098 2388 7104 2400
rect 7156 2428 7162 2440
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 7156 2400 8401 2428
rect 7156 2388 7162 2400
rect 8389 2397 8401 2400
rect 8435 2397 8447 2431
rect 9858 2428 9864 2440
rect 9819 2400 9864 2428
rect 8389 2391 8447 2397
rect 9858 2388 9864 2400
rect 9916 2428 9922 2440
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 9916 2400 10793 2428
rect 9916 2388 9922 2400
rect 10781 2397 10793 2400
rect 10827 2397 10839 2431
rect 10781 2391 10839 2397
rect 8754 2292 8760 2304
rect 8715 2264 8760 2292
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 11514 2292 11520 2304
rect 11475 2264 11520 2292
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 12802 2292 12808 2304
rect 12763 2264 12808 2292
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 3694 688 3700 740
rect 3752 728 3758 740
rect 4982 728 4988 740
rect 3752 700 4988 728
rect 3752 688 3758 700
rect 4982 688 4988 700
rect 5040 688 5046 740
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 8576 37272 8628 37324
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 10968 36907 11020 36916
rect 10968 36873 10977 36907
rect 10977 36873 11011 36907
rect 11011 36873 11020 36907
rect 10968 36864 11020 36873
rect 7196 36524 7248 36576
rect 7288 36524 7340 36576
rect 7564 36524 7616 36576
rect 8576 36703 8628 36712
rect 8576 36669 8585 36703
rect 8585 36669 8619 36703
rect 8619 36669 8628 36703
rect 8576 36660 8628 36669
rect 8392 36524 8444 36576
rect 11152 36524 11204 36576
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 10692 36320 10744 36372
rect 12348 36320 12400 36372
rect 6920 36252 6972 36304
rect 9772 36184 9824 36236
rect 11244 36227 11296 36236
rect 11244 36193 11253 36227
rect 11253 36193 11287 36227
rect 11287 36193 11296 36227
rect 11244 36184 11296 36193
rect 7196 36159 7248 36168
rect 7196 36125 7205 36159
rect 7205 36125 7239 36159
rect 7239 36125 7248 36159
rect 7196 36116 7248 36125
rect 7748 36091 7800 36100
rect 7748 36057 7757 36091
rect 7757 36057 7791 36091
rect 7791 36057 7800 36091
rect 7748 36048 7800 36057
rect 8576 35980 8628 36032
rect 9588 35980 9640 36032
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 7196 35776 7248 35828
rect 11336 35776 11388 35828
rect 12072 35776 12124 35828
rect 13728 35776 13780 35828
rect 7748 35751 7800 35760
rect 7748 35717 7757 35751
rect 7757 35717 7791 35751
rect 7791 35717 7800 35751
rect 7748 35708 7800 35717
rect 6920 35640 6972 35692
rect 7012 35504 7064 35556
rect 6736 35436 6788 35488
rect 7472 35436 7524 35488
rect 9496 35572 9548 35624
rect 10232 35615 10284 35624
rect 10232 35581 10241 35615
rect 10241 35581 10275 35615
rect 10275 35581 10284 35615
rect 10232 35572 10284 35581
rect 8760 35479 8812 35488
rect 8760 35445 8769 35479
rect 8769 35445 8803 35479
rect 8803 35445 8812 35479
rect 8760 35436 8812 35445
rect 9772 35479 9824 35488
rect 9772 35445 9781 35479
rect 9781 35445 9815 35479
rect 9815 35445 9824 35479
rect 9772 35436 9824 35445
rect 11336 35436 11388 35488
rect 11980 35436 12032 35488
rect 12992 35479 13044 35488
rect 12992 35445 13001 35479
rect 13001 35445 13035 35479
rect 13035 35445 13044 35479
rect 12992 35436 13044 35445
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 6920 35232 6972 35284
rect 12072 35232 12124 35284
rect 14188 35232 14240 35284
rect 7012 35207 7064 35216
rect 7012 35173 7021 35207
rect 7021 35173 7055 35207
rect 7055 35173 7064 35207
rect 7012 35164 7064 35173
rect 9864 35164 9916 35216
rect 6276 35096 6328 35148
rect 8300 35096 8352 35148
rect 11244 35096 11296 35148
rect 12440 35096 12492 35148
rect 7932 35028 7984 35080
rect 9404 35028 9456 35080
rect 11060 35028 11112 35080
rect 5264 34935 5316 34944
rect 5264 34901 5273 34935
rect 5273 34901 5307 34935
rect 5307 34901 5316 34935
rect 5264 34892 5316 34901
rect 10968 34892 11020 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 5448 34688 5500 34740
rect 6276 34731 6328 34740
rect 6276 34697 6285 34731
rect 6285 34697 6319 34731
rect 6319 34697 6328 34731
rect 6276 34688 6328 34697
rect 7012 34688 7064 34740
rect 8300 34688 8352 34740
rect 8484 34731 8536 34740
rect 8484 34697 8493 34731
rect 8493 34697 8527 34731
rect 8527 34697 8536 34731
rect 8484 34688 8536 34697
rect 13636 34731 13688 34740
rect 13636 34697 13645 34731
rect 13645 34697 13679 34731
rect 13679 34697 13688 34731
rect 13636 34688 13688 34697
rect 8760 34552 8812 34604
rect 10968 34620 11020 34672
rect 10876 34595 10928 34604
rect 10876 34561 10885 34595
rect 10885 34561 10919 34595
rect 10919 34561 10928 34595
rect 10876 34552 10928 34561
rect 12348 34552 12400 34604
rect 4160 34527 4212 34536
rect 4160 34493 4204 34527
rect 4204 34493 4212 34527
rect 4160 34484 4212 34493
rect 5172 34527 5224 34536
rect 5172 34493 5181 34527
rect 5181 34493 5215 34527
rect 5215 34493 5224 34527
rect 5172 34484 5224 34493
rect 5264 34484 5316 34536
rect 5632 34527 5684 34536
rect 5632 34493 5641 34527
rect 5641 34493 5675 34527
rect 5675 34493 5684 34527
rect 5632 34484 5684 34493
rect 6828 34527 6880 34536
rect 6828 34493 6837 34527
rect 6837 34493 6871 34527
rect 6871 34493 6880 34527
rect 6828 34484 6880 34493
rect 9864 34527 9916 34536
rect 9864 34493 9873 34527
rect 9873 34493 9907 34527
rect 9907 34493 9916 34527
rect 9864 34484 9916 34493
rect 11244 34484 11296 34536
rect 12440 34527 12492 34536
rect 12440 34493 12484 34527
rect 12484 34493 12492 34527
rect 12440 34484 12492 34493
rect 13912 34484 13964 34536
rect 6184 34348 6236 34400
rect 9036 34459 9088 34468
rect 9036 34425 9039 34459
rect 9039 34425 9073 34459
rect 9073 34425 9088 34459
rect 9036 34416 9088 34425
rect 10324 34391 10376 34400
rect 10324 34357 10333 34391
rect 10333 34357 10367 34391
rect 10367 34357 10376 34391
rect 10324 34348 10376 34357
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 6920 34144 6972 34196
rect 9404 34187 9456 34196
rect 9404 34153 9413 34187
rect 9413 34153 9447 34187
rect 9447 34153 9456 34187
rect 9404 34144 9456 34153
rect 13544 34187 13596 34196
rect 6184 34119 6236 34128
rect 6184 34085 6187 34119
rect 6187 34085 6221 34119
rect 6221 34085 6236 34119
rect 6184 34076 6236 34085
rect 7012 34119 7064 34128
rect 7012 34085 7021 34119
rect 7021 34085 7055 34119
rect 7055 34085 7064 34119
rect 7012 34076 7064 34085
rect 4528 34008 4580 34060
rect 6736 34051 6788 34060
rect 6736 34017 6745 34051
rect 6745 34017 6779 34051
rect 6779 34017 6788 34051
rect 7840 34076 7892 34128
rect 6736 34008 6788 34017
rect 5908 33940 5960 33992
rect 7932 33983 7984 33992
rect 7932 33949 7941 33983
rect 7941 33949 7975 33983
rect 7975 33949 7984 33983
rect 7932 33940 7984 33949
rect 8300 33872 8352 33924
rect 5264 33847 5316 33856
rect 5264 33813 5273 33847
rect 5273 33813 5307 33847
rect 5307 33813 5316 33847
rect 5264 33804 5316 33813
rect 5540 33804 5592 33856
rect 8208 33804 8260 33856
rect 9036 34076 9088 34128
rect 10140 34076 10192 34128
rect 11060 34076 11112 34128
rect 11520 34119 11572 34128
rect 11520 34085 11529 34119
rect 11529 34085 11563 34119
rect 11563 34085 11572 34119
rect 11520 34076 11572 34085
rect 13544 34153 13553 34187
rect 13553 34153 13587 34187
rect 13587 34153 13596 34187
rect 13544 34144 13596 34153
rect 11704 34076 11756 34128
rect 13544 34008 13596 34060
rect 9680 33983 9732 33992
rect 9680 33949 9689 33983
rect 9689 33949 9723 33983
rect 9723 33949 9732 33983
rect 9680 33940 9732 33949
rect 11980 33983 12032 33992
rect 11980 33949 11989 33983
rect 11989 33949 12023 33983
rect 12023 33949 12032 33983
rect 11980 33940 12032 33949
rect 10508 33804 10560 33856
rect 12532 33847 12584 33856
rect 12532 33813 12541 33847
rect 12541 33813 12575 33847
rect 12575 33813 12584 33847
rect 12532 33804 12584 33813
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 4528 33600 4580 33652
rect 5356 33600 5408 33652
rect 7840 33643 7892 33652
rect 7840 33609 7849 33643
rect 7849 33609 7883 33643
rect 7883 33609 7892 33643
rect 7840 33600 7892 33609
rect 8392 33600 8444 33652
rect 10140 33600 10192 33652
rect 11704 33643 11756 33652
rect 11704 33609 11713 33643
rect 11713 33609 11747 33643
rect 11747 33609 11756 33643
rect 11704 33600 11756 33609
rect 5908 33507 5960 33516
rect 5908 33473 5917 33507
rect 5917 33473 5951 33507
rect 5951 33473 5960 33507
rect 5908 33464 5960 33473
rect 7932 33464 7984 33516
rect 10324 33532 10376 33584
rect 10508 33507 10560 33516
rect 10508 33473 10517 33507
rect 10517 33473 10551 33507
rect 10551 33473 10560 33507
rect 10508 33464 10560 33473
rect 4068 33439 4120 33448
rect 4068 33405 4077 33439
rect 4077 33405 4111 33439
rect 4111 33405 4120 33439
rect 4068 33396 4120 33405
rect 5264 33439 5316 33448
rect 5264 33405 5273 33439
rect 5273 33405 5307 33439
rect 5307 33405 5316 33439
rect 5264 33396 5316 33405
rect 5632 33439 5684 33448
rect 5632 33405 5641 33439
rect 5641 33405 5675 33439
rect 5675 33405 5684 33439
rect 5632 33396 5684 33405
rect 5172 33328 5224 33380
rect 5540 33328 5592 33380
rect 7012 33371 7064 33380
rect 7012 33337 7021 33371
rect 7021 33337 7055 33371
rect 7055 33337 7064 33371
rect 7012 33328 7064 33337
rect 10140 33328 10192 33380
rect 3884 33303 3936 33312
rect 3884 33269 3893 33303
rect 3893 33269 3927 33303
rect 3927 33269 3936 33303
rect 3884 33260 3936 33269
rect 6184 33303 6236 33312
rect 6184 33269 6193 33303
rect 6193 33269 6227 33303
rect 6227 33269 6236 33303
rect 6184 33260 6236 33269
rect 11428 33303 11480 33312
rect 11428 33269 11437 33303
rect 11437 33269 11471 33303
rect 11471 33269 11480 33303
rect 11428 33260 11480 33269
rect 12256 33464 12308 33516
rect 12256 33328 12308 33380
rect 12532 33371 12584 33380
rect 12532 33337 12541 33371
rect 12541 33337 12575 33371
rect 12575 33337 12584 33371
rect 12532 33328 12584 33337
rect 13544 33303 13596 33312
rect 13544 33269 13553 33303
rect 13553 33269 13587 33303
rect 13587 33269 13596 33303
rect 13544 33260 13596 33269
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 4068 33056 4120 33108
rect 5448 33056 5500 33108
rect 5632 33099 5684 33108
rect 5632 33065 5641 33099
rect 5641 33065 5675 33099
rect 5675 33065 5684 33099
rect 5632 33056 5684 33065
rect 8300 33056 8352 33108
rect 9680 33056 9732 33108
rect 11520 33099 11572 33108
rect 11520 33065 11529 33099
rect 11529 33065 11563 33099
rect 11563 33065 11572 33099
rect 11520 33056 11572 33065
rect 6184 32988 6236 33040
rect 8024 33031 8076 33040
rect 8024 32997 8033 33031
rect 8033 32997 8067 33031
rect 8067 32997 8076 33031
rect 8024 32988 8076 32997
rect 10324 33031 10376 33040
rect 10324 32997 10333 33031
rect 10333 32997 10367 33031
rect 10367 32997 10376 33031
rect 10324 32988 10376 32997
rect 10876 33031 10928 33040
rect 10876 32997 10885 33031
rect 10885 32997 10919 33031
rect 10919 32997 10928 33031
rect 10876 32988 10928 32997
rect 12348 33056 12400 33108
rect 11888 33031 11940 33040
rect 11888 32997 11897 33031
rect 11897 32997 11931 33031
rect 11931 32997 11940 33031
rect 11888 32988 11940 32997
rect 4344 32920 4396 32972
rect 4988 32920 5040 32972
rect 13544 32920 13596 32972
rect 6092 32852 6144 32904
rect 7748 32852 7800 32904
rect 8300 32895 8352 32904
rect 8300 32861 8309 32895
rect 8309 32861 8343 32895
rect 8343 32861 8352 32895
rect 8300 32852 8352 32861
rect 9588 32852 9640 32904
rect 11520 32852 11572 32904
rect 12164 32852 12216 32904
rect 5172 32759 5224 32768
rect 5172 32725 5181 32759
rect 5181 32725 5215 32759
rect 5215 32725 5224 32759
rect 5172 32716 5224 32725
rect 7012 32759 7064 32768
rect 7012 32725 7021 32759
rect 7021 32725 7055 32759
rect 7055 32725 7064 32759
rect 7012 32716 7064 32725
rect 7380 32759 7432 32768
rect 7380 32725 7389 32759
rect 7389 32725 7423 32759
rect 7423 32725 7432 32759
rect 7380 32716 7432 32725
rect 12900 32716 12952 32768
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 4988 32555 5040 32564
rect 4988 32521 4997 32555
rect 4997 32521 5031 32555
rect 5031 32521 5040 32555
rect 4988 32512 5040 32521
rect 8024 32512 8076 32564
rect 10324 32512 10376 32564
rect 11428 32512 11480 32564
rect 11888 32512 11940 32564
rect 12348 32512 12400 32564
rect 12624 32512 12676 32564
rect 10048 32419 10100 32428
rect 10048 32385 10057 32419
rect 10057 32385 10091 32419
rect 10091 32385 10100 32419
rect 10048 32376 10100 32385
rect 10876 32376 10928 32428
rect 4528 32308 4580 32360
rect 5172 32351 5224 32360
rect 5172 32317 5181 32351
rect 5181 32317 5215 32351
rect 5215 32317 5224 32351
rect 5172 32308 5224 32317
rect 5632 32351 5684 32360
rect 5632 32317 5641 32351
rect 5641 32317 5675 32351
rect 5675 32317 5684 32351
rect 5632 32308 5684 32317
rect 6000 32308 6052 32360
rect 7380 32351 7432 32360
rect 7380 32317 7389 32351
rect 7389 32317 7423 32351
rect 7423 32317 7432 32351
rect 7380 32308 7432 32317
rect 12440 32351 12492 32360
rect 12440 32317 12484 32351
rect 12484 32317 12492 32351
rect 12440 32308 12492 32317
rect 6092 32240 6144 32292
rect 5540 32172 5592 32224
rect 6184 32172 6236 32224
rect 7104 32172 7156 32224
rect 8208 32240 8260 32292
rect 9864 32283 9916 32292
rect 9864 32249 9873 32283
rect 9873 32249 9907 32283
rect 9907 32249 9916 32283
rect 9864 32240 9916 32249
rect 9588 32172 9640 32224
rect 13544 32172 13596 32224
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 6092 31968 6144 32020
rect 6000 31943 6052 31952
rect 6000 31909 6009 31943
rect 6009 31909 6043 31943
rect 6043 31909 6052 31943
rect 6000 31900 6052 31909
rect 7012 31943 7064 31952
rect 7012 31909 7021 31943
rect 7021 31909 7055 31943
rect 7055 31909 7064 31943
rect 7012 31900 7064 31909
rect 7748 31968 7800 32020
rect 7932 31968 7984 32020
rect 9588 31968 9640 32020
rect 9680 31968 9732 32020
rect 12256 31968 12308 32020
rect 4068 31875 4120 31884
rect 4068 31841 4112 31875
rect 4112 31841 4120 31875
rect 5448 31875 5500 31884
rect 4068 31832 4120 31841
rect 5448 31841 5457 31875
rect 5457 31841 5491 31875
rect 5491 31841 5500 31875
rect 5448 31832 5500 31841
rect 5632 31832 5684 31884
rect 8760 31832 8812 31884
rect 9956 31875 10008 31884
rect 9956 31841 9965 31875
rect 9965 31841 9999 31875
rect 9999 31841 10008 31875
rect 9956 31832 10008 31841
rect 4252 31764 4304 31816
rect 11152 31832 11204 31884
rect 12164 31832 12216 31884
rect 5540 31696 5592 31748
rect 6552 31696 6604 31748
rect 9496 31628 9548 31680
rect 10600 31628 10652 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 5724 31467 5776 31476
rect 5724 31433 5733 31467
rect 5733 31433 5767 31467
rect 5767 31433 5776 31467
rect 5724 31424 5776 31433
rect 6552 31467 6604 31476
rect 6552 31433 6561 31467
rect 6561 31433 6595 31467
rect 6595 31433 6604 31467
rect 6552 31424 6604 31433
rect 7012 31467 7064 31476
rect 7012 31433 7021 31467
rect 7021 31433 7055 31467
rect 7055 31433 7064 31467
rect 7012 31424 7064 31433
rect 8300 31356 8352 31408
rect 7932 31288 7984 31340
rect 9588 31331 9640 31340
rect 9588 31297 9597 31331
rect 9597 31297 9631 31331
rect 9631 31297 9640 31331
rect 9588 31288 9640 31297
rect 10784 31331 10836 31340
rect 10784 31297 10793 31331
rect 10793 31297 10827 31331
rect 10827 31297 10836 31331
rect 10784 31288 10836 31297
rect 11980 31288 12032 31340
rect 5172 31263 5224 31272
rect 5172 31229 5181 31263
rect 5181 31229 5215 31263
rect 5215 31229 5224 31263
rect 5172 31220 5224 31229
rect 9036 31263 9088 31272
rect 9036 31229 9045 31263
rect 9045 31229 9079 31263
rect 9079 31229 9088 31263
rect 9036 31220 9088 31229
rect 9496 31263 9548 31272
rect 9496 31229 9505 31263
rect 9505 31229 9539 31263
rect 9539 31229 9548 31263
rect 9496 31220 9548 31229
rect 4068 31152 4120 31204
rect 5356 31152 5408 31204
rect 7748 31152 7800 31204
rect 9956 31152 10008 31204
rect 10600 31152 10652 31204
rect 4896 31127 4948 31136
rect 4896 31093 4905 31127
rect 4905 31093 4939 31127
rect 4939 31093 4948 31127
rect 4896 31084 4948 31093
rect 5448 31084 5500 31136
rect 6092 31127 6144 31136
rect 6092 31093 6101 31127
rect 6101 31093 6135 31127
rect 6135 31093 6144 31127
rect 6092 31084 6144 31093
rect 8760 31084 8812 31136
rect 9772 31084 9824 31136
rect 12164 31084 12216 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 7012 30880 7064 30932
rect 9036 30923 9088 30932
rect 9036 30889 9045 30923
rect 9045 30889 9079 30923
rect 9079 30889 9088 30923
rect 9036 30880 9088 30889
rect 10600 30923 10652 30932
rect 10600 30889 10609 30923
rect 10609 30889 10643 30923
rect 10643 30889 10652 30923
rect 10600 30880 10652 30889
rect 10784 30880 10836 30932
rect 4896 30812 4948 30864
rect 7840 30855 7892 30864
rect 7840 30821 7849 30855
rect 7849 30821 7883 30855
rect 7883 30821 7892 30855
rect 7840 30812 7892 30821
rect 10140 30812 10192 30864
rect 11612 30855 11664 30864
rect 11612 30821 11621 30855
rect 11621 30821 11655 30855
rect 11655 30821 11664 30855
rect 11612 30812 11664 30821
rect 5632 30744 5684 30796
rect 5816 30744 5868 30796
rect 6184 30744 6236 30796
rect 6460 30787 6512 30796
rect 6460 30753 6469 30787
rect 6469 30753 6503 30787
rect 6503 30753 6512 30787
rect 6460 30744 6512 30753
rect 4068 30676 4120 30728
rect 5356 30719 5408 30728
rect 5356 30685 5365 30719
rect 5365 30685 5399 30719
rect 5399 30685 5408 30719
rect 5356 30676 5408 30685
rect 8024 30676 8076 30728
rect 9680 30719 9732 30728
rect 9680 30685 9689 30719
rect 9689 30685 9723 30719
rect 9723 30685 9732 30719
rect 9680 30676 9732 30685
rect 11520 30719 11572 30728
rect 11520 30685 11529 30719
rect 11529 30685 11563 30719
rect 11563 30685 11572 30719
rect 11520 30676 11572 30685
rect 11980 30719 12032 30728
rect 11980 30685 11989 30719
rect 11989 30685 12023 30719
rect 12023 30685 12032 30719
rect 11980 30676 12032 30685
rect 5448 30608 5500 30660
rect 8300 30651 8352 30660
rect 5172 30540 5224 30592
rect 5908 30540 5960 30592
rect 8300 30617 8309 30651
rect 8309 30617 8343 30651
rect 8343 30617 8352 30651
rect 8300 30608 8352 30617
rect 7104 30583 7156 30592
rect 7104 30549 7113 30583
rect 7113 30549 7147 30583
rect 7147 30549 7156 30583
rect 7104 30540 7156 30549
rect 7748 30540 7800 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 4896 30336 4948 30388
rect 6460 30336 6512 30388
rect 7748 30379 7800 30388
rect 7748 30345 7757 30379
rect 7757 30345 7791 30379
rect 7791 30345 7800 30379
rect 7748 30336 7800 30345
rect 8024 30379 8076 30388
rect 8024 30345 8033 30379
rect 8033 30345 8067 30379
rect 8067 30345 8076 30379
rect 8024 30336 8076 30345
rect 11520 30379 11572 30388
rect 11520 30345 11529 30379
rect 11529 30345 11563 30379
rect 11563 30345 11572 30379
rect 11520 30336 11572 30345
rect 4068 30268 4120 30320
rect 8852 30268 8904 30320
rect 11612 30268 11664 30320
rect 5356 30243 5408 30252
rect 5356 30209 5365 30243
rect 5365 30209 5399 30243
rect 5399 30209 5408 30243
rect 5356 30200 5408 30209
rect 9588 30200 9640 30252
rect 6828 30175 6880 30184
rect 6828 30141 6837 30175
rect 6837 30141 6871 30175
rect 6871 30141 6880 30175
rect 6828 30132 6880 30141
rect 8300 30132 8352 30184
rect 5080 30107 5132 30116
rect 5080 30073 5089 30107
rect 5089 30073 5123 30107
rect 5123 30073 5132 30107
rect 5080 30064 5132 30073
rect 5172 30107 5224 30116
rect 5172 30073 5181 30107
rect 5181 30073 5215 30107
rect 5215 30073 5224 30107
rect 5172 30064 5224 30073
rect 7104 30064 7156 30116
rect 8392 30039 8444 30048
rect 8392 30005 8401 30039
rect 8401 30005 8435 30039
rect 8435 30005 8444 30039
rect 8392 29996 8444 30005
rect 9680 29996 9732 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 5080 29792 5132 29844
rect 5356 29792 5408 29844
rect 7840 29835 7892 29844
rect 7840 29801 7849 29835
rect 7849 29801 7883 29835
rect 7883 29801 7892 29835
rect 7840 29792 7892 29801
rect 8024 29792 8076 29844
rect 9588 29792 9640 29844
rect 11520 29792 11572 29844
rect 4804 29724 4856 29776
rect 6552 29724 6604 29776
rect 7104 29724 7156 29776
rect 10048 29724 10100 29776
rect 10692 29724 10744 29776
rect 3056 29699 3108 29708
rect 3056 29665 3074 29699
rect 3074 29665 3108 29699
rect 3056 29656 3108 29665
rect 12348 29699 12400 29708
rect 12348 29665 12366 29699
rect 12366 29665 12400 29699
rect 12348 29656 12400 29665
rect 4804 29631 4856 29640
rect 4804 29597 4813 29631
rect 4813 29597 4847 29631
rect 4847 29597 4856 29631
rect 4804 29588 4856 29597
rect 6184 29588 6236 29640
rect 7380 29588 7432 29640
rect 9956 29588 10008 29640
rect 10784 29588 10836 29640
rect 5356 29563 5408 29572
rect 4436 29452 4488 29504
rect 5356 29529 5365 29563
rect 5365 29529 5399 29563
rect 5399 29529 5408 29563
rect 5356 29520 5408 29529
rect 6368 29495 6420 29504
rect 6368 29461 6377 29495
rect 6377 29461 6411 29495
rect 6411 29461 6420 29495
rect 6368 29452 6420 29461
rect 10968 29452 11020 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 11060 29248 11112 29300
rect 12348 29248 12400 29300
rect 12992 29291 13044 29300
rect 12992 29257 13001 29291
rect 13001 29257 13035 29291
rect 13035 29257 13044 29291
rect 12992 29248 13044 29257
rect 5172 29180 5224 29232
rect 6552 29223 6604 29232
rect 6552 29189 6561 29223
rect 6561 29189 6595 29223
rect 6595 29189 6604 29223
rect 6552 29180 6604 29189
rect 4436 29112 4488 29164
rect 5356 29155 5408 29164
rect 5356 29121 5365 29155
rect 5365 29121 5399 29155
rect 5399 29121 5408 29155
rect 5356 29112 5408 29121
rect 7380 29155 7432 29164
rect 7380 29121 7389 29155
rect 7389 29121 7423 29155
rect 7423 29121 7432 29155
rect 7380 29112 7432 29121
rect 3516 29044 3568 29096
rect 4252 29044 4304 29096
rect 7012 29087 7064 29096
rect 7012 29053 7021 29087
rect 7021 29053 7055 29087
rect 7055 29053 7064 29087
rect 7012 29044 7064 29053
rect 7288 29087 7340 29096
rect 7288 29053 7297 29087
rect 7297 29053 7331 29087
rect 7331 29053 7340 29087
rect 7288 29044 7340 29053
rect 3056 29019 3108 29028
rect 3056 28985 3065 29019
rect 3065 28985 3099 29019
rect 3099 28985 3108 29019
rect 3056 28976 3108 28985
rect 4804 28976 4856 29028
rect 4712 28951 4764 28960
rect 4712 28917 4721 28951
rect 4721 28917 4755 28951
rect 4755 28917 4764 28951
rect 4712 28908 4764 28917
rect 4896 28908 4948 28960
rect 6368 28976 6420 29028
rect 8300 28976 8352 29028
rect 10968 29180 11020 29232
rect 10876 29155 10928 29164
rect 10876 29121 10885 29155
rect 10885 29121 10919 29155
rect 10919 29121 10928 29155
rect 10876 29112 10928 29121
rect 5540 28908 5592 28960
rect 8392 28951 8444 28960
rect 8392 28917 8401 28951
rect 8401 28917 8435 28951
rect 8435 28917 8444 28951
rect 10048 28976 10100 29028
rect 12440 29087 12492 29096
rect 12440 29053 12449 29087
rect 12449 29053 12483 29087
rect 12483 29053 12492 29087
rect 12440 29044 12492 29053
rect 13452 29087 13504 29096
rect 13452 29053 13496 29087
rect 13496 29053 13504 29087
rect 13452 29044 13504 29053
rect 11060 28976 11112 29028
rect 12992 28976 13044 29028
rect 8392 28908 8444 28917
rect 9772 28908 9824 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 4804 28704 4856 28756
rect 5724 28704 5776 28756
rect 6184 28747 6236 28756
rect 6184 28713 6193 28747
rect 6193 28713 6227 28747
rect 6227 28713 6236 28747
rect 6184 28704 6236 28713
rect 9956 28747 10008 28756
rect 9956 28713 9965 28747
rect 9965 28713 9999 28747
rect 9999 28713 10008 28747
rect 9956 28704 10008 28713
rect 11244 28704 11296 28756
rect 4712 28679 4764 28688
rect 4712 28645 4721 28679
rect 4721 28645 4755 28679
rect 4755 28645 4764 28679
rect 4712 28636 4764 28645
rect 7288 28679 7340 28688
rect 7288 28645 7297 28679
rect 7297 28645 7331 28679
rect 7331 28645 7340 28679
rect 7288 28636 7340 28645
rect 9588 28636 9640 28688
rect 11152 28636 11204 28688
rect 4804 28611 4856 28620
rect 4804 28577 4813 28611
rect 4813 28577 4847 28611
rect 4847 28577 4856 28611
rect 4804 28568 4856 28577
rect 6552 28611 6604 28620
rect 6552 28577 6561 28611
rect 6561 28577 6595 28611
rect 6595 28577 6604 28611
rect 6552 28568 6604 28577
rect 6736 28611 6788 28620
rect 6736 28577 6745 28611
rect 6745 28577 6779 28611
rect 6779 28577 6788 28611
rect 6736 28568 6788 28577
rect 8024 28611 8076 28620
rect 8024 28577 8033 28611
rect 8033 28577 8067 28611
rect 8067 28577 8076 28611
rect 8024 28568 8076 28577
rect 9772 28568 9824 28620
rect 10876 28611 10928 28620
rect 10876 28577 10885 28611
rect 10885 28577 10919 28611
rect 10919 28577 10928 28611
rect 10876 28568 10928 28577
rect 13636 28568 13688 28620
rect 6828 28543 6880 28552
rect 6828 28509 6837 28543
rect 6837 28509 6871 28543
rect 6871 28509 6880 28543
rect 6828 28500 6880 28509
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 12532 28500 12584 28552
rect 10784 28432 10836 28484
rect 12348 28475 12400 28484
rect 12348 28441 12357 28475
rect 12357 28441 12391 28475
rect 12391 28441 12400 28475
rect 12348 28432 12400 28441
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 4804 28160 4856 28212
rect 9772 28203 9824 28212
rect 9772 28169 9781 28203
rect 9781 28169 9815 28203
rect 9815 28169 9824 28203
rect 9772 28160 9824 28169
rect 11152 28203 11204 28212
rect 11152 28169 11161 28203
rect 11161 28169 11195 28203
rect 11195 28169 11204 28203
rect 11152 28160 11204 28169
rect 13636 28203 13688 28212
rect 13636 28169 13645 28203
rect 13645 28169 13679 28203
rect 13679 28169 13688 28203
rect 13636 28160 13688 28169
rect 3516 27820 3568 27872
rect 3884 27956 3936 28008
rect 8668 28092 8720 28144
rect 10968 28092 11020 28144
rect 13176 28092 13228 28144
rect 4896 28067 4948 28076
rect 4896 28033 4905 28067
rect 4905 28033 4939 28067
rect 4939 28033 4948 28067
rect 4896 28024 4948 28033
rect 5172 28024 5224 28076
rect 6552 28024 6604 28076
rect 6828 28024 6880 28076
rect 8024 28024 8076 28076
rect 11980 28024 12032 28076
rect 4988 27999 5040 28008
rect 4988 27965 4997 27999
rect 4997 27965 5031 27999
rect 5031 27965 5040 27999
rect 4988 27956 5040 27965
rect 7288 27956 7340 28008
rect 8944 27956 8996 28008
rect 9680 27956 9732 28008
rect 7472 27888 7524 27940
rect 8392 27931 8444 27940
rect 8392 27897 8401 27931
rect 8401 27897 8435 27931
rect 8435 27897 8444 27931
rect 8392 27888 8444 27897
rect 9772 27888 9824 27940
rect 5540 27820 5592 27872
rect 6828 27820 6880 27872
rect 7656 27820 7708 27872
rect 9404 27863 9456 27872
rect 9404 27829 9413 27863
rect 9413 27829 9447 27863
rect 9447 27829 9456 27863
rect 9404 27820 9456 27829
rect 10140 27820 10192 27872
rect 10324 27820 10376 27872
rect 11428 27820 11480 27872
rect 12716 27863 12768 27872
rect 12716 27829 12725 27863
rect 12725 27829 12759 27863
rect 12759 27829 12768 27863
rect 12716 27820 12768 27829
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 3516 27659 3568 27668
rect 3516 27625 3525 27659
rect 3525 27625 3559 27659
rect 3559 27625 3568 27659
rect 3516 27616 3568 27625
rect 4988 27616 5040 27668
rect 6736 27616 6788 27668
rect 8944 27659 8996 27668
rect 8944 27625 8953 27659
rect 8953 27625 8987 27659
rect 8987 27625 8996 27659
rect 8944 27616 8996 27625
rect 9404 27616 9456 27668
rect 5448 27548 5500 27600
rect 7288 27548 7340 27600
rect 9680 27616 9732 27668
rect 12532 27659 12584 27668
rect 12532 27625 12541 27659
rect 12541 27625 12575 27659
rect 12575 27625 12584 27659
rect 12532 27616 12584 27625
rect 13176 27616 13228 27668
rect 10048 27548 10100 27600
rect 10876 27548 10928 27600
rect 4160 27523 4212 27532
rect 4160 27489 4169 27523
rect 4169 27489 4203 27523
rect 4203 27489 4212 27523
rect 4160 27480 4212 27489
rect 4896 27480 4948 27532
rect 5172 27523 5224 27532
rect 5172 27489 5181 27523
rect 5181 27489 5215 27523
rect 5215 27489 5224 27523
rect 5172 27480 5224 27489
rect 6000 27523 6052 27532
rect 6000 27489 6009 27523
rect 6009 27489 6043 27523
rect 6043 27489 6052 27523
rect 6000 27480 6052 27489
rect 7380 27480 7432 27532
rect 7564 27480 7616 27532
rect 8392 27523 8444 27532
rect 8392 27489 8401 27523
rect 8401 27489 8435 27523
rect 8435 27489 8444 27523
rect 8392 27480 8444 27489
rect 11060 27480 11112 27532
rect 11612 27548 11664 27600
rect 12348 27548 12400 27600
rect 13084 27523 13136 27532
rect 13084 27489 13128 27523
rect 13128 27489 13136 27523
rect 13084 27480 13136 27489
rect 6184 27412 6236 27464
rect 8300 27412 8352 27464
rect 10140 27412 10192 27464
rect 10692 27412 10744 27464
rect 11520 27344 11572 27396
rect 9496 27319 9548 27328
rect 9496 27285 9505 27319
rect 9505 27285 9539 27319
rect 9539 27285 9548 27319
rect 9496 27276 9548 27285
rect 11336 27276 11388 27328
rect 12164 27276 12216 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 4160 27115 4212 27124
rect 4160 27081 4169 27115
rect 4169 27081 4203 27115
rect 4203 27081 4212 27115
rect 4160 27072 4212 27081
rect 5908 27115 5960 27124
rect 5908 27081 5917 27115
rect 5917 27081 5951 27115
rect 5951 27081 5960 27115
rect 5908 27072 5960 27081
rect 6184 27115 6236 27124
rect 6184 27081 6193 27115
rect 6193 27081 6227 27115
rect 6227 27081 6236 27115
rect 6184 27072 6236 27081
rect 6736 27072 6788 27124
rect 10048 27115 10100 27124
rect 10048 27081 10057 27115
rect 10057 27081 10091 27115
rect 10091 27081 10100 27115
rect 10048 27072 10100 27081
rect 11612 27115 11664 27124
rect 11612 27081 11621 27115
rect 11621 27081 11655 27115
rect 11655 27081 11664 27115
rect 11612 27072 11664 27081
rect 12440 27072 12492 27124
rect 13084 27115 13136 27124
rect 13084 27081 13093 27115
rect 13093 27081 13127 27115
rect 13127 27081 13136 27115
rect 13084 27072 13136 27081
rect 5264 27004 5316 27056
rect 4988 26911 5040 26920
rect 4988 26877 4997 26911
rect 4997 26877 5031 26911
rect 5031 26877 5040 26911
rect 4988 26868 5040 26877
rect 4804 26800 4856 26852
rect 6092 26800 6144 26852
rect 9680 26936 9732 26988
rect 10876 26936 10928 26988
rect 7932 26911 7984 26920
rect 7932 26877 7941 26911
rect 7941 26877 7975 26911
rect 7975 26877 7984 26911
rect 7932 26868 7984 26877
rect 8392 26868 8444 26920
rect 11428 26868 11480 26920
rect 10600 26843 10652 26852
rect 10600 26809 10609 26843
rect 10609 26809 10643 26843
rect 10643 26809 10652 26843
rect 10600 26800 10652 26809
rect 11244 26800 11296 26852
rect 4712 26732 4764 26784
rect 6000 26732 6052 26784
rect 7104 26732 7156 26784
rect 7380 26775 7432 26784
rect 7380 26741 7389 26775
rect 7389 26741 7423 26775
rect 7423 26741 7432 26775
rect 7380 26732 7432 26741
rect 8852 26732 8904 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 10140 26528 10192 26580
rect 10600 26528 10652 26580
rect 11520 26571 11572 26580
rect 11520 26537 11529 26571
rect 11529 26537 11563 26571
rect 11563 26537 11572 26571
rect 11520 26528 11572 26537
rect 5540 26503 5592 26512
rect 5540 26469 5549 26503
rect 5549 26469 5583 26503
rect 5583 26469 5592 26503
rect 5540 26460 5592 26469
rect 10692 26503 10744 26512
rect 10692 26469 10701 26503
rect 10701 26469 10735 26503
rect 10735 26469 10744 26503
rect 10692 26460 10744 26469
rect 11244 26503 11296 26512
rect 11244 26469 11253 26503
rect 11253 26469 11287 26503
rect 11287 26469 11296 26503
rect 11244 26460 11296 26469
rect 4896 26435 4948 26444
rect 4896 26401 4905 26435
rect 4905 26401 4939 26435
rect 4939 26401 4948 26435
rect 4896 26392 4948 26401
rect 6460 26392 6512 26444
rect 7196 26392 7248 26444
rect 7748 26392 7800 26444
rect 8116 26435 8168 26444
rect 8116 26401 8125 26435
rect 8125 26401 8159 26435
rect 8159 26401 8168 26435
rect 8116 26392 8168 26401
rect 8852 26392 8904 26444
rect 12072 26435 12124 26444
rect 12072 26401 12116 26435
rect 12116 26401 12124 26435
rect 12072 26392 12124 26401
rect 8760 26367 8812 26376
rect 8760 26333 8769 26367
rect 8769 26333 8803 26367
rect 8803 26333 8812 26367
rect 8760 26324 8812 26333
rect 10784 26324 10836 26376
rect 4988 26256 5040 26308
rect 6828 26299 6880 26308
rect 6828 26265 6837 26299
rect 6837 26265 6871 26299
rect 6871 26265 6880 26299
rect 6828 26256 6880 26265
rect 5540 26188 5592 26240
rect 5816 26231 5868 26240
rect 5816 26197 5825 26231
rect 5825 26197 5859 26231
rect 5859 26197 5868 26231
rect 5816 26188 5868 26197
rect 9588 26188 9640 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4896 26027 4948 26036
rect 4896 25993 4905 26027
rect 4905 25993 4939 26027
rect 4939 25993 4948 26027
rect 4896 25984 4948 25993
rect 6460 26027 6512 26036
rect 6460 25993 6469 26027
rect 6469 25993 6503 26027
rect 6503 25993 6512 26027
rect 6460 25984 6512 25993
rect 10600 25984 10652 26036
rect 10692 25984 10744 26036
rect 11980 25984 12032 26036
rect 12072 26027 12124 26036
rect 12072 25993 12081 26027
rect 12081 25993 12115 26027
rect 12115 25993 12124 26027
rect 12072 25984 12124 25993
rect 6092 25848 6144 25900
rect 9588 25848 9640 25900
rect 11520 25848 11572 25900
rect 5172 25780 5224 25832
rect 5816 25780 5868 25832
rect 6920 25780 6972 25832
rect 8024 25823 8076 25832
rect 8024 25789 8033 25823
rect 8033 25789 8067 25823
rect 8067 25789 8076 25823
rect 8024 25780 8076 25789
rect 5264 25687 5316 25696
rect 5264 25653 5273 25687
rect 5273 25653 5307 25687
rect 5307 25653 5316 25687
rect 11244 25780 11296 25832
rect 9404 25712 9456 25764
rect 8852 25687 8904 25696
rect 5264 25644 5316 25653
rect 8852 25653 8861 25687
rect 8861 25653 8895 25687
rect 8895 25653 8904 25687
rect 8852 25644 8904 25653
rect 9772 25644 9824 25696
rect 10048 25644 10100 25696
rect 10784 25644 10836 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 5540 25483 5592 25492
rect 5540 25449 5549 25483
rect 5549 25449 5583 25483
rect 5583 25449 5592 25483
rect 5540 25440 5592 25449
rect 5816 25440 5868 25492
rect 6920 25440 6972 25492
rect 8760 25440 8812 25492
rect 9404 25483 9456 25492
rect 9404 25449 9413 25483
rect 9413 25449 9447 25483
rect 9447 25449 9456 25483
rect 9404 25440 9456 25449
rect 10692 25440 10744 25492
rect 10784 25440 10836 25492
rect 7104 25372 7156 25424
rect 5816 25304 5868 25356
rect 6092 25347 6144 25356
rect 6092 25313 6101 25347
rect 6101 25313 6135 25347
rect 6135 25313 6144 25347
rect 6092 25304 6144 25313
rect 7288 25347 7340 25356
rect 7288 25313 7297 25347
rect 7297 25313 7331 25347
rect 7331 25313 7340 25347
rect 10048 25415 10100 25424
rect 10048 25381 10051 25415
rect 10051 25381 10085 25415
rect 10085 25381 10100 25415
rect 10048 25372 10100 25381
rect 10876 25415 10928 25424
rect 10876 25381 10885 25415
rect 10885 25381 10919 25415
rect 10919 25381 10928 25415
rect 10876 25372 10928 25381
rect 11244 25372 11296 25424
rect 7288 25304 7340 25313
rect 6184 25279 6236 25288
rect 6184 25245 6193 25279
rect 6193 25245 6227 25279
rect 6227 25245 6236 25279
rect 6184 25236 6236 25245
rect 4436 25211 4488 25220
rect 4436 25177 4445 25211
rect 4445 25177 4479 25211
rect 4479 25177 4488 25211
rect 4436 25168 4488 25177
rect 5448 25168 5500 25220
rect 5172 25100 5224 25152
rect 7840 25100 7892 25152
rect 8116 25100 8168 25152
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 6920 24896 6972 24948
rect 7288 24896 7340 24948
rect 5448 24871 5500 24880
rect 5448 24837 5457 24871
rect 5457 24837 5491 24871
rect 5491 24837 5500 24871
rect 5448 24828 5500 24837
rect 7564 24760 7616 24812
rect 7748 24803 7800 24812
rect 7748 24769 7757 24803
rect 7757 24769 7791 24803
rect 7791 24769 7800 24803
rect 7748 24760 7800 24769
rect 8208 24760 8260 24812
rect 8576 24760 8628 24812
rect 8760 24760 8812 24812
rect 10876 24803 10928 24812
rect 10876 24769 10885 24803
rect 10885 24769 10919 24803
rect 10919 24769 10928 24803
rect 10876 24760 10928 24769
rect 11244 24803 11296 24812
rect 11244 24769 11253 24803
rect 11253 24769 11287 24803
rect 11287 24769 11296 24803
rect 11244 24760 11296 24769
rect 3976 24735 4028 24744
rect 3976 24701 3985 24735
rect 3985 24701 4019 24735
rect 4019 24701 4028 24735
rect 3976 24692 4028 24701
rect 4344 24735 4396 24744
rect 4344 24701 4353 24735
rect 4353 24701 4387 24735
rect 4387 24701 4396 24735
rect 4344 24692 4396 24701
rect 5356 24735 5408 24744
rect 5356 24701 5362 24735
rect 5362 24701 5408 24735
rect 5356 24692 5408 24701
rect 6920 24692 6972 24744
rect 3148 24624 3200 24676
rect 4896 24624 4948 24676
rect 5172 24667 5224 24676
rect 5172 24633 5181 24667
rect 5181 24633 5215 24667
rect 5215 24633 5224 24667
rect 5172 24624 5224 24633
rect 6000 24624 6052 24676
rect 3976 24556 4028 24608
rect 5264 24556 5316 24608
rect 7104 24624 7156 24676
rect 10048 24624 10100 24676
rect 8576 24556 8628 24608
rect 9496 24556 9548 24608
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 2780 24352 2832 24404
rect 3148 24395 3200 24404
rect 3148 24361 3157 24395
rect 3157 24361 3191 24395
rect 3191 24361 3200 24395
rect 3148 24352 3200 24361
rect 3332 24352 3384 24404
rect 4436 24352 4488 24404
rect 5356 24352 5408 24404
rect 4160 24284 4212 24336
rect 2964 24259 3016 24268
rect 2964 24225 2973 24259
rect 2973 24225 3007 24259
rect 3007 24225 3016 24259
rect 2964 24216 3016 24225
rect 5724 24259 5776 24268
rect 5724 24225 5733 24259
rect 5733 24225 5767 24259
rect 5767 24225 5776 24259
rect 6828 24352 6880 24404
rect 7196 24395 7248 24404
rect 7196 24361 7205 24395
rect 7205 24361 7239 24395
rect 7239 24361 7248 24395
rect 7196 24352 7248 24361
rect 9680 24352 9732 24404
rect 11244 24327 11296 24336
rect 11244 24293 11253 24327
rect 11253 24293 11287 24327
rect 11287 24293 11296 24327
rect 11244 24284 11296 24293
rect 5724 24216 5776 24225
rect 7564 24216 7616 24268
rect 7840 24259 7892 24268
rect 7840 24225 7849 24259
rect 7849 24225 7883 24259
rect 7883 24225 7892 24259
rect 7840 24216 7892 24225
rect 8300 24259 8352 24268
rect 8300 24225 8309 24259
rect 8309 24225 8343 24259
rect 8343 24225 8352 24259
rect 8300 24216 8352 24225
rect 9680 24259 9732 24268
rect 9680 24225 9689 24259
rect 9689 24225 9723 24259
rect 9723 24225 9732 24259
rect 9680 24216 9732 24225
rect 10140 24259 10192 24268
rect 10140 24225 10149 24259
rect 10149 24225 10183 24259
rect 10183 24225 10192 24259
rect 10140 24216 10192 24225
rect 11060 24216 11112 24268
rect 4068 24148 4120 24200
rect 8576 24148 8628 24200
rect 4344 24080 4396 24132
rect 5540 24080 5592 24132
rect 6184 24080 6236 24132
rect 6828 24123 6880 24132
rect 6828 24089 6837 24123
rect 6837 24089 6871 24123
rect 6871 24089 6880 24123
rect 6828 24080 6880 24089
rect 8852 24080 8904 24132
rect 10140 24080 10192 24132
rect 10508 24080 10560 24132
rect 12348 24080 12400 24132
rect 5816 24012 5868 24064
rect 9312 24012 9364 24064
rect 10600 24012 10652 24064
rect 12716 24012 12768 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 2964 23808 3016 23860
rect 4344 23851 4396 23860
rect 4344 23817 4353 23851
rect 4353 23817 4387 23851
rect 4387 23817 4396 23851
rect 4344 23808 4396 23817
rect 6828 23808 6880 23860
rect 8208 23851 8260 23860
rect 8208 23817 8217 23851
rect 8217 23817 8251 23851
rect 8251 23817 8260 23851
rect 8208 23808 8260 23817
rect 9588 23808 9640 23860
rect 10140 23851 10192 23860
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 11060 23808 11112 23860
rect 12716 23851 12768 23860
rect 12716 23817 12725 23851
rect 12725 23817 12759 23851
rect 12759 23817 12768 23851
rect 12716 23808 12768 23817
rect 3332 23783 3384 23792
rect 3332 23749 3341 23783
rect 3341 23749 3375 23783
rect 3375 23749 3384 23783
rect 3332 23740 3384 23749
rect 7288 23783 7340 23792
rect 7288 23749 7312 23783
rect 7312 23749 7340 23783
rect 7288 23740 7340 23749
rect 8760 23740 8812 23792
rect 3976 23715 4028 23724
rect 3976 23681 3985 23715
rect 3985 23681 4019 23715
rect 4019 23681 4028 23715
rect 3976 23672 4028 23681
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 5540 23715 5592 23724
rect 4712 23672 4764 23681
rect 3240 23647 3292 23656
rect 3240 23613 3249 23647
rect 3249 23613 3283 23647
rect 3283 23613 3292 23647
rect 3240 23604 3292 23613
rect 3516 23647 3568 23656
rect 3516 23613 3525 23647
rect 3525 23613 3559 23647
rect 3559 23613 3568 23647
rect 3516 23604 3568 23613
rect 4988 23647 5040 23656
rect 4988 23613 4997 23647
rect 4997 23613 5031 23647
rect 5031 23613 5040 23647
rect 4988 23604 5040 23613
rect 5540 23681 5549 23715
rect 5549 23681 5583 23715
rect 5583 23681 5592 23715
rect 5540 23672 5592 23681
rect 7564 23672 7616 23724
rect 9312 23740 9364 23792
rect 12624 23783 12676 23792
rect 10508 23715 10560 23724
rect 10508 23681 10517 23715
rect 10517 23681 10551 23715
rect 10551 23681 10560 23715
rect 10508 23672 10560 23681
rect 12624 23749 12648 23783
rect 12648 23749 12676 23783
rect 12624 23740 12676 23749
rect 5724 23604 5776 23656
rect 3976 23536 4028 23588
rect 5172 23536 5224 23588
rect 7840 23604 7892 23656
rect 8576 23604 8628 23656
rect 11980 23604 12032 23656
rect 12532 23604 12584 23656
rect 9404 23579 9456 23588
rect 9404 23545 9413 23579
rect 9413 23545 9447 23579
rect 9447 23545 9456 23579
rect 9404 23536 9456 23545
rect 10508 23536 10560 23588
rect 12348 23536 12400 23588
rect 4896 23511 4948 23520
rect 4896 23477 4905 23511
rect 4905 23477 4939 23511
rect 4939 23477 4948 23511
rect 4896 23468 4948 23477
rect 7840 23468 7892 23520
rect 9680 23511 9732 23520
rect 9680 23477 9689 23511
rect 9689 23477 9723 23511
rect 9723 23477 9732 23511
rect 9680 23468 9732 23477
rect 13084 23511 13136 23520
rect 13084 23477 13093 23511
rect 13093 23477 13127 23511
rect 13127 23477 13136 23511
rect 13084 23468 13136 23477
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 4160 23264 4212 23316
rect 5540 23307 5592 23316
rect 5540 23273 5549 23307
rect 5549 23273 5583 23307
rect 5583 23273 5592 23307
rect 5540 23264 5592 23273
rect 5908 23264 5960 23316
rect 6828 23307 6880 23316
rect 2596 23171 2648 23180
rect 2596 23137 2605 23171
rect 2605 23137 2639 23171
rect 2639 23137 2648 23171
rect 2596 23128 2648 23137
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 2780 23128 2832 23137
rect 3976 23128 4028 23180
rect 4528 23128 4580 23180
rect 4988 23128 5040 23180
rect 5908 23128 5960 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 6276 23171 6328 23180
rect 6276 23137 6285 23171
rect 6285 23137 6319 23171
rect 6319 23137 6328 23171
rect 6276 23128 6328 23137
rect 6828 23273 6837 23307
rect 6837 23273 6871 23307
rect 6871 23273 6880 23307
rect 6828 23264 6880 23273
rect 7288 23264 7340 23316
rect 7564 23307 7616 23316
rect 7564 23273 7573 23307
rect 7573 23273 7607 23307
rect 7607 23273 7616 23307
rect 7564 23264 7616 23273
rect 8300 23264 8352 23316
rect 12532 23264 12584 23316
rect 10508 23239 10560 23248
rect 10508 23205 10517 23239
rect 10517 23205 10551 23239
rect 10551 23205 10560 23239
rect 10508 23196 10560 23205
rect 11980 23196 12032 23248
rect 6828 23128 6880 23180
rect 7932 23128 7984 23180
rect 8484 23171 8536 23180
rect 8484 23137 8493 23171
rect 8493 23137 8527 23171
rect 8527 23137 8536 23171
rect 8484 23128 8536 23137
rect 12072 23171 12124 23180
rect 12072 23137 12081 23171
rect 12081 23137 12115 23171
rect 12115 23137 12124 23171
rect 12072 23128 12124 23137
rect 8760 23103 8812 23112
rect 8760 23069 8769 23103
rect 8769 23069 8803 23103
rect 8803 23069 8812 23103
rect 8760 23060 8812 23069
rect 10416 23103 10468 23112
rect 10416 23069 10425 23103
rect 10425 23069 10459 23103
rect 10459 23069 10468 23103
rect 10416 23060 10468 23069
rect 11152 23060 11204 23112
rect 5632 22992 5684 23044
rect 2964 22924 3016 22976
rect 3516 22967 3568 22976
rect 3516 22933 3525 22967
rect 3525 22933 3559 22967
rect 3559 22933 3568 22967
rect 3516 22924 3568 22933
rect 11060 22924 11112 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2596 22720 2648 22772
rect 5816 22763 5868 22772
rect 5816 22729 5825 22763
rect 5825 22729 5859 22763
rect 5859 22729 5868 22763
rect 5816 22720 5868 22729
rect 5908 22720 5960 22772
rect 6276 22720 6328 22772
rect 7104 22720 7156 22772
rect 7932 22720 7984 22772
rect 12072 22720 12124 22772
rect 12440 22720 12492 22772
rect 12900 22720 12952 22772
rect 3976 22695 4028 22704
rect 3976 22661 3985 22695
rect 3985 22661 4019 22695
rect 4019 22661 4028 22695
rect 3976 22652 4028 22661
rect 7288 22652 7340 22704
rect 8484 22652 8536 22704
rect 4896 22627 4948 22636
rect 4896 22593 4905 22627
rect 4905 22593 4939 22627
rect 4939 22593 4948 22627
rect 4896 22584 4948 22593
rect 6092 22584 6144 22636
rect 6736 22584 6788 22636
rect 7196 22627 7248 22636
rect 7196 22593 7205 22627
rect 7205 22593 7239 22627
rect 7239 22593 7248 22627
rect 7196 22584 7248 22593
rect 8760 22584 8812 22636
rect 10968 22584 11020 22636
rect 11152 22627 11204 22636
rect 11152 22593 11161 22627
rect 11161 22593 11195 22627
rect 11195 22593 11204 22627
rect 11152 22584 11204 22593
rect 9680 22516 9732 22568
rect 10508 22516 10560 22568
rect 12164 22516 12216 22568
rect 13176 22516 13228 22568
rect 3148 22448 3200 22500
rect 3424 22491 3476 22500
rect 3424 22457 3433 22491
rect 3433 22457 3467 22491
rect 3467 22457 3476 22491
rect 3424 22448 3476 22457
rect 3884 22448 3936 22500
rect 5264 22448 5316 22500
rect 6920 22491 6972 22500
rect 6920 22457 6929 22491
rect 6929 22457 6963 22491
rect 6963 22457 6972 22491
rect 6920 22448 6972 22457
rect 4528 22380 4580 22432
rect 6828 22380 6880 22432
rect 7932 22380 7984 22432
rect 9496 22380 9548 22432
rect 10876 22448 10928 22500
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 2780 22176 2832 22228
rect 3424 22219 3476 22228
rect 3424 22185 3433 22219
rect 3433 22185 3467 22219
rect 3467 22185 3476 22219
rect 3424 22176 3476 22185
rect 4896 22176 4948 22228
rect 5816 22176 5868 22228
rect 6828 22176 6880 22228
rect 7288 22176 7340 22228
rect 8760 22176 8812 22228
rect 9496 22176 9548 22228
rect 5264 22108 5316 22160
rect 5540 22108 5592 22160
rect 3056 22083 3108 22092
rect 3056 22049 3074 22083
rect 3074 22049 3108 22083
rect 3056 22040 3108 22049
rect 2228 21972 2280 22024
rect 3424 21972 3476 22024
rect 4988 22015 5040 22024
rect 4988 21981 4997 22015
rect 4997 21981 5031 22015
rect 5031 21981 5040 22015
rect 4988 21972 5040 21981
rect 6184 22108 6236 22160
rect 6920 22108 6972 22160
rect 7932 22108 7984 22160
rect 9680 22108 9732 22160
rect 10876 22176 10928 22228
rect 11612 22151 11664 22160
rect 11612 22117 11621 22151
rect 11621 22117 11655 22151
rect 11655 22117 11664 22151
rect 11612 22108 11664 22117
rect 11980 22108 12032 22160
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 8300 22040 8352 22092
rect 8576 22040 8628 22092
rect 13452 22108 13504 22160
rect 5632 21904 5684 21956
rect 8116 21972 8168 22024
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 11980 21972 12032 22024
rect 12164 22015 12216 22024
rect 12164 21981 12173 22015
rect 12173 21981 12207 22015
rect 12207 21981 12216 22015
rect 12164 21972 12216 21981
rect 13820 21972 13872 22024
rect 7564 21904 7616 21956
rect 10968 21904 11020 21956
rect 12532 21904 12584 21956
rect 4804 21836 4856 21888
rect 11520 21836 11572 21888
rect 12348 21836 12400 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 4988 21632 5040 21684
rect 5264 21632 5316 21684
rect 7932 21632 7984 21684
rect 8760 21632 8812 21684
rect 3424 21564 3476 21616
rect 4712 21539 4764 21548
rect 4712 21505 4721 21539
rect 4721 21505 4755 21539
rect 4755 21505 4764 21539
rect 4712 21496 4764 21505
rect 4988 21539 5040 21548
rect 4988 21505 4997 21539
rect 4997 21505 5031 21539
rect 5031 21505 5040 21539
rect 4988 21496 5040 21505
rect 7656 21428 7708 21480
rect 8392 21471 8444 21480
rect 8392 21437 8401 21471
rect 8401 21437 8435 21471
rect 8435 21437 8444 21471
rect 8392 21428 8444 21437
rect 4804 21403 4856 21412
rect 4804 21369 4813 21403
rect 4813 21369 4847 21403
rect 4847 21369 4856 21403
rect 4804 21360 4856 21369
rect 8668 21403 8720 21412
rect 8668 21369 8677 21403
rect 8677 21369 8711 21403
rect 8711 21369 8720 21403
rect 8668 21360 8720 21369
rect 11612 21632 11664 21684
rect 11980 21632 12032 21684
rect 13452 21675 13504 21684
rect 13452 21641 13461 21675
rect 13461 21641 13495 21675
rect 13495 21641 13504 21675
rect 13452 21632 13504 21641
rect 13820 21675 13872 21684
rect 13820 21641 13829 21675
rect 13829 21641 13863 21675
rect 13863 21641 13872 21675
rect 13820 21632 13872 21641
rect 9680 21564 9732 21616
rect 12164 21496 12216 21548
rect 9588 21471 9640 21480
rect 9588 21437 9597 21471
rect 9597 21437 9631 21471
rect 9631 21437 9640 21471
rect 9588 21428 9640 21437
rect 10784 21428 10836 21480
rect 11336 21428 11388 21480
rect 9956 21360 10008 21412
rect 12532 21403 12584 21412
rect 12532 21369 12541 21403
rect 12541 21369 12575 21403
rect 12575 21369 12584 21403
rect 12532 21360 12584 21369
rect 12624 21403 12676 21412
rect 12624 21369 12633 21403
rect 12633 21369 12667 21403
rect 12667 21369 12676 21403
rect 12624 21360 12676 21369
rect 3056 21335 3108 21344
rect 3056 21301 3065 21335
rect 3065 21301 3099 21335
rect 3099 21301 3108 21335
rect 3056 21292 3108 21301
rect 3516 21292 3568 21344
rect 5908 21292 5960 21344
rect 6828 21292 6880 21344
rect 7288 21292 7340 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 7656 21088 7708 21140
rect 8116 21131 8168 21140
rect 8116 21097 8125 21131
rect 8125 21097 8159 21131
rect 8159 21097 8168 21131
rect 8116 21088 8168 21097
rect 8668 21088 8720 21140
rect 12624 21088 12676 21140
rect 13176 21088 13228 21140
rect 7196 21063 7248 21072
rect 7196 21029 7205 21063
rect 7205 21029 7239 21063
rect 7239 21029 7248 21063
rect 7196 21020 7248 21029
rect 7380 21020 7432 21072
rect 4804 20995 4856 21004
rect 4804 20961 4813 20995
rect 4813 20961 4847 20995
rect 4847 20961 4856 20995
rect 4804 20952 4856 20961
rect 6092 20952 6144 21004
rect 6368 20952 6420 21004
rect 9956 21020 10008 21072
rect 11520 21020 11572 21072
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 6552 20884 6604 20936
rect 8208 20952 8260 21004
rect 13084 20995 13136 21004
rect 13084 20961 13102 20995
rect 13102 20961 13136 20995
rect 8392 20884 8444 20936
rect 13084 20952 13136 20961
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 11152 20884 11204 20936
rect 12164 20927 12216 20936
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 12532 20884 12584 20936
rect 13084 20816 13136 20868
rect 9588 20748 9640 20800
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 4436 20544 4488 20596
rect 4804 20544 4856 20596
rect 6552 20587 6604 20596
rect 6552 20553 6561 20587
rect 6561 20553 6595 20587
rect 6595 20553 6604 20587
rect 6552 20544 6604 20553
rect 4988 20519 5040 20528
rect 4988 20485 4997 20519
rect 4997 20485 5031 20519
rect 5031 20485 5040 20519
rect 4988 20476 5040 20485
rect 8300 20544 8352 20596
rect 8760 20587 8812 20596
rect 8760 20553 8769 20587
rect 8769 20553 8803 20587
rect 8803 20553 8812 20587
rect 8760 20544 8812 20553
rect 9312 20544 9364 20596
rect 11520 20544 11572 20596
rect 12440 20544 12492 20596
rect 13084 20544 13136 20596
rect 8668 20408 8720 20460
rect 10968 20476 11020 20528
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 4528 20315 4580 20324
rect 4528 20281 4537 20315
rect 4537 20281 4571 20315
rect 4571 20281 4580 20315
rect 4528 20272 4580 20281
rect 5540 20272 5592 20324
rect 6368 20272 6420 20324
rect 9680 20340 9732 20392
rect 12532 20383 12584 20392
rect 12532 20349 12534 20383
rect 12534 20349 12584 20383
rect 12532 20340 12584 20349
rect 13452 20383 13504 20392
rect 13452 20349 13496 20383
rect 13496 20349 13504 20383
rect 13912 20383 13964 20392
rect 13452 20340 13504 20349
rect 13912 20349 13921 20383
rect 13921 20349 13955 20383
rect 13955 20349 13964 20383
rect 13912 20340 13964 20349
rect 7748 20272 7800 20324
rect 8208 20272 8260 20324
rect 9312 20315 9364 20324
rect 9312 20281 9315 20315
rect 9315 20281 9349 20315
rect 9349 20281 9364 20315
rect 9312 20272 9364 20281
rect 10968 20272 11020 20324
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 2872 20000 2924 20052
rect 6184 20000 6236 20052
rect 6828 20000 6880 20052
rect 3148 19864 3200 19916
rect 4988 19932 5040 19984
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 9680 20000 9732 20052
rect 10968 20000 11020 20052
rect 11980 20000 12032 20052
rect 10232 19932 10284 19984
rect 11428 19932 11480 19984
rect 12072 19932 12124 19984
rect 7656 19907 7708 19916
rect 4988 19839 5040 19848
rect 4988 19805 4997 19839
rect 4997 19805 5031 19839
rect 5031 19805 5040 19839
rect 4988 19796 5040 19805
rect 6276 19796 6328 19848
rect 7656 19873 7665 19907
rect 7665 19873 7699 19907
rect 7699 19873 7708 19907
rect 7656 19864 7708 19873
rect 8392 19864 8444 19916
rect 10048 19864 10100 19916
rect 7012 19796 7064 19848
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 10876 19839 10928 19848
rect 10876 19805 10885 19839
rect 10885 19805 10919 19839
rect 10919 19805 10928 19839
rect 10876 19796 10928 19805
rect 8484 19728 8536 19780
rect 5264 19703 5316 19712
rect 5264 19669 5273 19703
rect 5273 19669 5307 19703
rect 5307 19669 5316 19703
rect 6092 19703 6144 19712
rect 5264 19660 5316 19669
rect 6092 19669 6101 19703
rect 6101 19669 6135 19703
rect 6135 19669 6144 19703
rect 6092 19660 6144 19669
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 3148 19456 3200 19508
rect 6276 19499 6328 19508
rect 6276 19465 6285 19499
rect 6285 19465 6319 19499
rect 6319 19465 6328 19499
rect 6276 19456 6328 19465
rect 10968 19499 11020 19508
rect 10968 19465 10977 19499
rect 10977 19465 11011 19499
rect 11011 19465 11020 19499
rect 10968 19456 11020 19465
rect 5264 19431 5316 19440
rect 5264 19397 5273 19431
rect 5273 19397 5307 19431
rect 5307 19397 5316 19431
rect 5264 19388 5316 19397
rect 8484 19431 8536 19440
rect 8484 19397 8493 19431
rect 8493 19397 8527 19431
rect 8527 19397 8536 19431
rect 8484 19388 8536 19397
rect 4896 19320 4948 19372
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 5264 19252 5316 19304
rect 6092 19320 6144 19372
rect 7472 19320 7524 19372
rect 7932 19320 7984 19372
rect 7656 19252 7708 19304
rect 6920 19184 6972 19236
rect 7564 19227 7616 19236
rect 7564 19193 7573 19227
rect 7573 19193 7607 19227
rect 7607 19193 7616 19227
rect 7564 19184 7616 19193
rect 7932 19184 7984 19236
rect 8760 19252 8812 19304
rect 9772 19252 9824 19304
rect 10048 19252 10100 19304
rect 9588 19184 9640 19236
rect 4344 19159 4396 19168
rect 4344 19125 4353 19159
rect 4353 19125 4387 19159
rect 4387 19125 4396 19159
rect 4344 19116 4396 19125
rect 5448 19116 5500 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 6184 19116 6236 19168
rect 6644 19116 6696 19168
rect 6828 19116 6880 19168
rect 8300 19116 8352 19168
rect 9772 19159 9824 19168
rect 9772 19125 9781 19159
rect 9781 19125 9815 19159
rect 9815 19125 9824 19159
rect 9772 19116 9824 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 4160 18912 4212 18964
rect 6092 18955 6144 18964
rect 6092 18921 6101 18955
rect 6101 18921 6135 18955
rect 6135 18921 6144 18955
rect 6092 18912 6144 18921
rect 7012 18912 7064 18964
rect 10232 18912 10284 18964
rect 6828 18844 6880 18896
rect 8760 18844 8812 18896
rect 4988 18819 5040 18828
rect 4988 18785 4997 18819
rect 4997 18785 5031 18819
rect 5031 18785 5040 18819
rect 4988 18776 5040 18785
rect 5264 18776 5316 18828
rect 5816 18776 5868 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 5448 18708 5500 18760
rect 6184 18708 6236 18760
rect 6920 18776 6972 18828
rect 8208 18819 8260 18828
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 6644 18708 6696 18760
rect 4804 18683 4856 18692
rect 4804 18649 4813 18683
rect 4813 18649 4847 18683
rect 4847 18649 4856 18683
rect 4804 18640 4856 18649
rect 6828 18640 6880 18692
rect 7012 18640 7064 18692
rect 8392 18640 8444 18692
rect 10692 18819 10744 18828
rect 10692 18785 10701 18819
rect 10701 18785 10735 18819
rect 10735 18785 10744 18819
rect 10692 18776 10744 18785
rect 9588 18708 9640 18760
rect 11520 18708 11572 18760
rect 5816 18615 5868 18624
rect 5816 18581 5825 18615
rect 5825 18581 5859 18615
rect 5859 18581 5868 18615
rect 5816 18572 5868 18581
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 2872 18411 2924 18420
rect 2872 18377 2881 18411
rect 2881 18377 2915 18411
rect 2915 18377 2924 18411
rect 2872 18368 2924 18377
rect 4988 18368 5040 18420
rect 6276 18368 6328 18420
rect 7932 18368 7984 18420
rect 8760 18368 8812 18420
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 4068 18300 4120 18352
rect 4804 18343 4856 18352
rect 4804 18309 4813 18343
rect 4813 18309 4847 18343
rect 4847 18309 4856 18343
rect 4804 18300 4856 18309
rect 5816 18300 5868 18352
rect 2872 18164 2924 18216
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 5448 18207 5500 18216
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 7196 18164 7248 18216
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 5356 18096 5408 18148
rect 7380 18139 7432 18148
rect 7380 18105 7389 18139
rect 7389 18105 7423 18139
rect 7423 18105 7432 18139
rect 11060 18164 11112 18216
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 7380 18096 7432 18105
rect 10048 18096 10100 18148
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5080 18028 5132 18037
rect 11152 18028 11204 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 6184 17824 6236 17876
rect 6828 17824 6880 17876
rect 5264 17799 5316 17808
rect 5264 17765 5267 17799
rect 5267 17765 5301 17799
rect 5301 17765 5316 17799
rect 5264 17756 5316 17765
rect 3148 17688 3200 17740
rect 5080 17688 5132 17740
rect 7288 17688 7340 17740
rect 8208 17824 8260 17876
rect 8576 17867 8628 17876
rect 8576 17833 8585 17867
rect 8585 17833 8619 17867
rect 8619 17833 8628 17867
rect 8576 17824 8628 17833
rect 9404 17867 9456 17876
rect 9404 17833 9413 17867
rect 9413 17833 9447 17867
rect 9447 17833 9456 17867
rect 9404 17824 9456 17833
rect 11060 17824 11112 17876
rect 11428 17824 11480 17876
rect 10048 17799 10100 17808
rect 10048 17765 10051 17799
rect 10051 17765 10085 17799
rect 10085 17765 10100 17799
rect 10048 17756 10100 17765
rect 11520 17799 11572 17808
rect 11520 17765 11529 17799
rect 11529 17765 11563 17799
rect 11563 17765 11572 17799
rect 11520 17756 11572 17765
rect 7012 17620 7064 17672
rect 8116 17688 8168 17740
rect 9680 17731 9732 17740
rect 9680 17697 9689 17731
rect 9689 17697 9723 17731
rect 9723 17697 9732 17731
rect 9680 17688 9732 17697
rect 8024 17663 8076 17672
rect 8024 17629 8033 17663
rect 8033 17629 8067 17663
rect 8067 17629 8076 17663
rect 8024 17620 8076 17629
rect 12808 17620 12860 17672
rect 4896 17484 4948 17536
rect 5448 17484 5500 17536
rect 5724 17484 5776 17536
rect 7196 17484 7248 17536
rect 12164 17484 12216 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 3148 17280 3200 17332
rect 4252 17323 4304 17332
rect 4252 17289 4261 17323
rect 4261 17289 4295 17323
rect 4295 17289 4304 17323
rect 4252 17280 4304 17289
rect 5080 17280 5132 17332
rect 5356 17280 5408 17332
rect 7012 17280 7064 17332
rect 7380 17323 7432 17332
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 5816 17212 5868 17264
rect 7288 17212 7340 17264
rect 4068 17144 4120 17196
rect 5264 17187 5316 17196
rect 4252 17076 4304 17128
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 8208 17144 8260 17196
rect 5632 17076 5684 17128
rect 7380 17076 7432 17128
rect 7932 17076 7984 17128
rect 9128 17119 9180 17128
rect 9128 17085 9137 17119
rect 9137 17085 9171 17119
rect 9171 17085 9180 17119
rect 9128 17076 9180 17085
rect 6000 17008 6052 17060
rect 10048 17280 10100 17332
rect 11336 17323 11388 17332
rect 11336 17289 11345 17323
rect 11345 17289 11379 17323
rect 11379 17289 11388 17323
rect 11336 17280 11388 17289
rect 11520 17280 11572 17332
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 9864 17076 9916 17128
rect 11336 17076 11388 17128
rect 12164 17008 12216 17060
rect 3976 16940 4028 16992
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 11060 16940 11112 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 4068 16736 4120 16788
rect 5816 16779 5868 16788
rect 5816 16745 5825 16779
rect 5825 16745 5859 16779
rect 5859 16745 5868 16779
rect 5816 16736 5868 16745
rect 6828 16736 6880 16788
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 9680 16736 9732 16788
rect 10048 16736 10100 16788
rect 2872 16600 2924 16652
rect 5356 16668 5408 16720
rect 5908 16668 5960 16720
rect 7932 16668 7984 16720
rect 8208 16711 8260 16720
rect 8208 16677 8211 16711
rect 8211 16677 8245 16711
rect 8245 16677 8260 16711
rect 8208 16668 8260 16677
rect 8576 16668 8628 16720
rect 10692 16711 10744 16720
rect 10692 16677 10701 16711
rect 10701 16677 10735 16711
rect 10735 16677 10744 16711
rect 10692 16668 10744 16677
rect 11428 16736 11480 16788
rect 12164 16668 12216 16720
rect 12808 16711 12860 16720
rect 12808 16677 12817 16711
rect 12817 16677 12851 16711
rect 12851 16677 12860 16711
rect 12808 16668 12860 16677
rect 5448 16643 5500 16652
rect 4804 16532 4856 16584
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 7380 16600 7432 16652
rect 8024 16600 8076 16652
rect 8300 16600 8352 16652
rect 9588 16600 9640 16652
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 11152 16507 11204 16516
rect 11152 16473 11161 16507
rect 11161 16473 11195 16507
rect 11195 16473 11204 16507
rect 12624 16532 12676 16584
rect 11152 16464 11204 16473
rect 4896 16396 4948 16448
rect 5632 16396 5684 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 2872 16192 2924 16244
rect 3976 16235 4028 16244
rect 3976 16201 3985 16235
rect 3985 16201 4019 16235
rect 4019 16201 4028 16235
rect 3976 16192 4028 16201
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 7380 16235 7432 16244
rect 7380 16201 7389 16235
rect 7389 16201 7423 16235
rect 7423 16201 7432 16235
rect 7380 16192 7432 16201
rect 8576 16235 8628 16244
rect 8576 16201 8585 16235
rect 8585 16201 8619 16235
rect 8619 16201 8628 16235
rect 8576 16192 8628 16201
rect 8760 16192 8812 16244
rect 10600 16192 10652 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 12624 16192 12676 16244
rect 3976 15988 4028 16040
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 8852 16056 8904 16108
rect 5816 15963 5868 15972
rect 5816 15929 5825 15963
rect 5825 15929 5859 15963
rect 5859 15929 5868 15963
rect 5816 15920 5868 15929
rect 6552 15920 6604 15972
rect 7104 15963 7156 15972
rect 7104 15929 7113 15963
rect 7113 15929 7147 15963
rect 7147 15929 7156 15963
rect 7104 15920 7156 15929
rect 7748 15920 7800 15972
rect 8392 15920 8444 15972
rect 12716 16056 12768 16108
rect 9956 15920 10008 15972
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 10876 15852 10928 15904
rect 12808 15988 12860 16040
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 5356 15648 5408 15700
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 7840 15648 7892 15700
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 8668 15691 8720 15700
rect 8668 15657 8677 15691
rect 8677 15657 8711 15691
rect 8711 15657 8720 15691
rect 8668 15648 8720 15657
rect 8852 15648 8904 15700
rect 10600 15648 10652 15700
rect 5264 15580 5316 15632
rect 5448 15580 5500 15632
rect 5632 15580 5684 15632
rect 7104 15555 7156 15564
rect 7104 15521 7113 15555
rect 7113 15521 7147 15555
rect 7147 15521 7156 15555
rect 7104 15512 7156 15521
rect 9956 15580 10008 15632
rect 11060 15580 11112 15632
rect 11520 15623 11572 15632
rect 11520 15589 11529 15623
rect 11529 15589 11563 15623
rect 11563 15589 11572 15623
rect 11520 15580 11572 15589
rect 11704 15580 11756 15632
rect 8024 15512 8076 15564
rect 8484 15555 8536 15564
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 8484 15512 8536 15521
rect 9772 15512 9824 15564
rect 12256 15512 12308 15564
rect 12992 15555 13044 15564
rect 12992 15521 13036 15555
rect 13036 15521 13044 15555
rect 12992 15512 13044 15521
rect 5816 15444 5868 15496
rect 12348 15444 12400 15496
rect 6092 15351 6144 15360
rect 6092 15317 6101 15351
rect 6101 15317 6135 15351
rect 6135 15317 6144 15351
rect 6092 15308 6144 15317
rect 10600 15351 10652 15360
rect 10600 15317 10609 15351
rect 10609 15317 10643 15351
rect 10643 15317 10652 15351
rect 10600 15308 10652 15317
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 12808 15308 12860 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 5448 15104 5500 15156
rect 8024 15147 8076 15156
rect 4160 14900 4212 14952
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5264 14900 5316 14909
rect 5632 14900 5684 14952
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 8760 15147 8812 15156
rect 8760 15113 8769 15147
rect 8769 15113 8803 15147
rect 8803 15113 8812 15147
rect 8760 15104 8812 15113
rect 9956 15104 10008 15156
rect 10600 15147 10652 15156
rect 10600 15113 10609 15147
rect 10609 15113 10643 15147
rect 10643 15113 10652 15147
rect 10600 15104 10652 15113
rect 11704 15147 11756 15156
rect 11704 15113 11713 15147
rect 11713 15113 11747 15147
rect 11747 15113 11756 15147
rect 11704 15104 11756 15113
rect 13544 15104 13596 15156
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 8392 14968 8444 15020
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 10968 14968 11020 15020
rect 12716 14900 12768 14952
rect 13268 14900 13320 14952
rect 8760 14832 8812 14884
rect 10600 14832 10652 14884
rect 11060 14832 11112 14884
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 6644 14764 6696 14816
rect 6828 14764 6880 14816
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 9864 14807 9916 14816
rect 9864 14773 9873 14807
rect 9873 14773 9907 14807
rect 9907 14773 9916 14807
rect 9864 14764 9916 14773
rect 11980 14764 12032 14816
rect 12992 14807 13044 14816
rect 12992 14773 13001 14807
rect 13001 14773 13035 14807
rect 13035 14773 13044 14807
rect 12992 14764 13044 14773
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 5264 14560 5316 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 7104 14560 7156 14612
rect 6644 14492 6696 14544
rect 7748 14492 7800 14544
rect 5080 14467 5132 14476
rect 5080 14433 5098 14467
rect 5098 14433 5132 14467
rect 5080 14424 5132 14433
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 8484 14560 8536 14612
rect 8668 14560 8720 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 9772 14560 9824 14612
rect 11520 14603 11572 14612
rect 11520 14569 11529 14603
rect 11529 14569 11563 14603
rect 11563 14569 11572 14603
rect 11520 14560 11572 14569
rect 9864 14492 9916 14544
rect 11152 14492 11204 14544
rect 12440 14492 12492 14544
rect 11060 14467 11112 14476
rect 11060 14433 11069 14467
rect 11069 14433 11103 14467
rect 11103 14433 11112 14467
rect 11060 14424 11112 14433
rect 6460 14399 6512 14408
rect 6460 14365 6469 14399
rect 6469 14365 6503 14399
rect 6503 14365 6512 14399
rect 6460 14356 6512 14365
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 8300 14356 8352 14408
rect 11612 14356 11664 14408
rect 12808 14356 12860 14408
rect 4252 14220 4304 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 4068 14016 4120 14068
rect 4436 14059 4488 14068
rect 4436 14025 4445 14059
rect 4445 14025 4479 14059
rect 4479 14025 4488 14059
rect 4436 14016 4488 14025
rect 3424 13991 3476 14000
rect 3424 13957 3433 13991
rect 3433 13957 3467 13991
rect 3467 13957 3476 13991
rect 3424 13948 3476 13957
rect 4160 13880 4212 13932
rect 5080 14016 5132 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 7012 14016 7064 14068
rect 8116 14016 8168 14068
rect 10324 14016 10376 14068
rect 10600 14016 10652 14068
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 11612 14059 11664 14068
rect 11612 14025 11621 14059
rect 11621 14025 11655 14059
rect 11655 14025 11664 14059
rect 11612 14016 11664 14025
rect 11980 14016 12032 14068
rect 12808 14016 12860 14068
rect 5264 13880 5316 13932
rect 6920 13880 6972 13932
rect 4068 13812 4120 13864
rect 5540 13812 5592 13864
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 8116 13812 8168 13864
rect 8760 13812 8812 13864
rect 12440 13880 12492 13932
rect 5264 13787 5316 13796
rect 5264 13753 5267 13787
rect 5267 13753 5301 13787
rect 5301 13753 5316 13787
rect 6920 13787 6972 13796
rect 5264 13744 5316 13753
rect 6920 13753 6929 13787
rect 6929 13753 6963 13787
rect 6963 13753 6972 13787
rect 6920 13744 6972 13753
rect 7012 13787 7064 13796
rect 7012 13753 7021 13787
rect 7021 13753 7055 13787
rect 7055 13753 7064 13787
rect 10232 13787 10284 13796
rect 7012 13744 7064 13753
rect 10232 13753 10241 13787
rect 10241 13753 10275 13787
rect 10275 13753 10284 13787
rect 10232 13744 10284 13753
rect 10324 13787 10376 13796
rect 10324 13753 10333 13787
rect 10333 13753 10367 13787
rect 10367 13753 10376 13787
rect 10324 13744 10376 13753
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 4252 13447 4304 13456
rect 4252 13413 4261 13447
rect 4261 13413 4295 13447
rect 4295 13413 4304 13447
rect 4252 13404 4304 13413
rect 4344 13447 4396 13456
rect 4344 13413 4353 13447
rect 4353 13413 4387 13447
rect 4387 13413 4396 13447
rect 4344 13404 4396 13413
rect 5448 13404 5500 13456
rect 4988 13336 5040 13388
rect 6092 13404 6144 13456
rect 6644 13472 6696 13524
rect 6920 13472 6972 13524
rect 8760 13472 8812 13524
rect 10232 13472 10284 13524
rect 7656 13404 7708 13456
rect 9864 13447 9916 13456
rect 9864 13413 9873 13447
rect 9873 13413 9907 13447
rect 9907 13413 9916 13447
rect 9864 13404 9916 13413
rect 11152 13336 11204 13388
rect 5632 13268 5684 13320
rect 5816 13268 5868 13320
rect 7564 13268 7616 13320
rect 8668 13268 8720 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 10508 13268 10560 13320
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 4252 12928 4304 12980
rect 6092 12928 6144 12980
rect 7656 12971 7708 12980
rect 7656 12937 7665 12971
rect 7665 12937 7699 12971
rect 7699 12937 7708 12971
rect 7656 12928 7708 12937
rect 8668 12928 8720 12980
rect 9772 12928 9824 12980
rect 11060 12928 11112 12980
rect 11152 12928 11204 12980
rect 12532 12928 12584 12980
rect 4344 12860 4396 12912
rect 5816 12903 5868 12912
rect 5816 12869 5825 12903
rect 5825 12869 5859 12903
rect 5859 12869 5868 12903
rect 5816 12860 5868 12869
rect 4988 12792 5040 12844
rect 8208 12792 8260 12844
rect 5080 12724 5132 12776
rect 5264 12699 5316 12708
rect 5264 12665 5273 12699
rect 5273 12665 5307 12699
rect 5307 12665 5316 12699
rect 5264 12656 5316 12665
rect 5448 12656 5500 12708
rect 7656 12656 7708 12708
rect 5908 12588 5960 12640
rect 6184 12588 6236 12640
rect 8208 12588 8260 12640
rect 9864 12792 9916 12844
rect 11152 12767 11204 12776
rect 11152 12733 11170 12767
rect 11170 12733 11204 12767
rect 11152 12724 11204 12733
rect 8760 12656 8812 12708
rect 9588 12699 9640 12708
rect 9588 12665 9597 12699
rect 9597 12665 9631 12699
rect 9631 12665 9640 12699
rect 9588 12656 9640 12665
rect 10232 12699 10284 12708
rect 10232 12665 10241 12699
rect 10241 12665 10275 12699
rect 10275 12665 10284 12699
rect 10232 12656 10284 12665
rect 11336 12588 11388 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 4988 12384 5040 12436
rect 5264 12384 5316 12436
rect 5632 12384 5684 12436
rect 6184 12316 6236 12368
rect 7104 12384 7156 12436
rect 7656 12384 7708 12436
rect 7932 12384 7984 12436
rect 9956 12384 10008 12436
rect 10508 12384 10560 12436
rect 7288 12316 7340 12368
rect 8116 12316 8168 12368
rect 8576 12316 8628 12368
rect 9496 12316 9548 12368
rect 11428 12359 11480 12368
rect 11428 12325 11437 12359
rect 11437 12325 11471 12359
rect 11471 12325 11480 12359
rect 11428 12316 11480 12325
rect 4712 12248 4764 12300
rect 12808 12291 12860 12300
rect 12808 12257 12852 12291
rect 12852 12257 12860 12291
rect 12808 12248 12860 12257
rect 5632 12180 5684 12232
rect 7840 12180 7892 12232
rect 9404 12180 9456 12232
rect 11336 12223 11388 12232
rect 7656 12112 7708 12164
rect 8024 12112 8076 12164
rect 10232 12112 10284 12164
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 9588 12044 9640 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 5356 11840 5408 11892
rect 4712 11772 4764 11824
rect 5172 11815 5224 11824
rect 5172 11781 5181 11815
rect 5181 11781 5215 11815
rect 5215 11781 5224 11815
rect 5172 11772 5224 11781
rect 5816 11840 5868 11892
rect 6184 11840 6236 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 8760 11840 8812 11892
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 11336 11840 11388 11892
rect 11428 11840 11480 11892
rect 12808 11840 12860 11892
rect 7932 11772 7984 11824
rect 9128 11704 9180 11756
rect 10508 11704 10560 11756
rect 11060 11704 11112 11756
rect 6092 11636 6144 11688
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 11244 11679 11296 11688
rect 11244 11645 11288 11679
rect 11288 11645 11296 11679
rect 11244 11636 11296 11645
rect 12624 11636 12676 11688
rect 12992 11636 13044 11688
rect 7932 11568 7984 11620
rect 10416 11611 10468 11620
rect 5632 11500 5684 11552
rect 9680 11500 9732 11552
rect 10416 11577 10425 11611
rect 10425 11577 10459 11611
rect 10459 11577 10468 11611
rect 10416 11568 10468 11577
rect 10784 11500 10836 11552
rect 11244 11500 11296 11552
rect 12440 11500 12492 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 6184 11296 6236 11348
rect 4068 11160 4120 11212
rect 4804 11160 4856 11212
rect 5816 11160 5868 11212
rect 6552 11203 6604 11212
rect 6552 11169 6561 11203
rect 6561 11169 6595 11203
rect 6595 11169 6604 11203
rect 6552 11160 6604 11169
rect 7104 11296 7156 11348
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 12072 11296 12124 11348
rect 7748 11228 7800 11280
rect 7932 11228 7984 11280
rect 9496 11228 9548 11280
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 12532 11160 12584 11212
rect 8300 11092 8352 11144
rect 10232 11092 10284 11144
rect 10968 11092 11020 11144
rect 5356 11024 5408 11076
rect 5816 11024 5868 11076
rect 7748 11067 7800 11076
rect 7748 11033 7757 11067
rect 7757 11033 7791 11067
rect 7791 11033 7800 11067
rect 7748 11024 7800 11033
rect 5632 10956 5684 11008
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 11060 10956 11112 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 4068 10795 4120 10804
rect 4068 10761 4077 10795
rect 4077 10761 4111 10795
rect 4111 10761 4120 10795
rect 4068 10752 4120 10761
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 6552 10752 6604 10804
rect 7932 10795 7984 10804
rect 7932 10761 7941 10795
rect 7941 10761 7975 10795
rect 7975 10761 7984 10795
rect 7932 10752 7984 10761
rect 8760 10752 8812 10804
rect 9496 10795 9548 10804
rect 9496 10761 9505 10795
rect 9505 10761 9539 10795
rect 9539 10761 9548 10795
rect 9496 10752 9548 10761
rect 11152 10752 11204 10804
rect 12532 10752 12584 10804
rect 13176 10752 13228 10804
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 7104 10616 7156 10668
rect 9312 10684 9364 10736
rect 8024 10616 8076 10668
rect 8760 10616 8812 10668
rect 9404 10616 9456 10668
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 5264 10523 5316 10532
rect 5264 10489 5273 10523
rect 5273 10489 5307 10523
rect 5307 10489 5316 10523
rect 5264 10480 5316 10489
rect 5448 10480 5500 10532
rect 7012 10523 7064 10532
rect 7012 10489 7021 10523
rect 7021 10489 7055 10523
rect 7055 10489 7064 10523
rect 7012 10480 7064 10489
rect 8668 10523 8720 10532
rect 8668 10489 8677 10523
rect 8677 10489 8711 10523
rect 8711 10489 8720 10523
rect 8668 10480 8720 10489
rect 10140 10523 10192 10532
rect 10140 10489 10149 10523
rect 10149 10489 10183 10523
rect 10183 10489 10192 10523
rect 10140 10480 10192 10489
rect 10600 10412 10652 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 10600 10251 10652 10260
rect 10600 10217 10609 10251
rect 10609 10217 10643 10251
rect 10643 10217 10652 10251
rect 10600 10208 10652 10217
rect 6276 10140 6328 10192
rect 7472 10183 7524 10192
rect 7472 10149 7481 10183
rect 7481 10149 7515 10183
rect 7515 10149 7524 10183
rect 7472 10140 7524 10149
rect 8024 10183 8076 10192
rect 8024 10149 8033 10183
rect 8033 10149 8067 10183
rect 8067 10149 8076 10183
rect 8024 10140 8076 10149
rect 10048 10183 10100 10192
rect 10048 10149 10051 10183
rect 10051 10149 10085 10183
rect 10085 10149 10100 10183
rect 10048 10140 10100 10149
rect 10140 10140 10192 10192
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 7012 10072 7064 10124
rect 10416 10072 10468 10124
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 7564 10004 7616 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 7932 9664 7984 9716
rect 10042 9664 10094 9716
rect 10416 9664 10468 9716
rect 7472 9596 7524 9648
rect 5448 9460 5500 9512
rect 7012 9460 7064 9512
rect 9680 9528 9732 9580
rect 8576 9503 8628 9512
rect 6276 9392 6328 9444
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 9864 9460 9916 9512
rect 10416 9503 10468 9512
rect 6184 9324 6236 9376
rect 9588 9392 9640 9444
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 4712 9120 4764 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 5540 9120 5592 9172
rect 6920 9120 6972 9172
rect 8576 9120 8628 9172
rect 8760 9163 8812 9172
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 9772 9120 9824 9172
rect 5632 9052 5684 9104
rect 7748 9052 7800 9104
rect 7932 9052 7984 9104
rect 10416 9052 10468 9104
rect 4344 9027 4396 9036
rect 4344 8993 4388 9027
rect 4388 8993 4396 9027
rect 4344 8984 4396 8993
rect 5264 8984 5316 9036
rect 5724 8984 5776 9036
rect 4528 8916 4580 8968
rect 6184 8984 6236 9036
rect 7012 8984 7064 9036
rect 9956 8984 10008 9036
rect 10140 8984 10192 9036
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 10232 8891 10284 8900
rect 10232 8857 10241 8891
rect 10241 8857 10275 8891
rect 10275 8857 10284 8891
rect 10232 8848 10284 8857
rect 4068 8780 4120 8832
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4344 8619 4396 8628
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 4436 8576 4488 8628
rect 4804 8576 4856 8628
rect 5816 8576 5868 8628
rect 10692 8576 10744 8628
rect 7748 8551 7800 8560
rect 7748 8517 7757 8551
rect 7757 8517 7791 8551
rect 7791 8517 7800 8551
rect 7748 8508 7800 8517
rect 7104 8440 7156 8492
rect 7932 8440 7984 8492
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 5816 8372 5868 8424
rect 6000 8372 6052 8424
rect 8668 8372 8720 8424
rect 8852 8440 8904 8492
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 8116 8304 8168 8356
rect 8852 8304 8904 8356
rect 9956 8304 10008 8356
rect 12256 8304 12308 8356
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 6184 7964 6236 8016
rect 8116 8007 8168 8016
rect 8116 7973 8125 8007
rect 8125 7973 8159 8007
rect 8159 7973 8168 8007
rect 8116 7964 8168 7973
rect 10048 8007 10100 8016
rect 10048 7973 10051 8007
rect 10051 7973 10085 8007
rect 10085 7973 10100 8007
rect 10048 7964 10100 7973
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 5632 7896 5684 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 6092 7828 6144 7880
rect 5540 7692 5592 7744
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7840 7828 7892 7880
rect 8760 7828 8812 7880
rect 11060 7828 11112 7880
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 5632 7488 5684 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 9680 7488 9732 7540
rect 5080 7420 5132 7472
rect 6092 7352 6144 7404
rect 7012 7352 7064 7404
rect 8852 7352 8904 7404
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 6920 7216 6972 7268
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 7748 7216 7800 7268
rect 10048 7420 10100 7472
rect 11704 7420 11756 7472
rect 11152 7284 11204 7336
rect 7288 7148 7340 7200
rect 7840 7148 7892 7200
rect 10140 7191 10192 7200
rect 10140 7157 10149 7191
rect 10149 7157 10183 7191
rect 10183 7157 10192 7191
rect 10140 7148 10192 7157
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 5632 6944 5684 6996
rect 7748 6944 7800 6996
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 10140 6944 10192 6996
rect 10416 6944 10468 6996
rect 5448 6876 5500 6928
rect 4620 6808 4672 6860
rect 5540 6808 5592 6860
rect 6552 6876 6604 6928
rect 10048 6919 10100 6928
rect 10048 6885 10051 6919
rect 10051 6885 10085 6919
rect 10085 6885 10100 6919
rect 10048 6876 10100 6885
rect 6920 6808 6972 6860
rect 9864 6808 9916 6860
rect 11336 6808 11388 6860
rect 5632 6740 5684 6792
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 6184 6604 6236 6656
rect 7012 6604 7064 6656
rect 8760 6604 8812 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 4344 6400 4396 6452
rect 4620 6400 4672 6452
rect 6552 6443 6604 6452
rect 6552 6409 6561 6443
rect 6561 6409 6595 6443
rect 6595 6409 6604 6443
rect 6552 6400 6604 6409
rect 7748 6400 7800 6452
rect 8300 6400 8352 6452
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 10048 6400 10100 6452
rect 11336 6400 11388 6452
rect 11520 6400 11572 6452
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 10968 6264 11020 6316
rect 3056 6196 3108 6248
rect 5540 6196 5592 6248
rect 6920 6171 6972 6180
rect 6920 6137 6929 6171
rect 6929 6137 6963 6171
rect 6963 6137 6972 6171
rect 6920 6128 6972 6137
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 8760 6128 8812 6137
rect 10416 6171 10468 6180
rect 10416 6137 10425 6171
rect 10425 6137 10459 6171
rect 10459 6137 10468 6171
rect 10968 6171 11020 6180
rect 10416 6128 10468 6137
rect 10968 6137 10977 6171
rect 10977 6137 11011 6171
rect 11011 6137 11020 6171
rect 10968 6128 11020 6137
rect 5632 6103 5684 6112
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 5632 5856 5684 5908
rect 6920 5856 6972 5908
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 5724 5788 5776 5840
rect 7012 5831 7064 5840
rect 7012 5797 7021 5831
rect 7021 5797 7055 5831
rect 7055 5797 7064 5831
rect 7012 5788 7064 5797
rect 7104 5788 7156 5840
rect 8024 5788 8076 5840
rect 8944 5788 8996 5840
rect 10600 5788 10652 5840
rect 5632 5652 5684 5704
rect 6552 5720 6604 5772
rect 10968 5720 11020 5772
rect 11980 5720 12032 5772
rect 6828 5652 6880 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10968 5516 11020 5568
rect 11520 5516 11572 5568
rect 12072 5516 12124 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 6276 5355 6328 5364
rect 6276 5321 6285 5355
rect 6285 5321 6319 5355
rect 6319 5321 6328 5355
rect 6276 5312 6328 5321
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 8024 5312 8076 5364
rect 10600 5312 10652 5364
rect 11980 5312 12032 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 7932 5244 7984 5296
rect 8576 5244 8628 5296
rect 11244 5287 11296 5296
rect 5632 5176 5684 5228
rect 6644 5176 6696 5228
rect 7104 5176 7156 5228
rect 9772 5219 9824 5228
rect 6276 5108 6328 5160
rect 6828 5108 6880 5160
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 7932 5108 7984 5160
rect 8484 5108 8536 5160
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 10140 5176 10192 5228
rect 11244 5253 11253 5287
rect 11253 5253 11287 5287
rect 11287 5253 11296 5287
rect 11244 5244 11296 5253
rect 13452 5244 13504 5296
rect 11244 5108 11296 5160
rect 12900 5108 12952 5160
rect 8392 5083 8444 5092
rect 8392 5049 8401 5083
rect 8401 5049 8435 5083
rect 8435 5049 8444 5083
rect 8392 5040 8444 5049
rect 6092 4972 6144 5024
rect 9956 4972 10008 5024
rect 12440 4972 12492 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 5264 4811 5316 4820
rect 5264 4777 5273 4811
rect 5273 4777 5307 4811
rect 5307 4777 5316 4811
rect 5264 4768 5316 4777
rect 7656 4811 7708 4820
rect 7656 4777 7665 4811
rect 7665 4777 7699 4811
rect 7699 4777 7708 4811
rect 7656 4768 7708 4777
rect 9220 4811 9272 4820
rect 9220 4777 9229 4811
rect 9229 4777 9263 4811
rect 9263 4777 9272 4811
rect 9220 4768 9272 4777
rect 5632 4700 5684 4752
rect 6184 4700 6236 4752
rect 6920 4700 6972 4752
rect 10048 4700 10100 4752
rect 8024 4675 8076 4684
rect 8024 4641 8033 4675
rect 8033 4641 8067 4675
rect 8067 4641 8076 4675
rect 8024 4632 8076 4641
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 12256 4632 12308 4684
rect 13360 4632 13412 4684
rect 8760 4607 8812 4616
rect 8760 4573 8769 4607
rect 8769 4573 8803 4607
rect 8803 4573 8812 4607
rect 8760 4564 8812 4573
rect 10140 4607 10192 4616
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 6184 4428 6236 4480
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10508 4564 10560 4616
rect 13820 4496 13872 4548
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 12164 4428 12216 4480
rect 14648 4428 14700 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 7932 4267 7984 4276
rect 7932 4233 7941 4267
rect 7941 4233 7975 4267
rect 7975 4233 7984 4267
rect 7932 4224 7984 4233
rect 11244 4267 11296 4276
rect 11244 4233 11253 4267
rect 11253 4233 11287 4267
rect 11287 4233 11296 4267
rect 11244 4224 11296 4233
rect 12256 4267 12308 4276
rect 12256 4233 12265 4267
rect 12265 4233 12299 4267
rect 12299 4233 12308 4267
rect 12256 4224 12308 4233
rect 13360 4267 13412 4276
rect 13360 4233 13369 4267
rect 13369 4233 13403 4267
rect 13403 4233 13412 4267
rect 13360 4224 13412 4233
rect 4896 4088 4948 4140
rect 2872 4020 2924 4072
rect 4068 4020 4120 4072
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 5724 4088 5776 4140
rect 6644 4088 6696 4140
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 7748 4088 7800 4140
rect 9680 4131 9732 4140
rect 5080 3952 5132 4004
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 6920 3995 6972 4004
rect 6920 3961 6929 3995
rect 6929 3961 6963 3995
rect 6963 3961 6972 3995
rect 6920 3952 6972 3961
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 10968 4088 11020 4140
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 12532 4020 12584 4072
rect 13544 4063 13596 4072
rect 13544 4029 13588 4063
rect 13588 4029 13596 4063
rect 13544 4020 13596 4029
rect 5540 3884 5592 3936
rect 5632 3884 5684 3936
rect 6092 3884 6144 3936
rect 6736 3884 6788 3936
rect 7748 3884 7800 3936
rect 9496 3884 9548 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 10692 3884 10744 3936
rect 12900 3884 12952 3936
rect 13084 3884 13136 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 8760 3680 8812 3732
rect 10416 3680 10468 3732
rect 12348 3680 12400 3732
rect 6276 3655 6328 3664
rect 6276 3621 6279 3655
rect 6279 3621 6313 3655
rect 6313 3621 6328 3655
rect 6276 3612 6328 3621
rect 7656 3612 7708 3664
rect 8024 3612 8076 3664
rect 8392 3612 8444 3664
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 11428 3655 11480 3664
rect 9864 3612 9916 3621
rect 11428 3621 11437 3655
rect 11437 3621 11471 3655
rect 11471 3621 11480 3655
rect 11428 3612 11480 3621
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 4896 3587 4948 3596
rect 4896 3553 4905 3587
rect 4905 3553 4939 3587
rect 4939 3553 4948 3587
rect 4896 3544 4948 3553
rect 6828 3544 6880 3596
rect 7840 3587 7892 3596
rect 7840 3553 7849 3587
rect 7849 3553 7883 3587
rect 7883 3553 7892 3587
rect 7840 3544 7892 3553
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 13452 3587 13504 3596
rect 13452 3553 13461 3587
rect 13461 3553 13495 3587
rect 13495 3553 13504 3587
rect 13452 3544 13504 3553
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 9956 3476 10008 3528
rect 11060 3476 11112 3528
rect 11796 3476 11848 3528
rect 13084 3476 13136 3528
rect 6184 3408 6236 3460
rect 10048 3408 10100 3460
rect 10968 3408 11020 3460
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 10508 3340 10560 3392
rect 13636 3383 13688 3392
rect 13636 3349 13645 3383
rect 13645 3349 13679 3383
rect 13679 3349 13688 3383
rect 13636 3340 13688 3349
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 5448 3136 5500 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 7748 3179 7800 3188
rect 4620 3068 4672 3120
rect 4896 3068 4948 3120
rect 7748 3145 7757 3179
rect 7757 3145 7791 3179
rect 7791 3145 7800 3179
rect 7748 3136 7800 3145
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 9864 3179 9916 3188
rect 4436 3000 4488 3052
rect 5724 3000 5776 3052
rect 6644 3000 6696 3052
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 388 2864 440 2916
rect 5356 2907 5408 2916
rect 3516 2796 3568 2848
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12716 3136 12768 3188
rect 13268 3136 13320 3188
rect 10968 3111 11020 3120
rect 10968 3077 10977 3111
rect 10977 3077 11011 3111
rect 11011 3077 11020 3111
rect 10968 3068 11020 3077
rect 11336 3068 11388 3120
rect 13452 3111 13504 3120
rect 13452 3077 13461 3111
rect 13461 3077 13495 3111
rect 13495 3077 13504 3111
rect 13452 3068 13504 3077
rect 8760 3000 8812 3052
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 12716 2932 12768 2984
rect 13544 2975 13596 2984
rect 13544 2941 13588 2975
rect 13588 2941 13596 2975
rect 13544 2932 13596 2941
rect 10048 2864 10100 2916
rect 7288 2796 7340 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 4436 2592 4488 2644
rect 5908 2592 5960 2644
rect 6736 2635 6788 2644
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 4252 2499 4304 2508
rect 5264 2524 5316 2576
rect 6000 2567 6052 2576
rect 6000 2533 6009 2567
rect 6009 2533 6043 2567
rect 6043 2533 6052 2567
rect 6000 2524 6052 2533
rect 7104 2592 7156 2644
rect 7840 2592 7892 2644
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 11060 2592 11112 2644
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 10508 2567 10560 2576
rect 10508 2533 10517 2567
rect 10517 2533 10551 2567
rect 10551 2533 10560 2567
rect 10508 2524 10560 2533
rect 4252 2465 4296 2499
rect 4296 2465 4304 2499
rect 4252 2456 4304 2465
rect 5908 2499 5960 2508
rect 5908 2465 5917 2499
rect 5917 2465 5951 2499
rect 5951 2465 5960 2499
rect 5908 2456 5960 2465
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 11244 2456 11296 2508
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 12808 2295 12860 2304
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 12808 2252 12860 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 3700 688 3752 740
rect 4988 688 5040 740
<< metal2 >>
rect 294 39520 350 40000
rect 846 39520 902 40000
rect 1490 39520 1546 40000
rect 2134 39522 2190 40000
rect 2134 39520 2268 39522
rect 2686 39520 2742 40000
rect 3330 39520 3386 40000
rect 3974 39520 4030 40000
rect 4526 39520 4582 40000
rect 5170 39520 5226 40000
rect 5814 39520 5870 40000
rect 6366 39520 6422 40000
rect 7010 39520 7066 40000
rect 7654 39520 7710 40000
rect 8298 39520 8354 40000
rect 8850 39520 8906 40000
rect 9494 39520 9550 40000
rect 10138 39520 10194 40000
rect 10690 39520 10746 40000
rect 11334 39520 11390 40000
rect 11978 39520 12034 40000
rect 12530 39520 12586 40000
rect 13174 39520 13230 40000
rect 13818 39520 13874 40000
rect 14370 39520 14426 40000
rect 15014 39520 15070 40000
rect 15658 39520 15714 40000
rect 308 34785 336 39520
rect 294 34776 350 34785
rect 294 34711 350 34720
rect 860 34649 888 39520
rect 1504 35601 1532 39520
rect 2148 39494 2268 39520
rect 1490 35592 1546 35601
rect 1490 35527 1546 35536
rect 846 34640 902 34649
rect 846 34575 902 34584
rect 2240 22030 2268 39494
rect 2700 27577 2728 39520
rect 3344 35057 3372 39520
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3330 35048 3386 35057
rect 3330 34983 3386 34992
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3146 34776 3202 34785
rect 3622 34768 3918 34788
rect 3988 34762 4016 39520
rect 4540 35136 4568 39520
rect 5184 35714 5212 39520
rect 4448 35108 4568 35136
rect 4632 35686 5212 35714
rect 3988 34734 4384 34762
rect 3146 34711 3202 34720
rect 3056 29708 3108 29714
rect 3056 29650 3108 29656
rect 3068 29073 3096 29650
rect 3160 29209 3188 34711
rect 3514 34640 3570 34649
rect 3514 34575 3570 34584
rect 4158 34640 4214 34649
rect 4158 34575 4214 34584
rect 3146 29200 3202 29209
rect 3146 29135 3202 29144
rect 3054 29064 3110 29073
rect 3054 28999 3056 29008
rect 3108 28999 3110 29008
rect 3056 28970 3108 28976
rect 3160 27690 3188 29135
rect 3528 29102 3556 34575
rect 4172 34542 4200 34575
rect 4160 34536 4212 34542
rect 4160 34478 4212 34484
rect 4066 33960 4122 33969
rect 4066 33895 4122 33904
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3882 33552 3938 33561
rect 3882 33487 3938 33496
rect 3896 33318 3924 33487
rect 4080 33454 4108 33895
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 4250 33416 4306 33425
rect 3884 33312 3936 33318
rect 3884 33254 3936 33260
rect 4080 33114 4108 33390
rect 4250 33351 4306 33360
rect 4068 33108 4120 33114
rect 4068 33050 4120 33056
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 4080 31210 4108 31826
rect 4264 31822 4292 33351
rect 4356 32978 4384 34734
rect 4448 33017 4476 35108
rect 4526 35048 4582 35057
rect 4526 34983 4582 34992
rect 4540 34066 4568 34983
rect 4528 34060 4580 34066
rect 4528 34002 4580 34008
rect 4540 33658 4568 34002
rect 4528 33652 4580 33658
rect 4528 33594 4580 33600
rect 4434 33008 4490 33017
rect 4344 32972 4396 32978
rect 4434 32943 4490 32952
rect 4344 32914 4396 32920
rect 4528 32360 4580 32366
rect 4528 32302 4580 32308
rect 4252 31816 4304 31822
rect 4252 31758 4304 31764
rect 4068 31204 4120 31210
rect 4068 31146 4120 31152
rect 4068 30728 4120 30734
rect 4068 30670 4120 30676
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 4080 30326 4108 30670
rect 4068 30320 4120 30326
rect 4068 30262 4120 30268
rect 4540 29617 4568 32302
rect 4526 29608 4582 29617
rect 4526 29543 4582 29552
rect 4436 29504 4488 29510
rect 4436 29446 4488 29452
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 4448 29170 4476 29446
rect 4436 29164 4488 29170
rect 4436 29106 4488 29112
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 4252 29096 4304 29102
rect 4252 29038 4304 29044
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3884 28008 3936 28014
rect 3936 27968 4016 27996
rect 3884 27950 3936 27956
rect 3516 27872 3568 27878
rect 3516 27814 3568 27820
rect 3068 27662 3188 27690
rect 3528 27674 3556 27814
rect 3516 27668 3568 27674
rect 2686 27568 2742 27577
rect 2686 27503 2742 27512
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2792 23304 2820 24346
rect 2962 24304 3018 24313
rect 2962 24239 2964 24248
rect 3016 24239 3018 24248
rect 2964 24210 3016 24216
rect 2976 23866 3004 24210
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 2608 23276 2820 23304
rect 2608 23186 2636 23276
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2608 22778 2636 23122
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2792 22234 2820 23122
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2780 22228 2832 22234
rect 2780 22170 2832 22176
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 2870 20088 2926 20097
rect 2870 20023 2872 20032
rect 2924 20023 2926 20032
rect 2872 19994 2924 20000
rect 2870 18728 2926 18737
rect 2870 18663 2926 18672
rect 2884 18426 2912 18663
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2884 18222 2912 18362
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2884 16250 2912 16594
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2884 16017 2912 16186
rect 2870 16008 2926 16017
rect 2870 15943 2926 15952
rect 2976 10169 3004 22918
rect 3068 22098 3096 27662
rect 3516 27610 3568 27616
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3988 24750 4016 27968
rect 4160 27532 4212 27538
rect 4160 27474 4212 27480
rect 4172 27130 4200 27474
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 3976 24744 4028 24750
rect 3976 24686 4028 24692
rect 3148 24676 3200 24682
rect 3148 24618 3200 24624
rect 3160 24410 3188 24618
rect 3988 24614 4016 24686
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3148 24404 3200 24410
rect 3148 24346 3200 24352
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3344 23798 3372 24346
rect 4160 24336 4212 24342
rect 4160 24278 4212 24284
rect 4068 24200 4120 24206
rect 3974 24168 4030 24177
rect 4068 24142 4120 24148
rect 3974 24103 4030 24112
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3332 23792 3384 23798
rect 3238 23760 3294 23769
rect 3332 23734 3384 23740
rect 3988 23730 4016 24103
rect 3238 23695 3294 23704
rect 3976 23724 4028 23730
rect 3252 23662 3280 23695
rect 3976 23666 4028 23672
rect 3240 23656 3292 23662
rect 3240 23598 3292 23604
rect 3516 23656 3568 23662
rect 3516 23598 3568 23604
rect 3528 22982 3556 23598
rect 3976 23588 4028 23594
rect 3976 23530 4028 23536
rect 3988 23186 4016 23530
rect 3976 23180 4028 23186
rect 3976 23122 4028 23128
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3146 22536 3202 22545
rect 3146 22471 3148 22480
rect 3200 22471 3202 22480
rect 3424 22500 3476 22506
rect 3148 22442 3200 22448
rect 3424 22442 3476 22448
rect 3436 22234 3464 22442
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3056 22092 3108 22098
rect 3056 22034 3108 22040
rect 3068 21350 3096 22034
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3436 21622 3464 21966
rect 3424 21616 3476 21622
rect 3424 21558 3476 21564
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 2962 10160 3018 10169
rect 2962 10095 3018 10104
rect 3068 6254 3096 21286
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3160 19514 3188 19858
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3146 17776 3202 17785
rect 3146 17711 3148 17720
rect 3200 17711 3202 17720
rect 3148 17682 3200 17688
rect 3160 17338 3188 17682
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3436 15065 3464 21558
rect 3528 21350 3556 22918
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3976 22704 4028 22710
rect 3974 22672 3976 22681
rect 4028 22672 4030 22681
rect 3974 22607 4030 22616
rect 4080 22522 4108 24142
rect 4172 23322 4200 24278
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4172 22817 4200 23258
rect 4158 22808 4214 22817
rect 4158 22743 4214 22752
rect 3896 22506 4108 22522
rect 3884 22500 4108 22506
rect 3936 22494 4108 22500
rect 3884 22442 3936 22448
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18970 4200 19246
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 3974 18864 4030 18873
rect 3974 18799 4030 18808
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3988 18222 4016 18799
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 4080 17202 4108 18294
rect 4264 17490 4292 29038
rect 4436 25220 4488 25226
rect 4436 25162 4488 25168
rect 4344 24744 4396 24750
rect 4342 24712 4344 24721
rect 4396 24712 4398 24721
rect 4342 24647 4398 24656
rect 4448 24410 4476 25162
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4540 24290 4568 29543
rect 4448 24262 4568 24290
rect 4344 24132 4396 24138
rect 4344 24074 4396 24080
rect 4356 23866 4384 24074
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 4448 21026 4476 24262
rect 4528 23180 4580 23186
rect 4528 23122 4580 23128
rect 4540 22438 4568 23122
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4540 22137 4568 22374
rect 4526 22128 4582 22137
rect 4526 22063 4582 22072
rect 4632 21128 4660 35686
rect 5446 35592 5502 35601
rect 5446 35527 5502 35536
rect 5264 34944 5316 34950
rect 5264 34886 5316 34892
rect 5170 34640 5226 34649
rect 5170 34575 5226 34584
rect 5184 34542 5212 34575
rect 5276 34542 5304 34886
rect 5460 34746 5488 35527
rect 5448 34740 5500 34746
rect 5448 34682 5500 34688
rect 5172 34536 5224 34542
rect 5172 34478 5224 34484
rect 5264 34536 5316 34542
rect 5264 34478 5316 34484
rect 5632 34536 5684 34542
rect 5632 34478 5684 34484
rect 5264 33856 5316 33862
rect 5540 33856 5592 33862
rect 5264 33798 5316 33804
rect 5460 33816 5540 33844
rect 5276 33454 5304 33798
rect 5356 33652 5408 33658
rect 5356 33594 5408 33600
rect 5264 33448 5316 33454
rect 5262 33416 5264 33425
rect 5316 33416 5318 33425
rect 5172 33380 5224 33386
rect 5262 33351 5318 33360
rect 5172 33322 5224 33328
rect 4988 32972 5040 32978
rect 4988 32914 5040 32920
rect 5000 32570 5028 32914
rect 5184 32774 5212 33322
rect 5172 32768 5224 32774
rect 5172 32710 5224 32716
rect 4988 32564 5040 32570
rect 4988 32506 5040 32512
rect 5000 31929 5028 32506
rect 5184 32366 5212 32710
rect 5172 32360 5224 32366
rect 5172 32302 5224 32308
rect 4986 31920 5042 31929
rect 4986 31855 5042 31864
rect 5184 31736 5212 32302
rect 5368 31793 5396 33594
rect 5460 33368 5488 33816
rect 5540 33798 5592 33804
rect 5644 33454 5672 34478
rect 5632 33448 5684 33454
rect 5632 33390 5684 33396
rect 5540 33380 5592 33386
rect 5460 33340 5540 33368
rect 5460 33114 5488 33340
rect 5540 33322 5592 33328
rect 5644 33114 5672 33390
rect 5448 33108 5500 33114
rect 5448 33050 5500 33056
rect 5632 33108 5684 33114
rect 5632 33050 5684 33056
rect 5644 32366 5672 33050
rect 5828 32450 5856 39520
rect 6380 37754 6408 39520
rect 6380 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6276 35148 6328 35154
rect 6276 35090 6328 35096
rect 6288 35057 6316 35090
rect 6274 35048 6330 35057
rect 6274 34983 6330 34992
rect 6288 34746 6316 34983
rect 6276 34740 6328 34746
rect 6276 34682 6328 34688
rect 6184 34400 6236 34406
rect 6184 34342 6236 34348
rect 6196 34134 6224 34342
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6184 34128 6236 34134
rect 6184 34070 6236 34076
rect 5908 33992 5960 33998
rect 5908 33934 5960 33940
rect 5920 33522 5948 33934
rect 5908 33516 5960 33522
rect 5908 33458 5960 33464
rect 6196 33318 6224 34070
rect 6184 33312 6236 33318
rect 6184 33254 6236 33260
rect 6196 33046 6224 33254
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6184 33040 6236 33046
rect 6184 32982 6236 32988
rect 6092 32904 6144 32910
rect 6092 32846 6144 32852
rect 5828 32422 5948 32450
rect 5632 32360 5684 32366
rect 5632 32302 5684 32308
rect 5540 32224 5592 32230
rect 5540 32166 5592 32172
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 5354 31784 5410 31793
rect 5184 31708 5304 31736
rect 5354 31719 5410 31728
rect 5172 31272 5224 31278
rect 5172 31214 5224 31220
rect 4896 31136 4948 31142
rect 4896 31078 4948 31084
rect 4908 30870 4936 31078
rect 4896 30864 4948 30870
rect 4896 30806 4948 30812
rect 4908 30394 4936 30806
rect 5184 30598 5212 31214
rect 5172 30592 5224 30598
rect 5172 30534 5224 30540
rect 4896 30388 4948 30394
rect 4896 30330 4948 30336
rect 5184 30122 5212 30534
rect 5080 30116 5132 30122
rect 5080 30058 5132 30064
rect 5172 30116 5224 30122
rect 5172 30058 5224 30064
rect 5092 29850 5120 30058
rect 5080 29844 5132 29850
rect 5080 29786 5132 29792
rect 4804 29776 4856 29782
rect 4724 29724 4804 29730
rect 4724 29718 4856 29724
rect 4724 29702 4844 29718
rect 4724 28966 4752 29702
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4816 29034 4844 29582
rect 5172 29232 5224 29238
rect 5172 29174 5224 29180
rect 5078 29064 5134 29073
rect 4804 29028 4856 29034
rect 5078 28999 5134 29008
rect 4804 28970 4856 28976
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4724 28694 4752 28902
rect 4816 28762 4844 28970
rect 4896 28960 4948 28966
rect 4896 28902 4948 28908
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 4712 28688 4764 28694
rect 4908 28642 4936 28902
rect 4712 28630 4764 28636
rect 4816 28626 4936 28642
rect 4804 28620 4936 28626
rect 4856 28614 4936 28620
rect 4804 28562 4856 28568
rect 4816 28218 4844 28562
rect 4804 28212 4856 28218
rect 4804 28154 4856 28160
rect 4896 28076 4948 28082
rect 4896 28018 4948 28024
rect 4908 27538 4936 28018
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 5000 27674 5028 27950
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 4896 27532 4948 27538
rect 4816 27492 4896 27520
rect 4816 26858 4844 27492
rect 4896 27474 4948 27480
rect 4894 27432 4950 27441
rect 4894 27367 4950 27376
rect 4804 26852 4856 26858
rect 4804 26794 4856 26800
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4724 23730 4752 26726
rect 4908 26450 4936 27367
rect 4988 26920 5040 26926
rect 4988 26862 5040 26868
rect 4896 26444 4948 26450
rect 4896 26386 4948 26392
rect 4908 26042 4936 26386
rect 5000 26314 5028 26862
rect 4988 26308 5040 26314
rect 4988 26250 5040 26256
rect 4896 26036 4948 26042
rect 4896 25978 4948 25984
rect 4896 24676 4948 24682
rect 4896 24618 4948 24624
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4908 23644 4936 24618
rect 4988 23656 5040 23662
rect 4908 23616 4988 23644
rect 4988 23598 5040 23604
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4710 22672 4766 22681
rect 4908 22642 4936 23462
rect 5000 23186 5028 23598
rect 5092 23474 5120 28999
rect 5184 28082 5212 29174
rect 5172 28076 5224 28082
rect 5172 28018 5224 28024
rect 5172 27532 5224 27538
rect 5172 27474 5224 27480
rect 5184 25838 5212 27474
rect 5276 27062 5304 31708
rect 5356 31204 5408 31210
rect 5356 31146 5408 31152
rect 5368 30734 5396 31146
rect 5460 31142 5488 31826
rect 5552 31754 5580 32166
rect 5644 31906 5672 32302
rect 5644 31890 5764 31906
rect 5632 31884 5764 31890
rect 5684 31878 5764 31884
rect 5632 31826 5684 31832
rect 5630 31784 5686 31793
rect 5540 31748 5592 31754
rect 5630 31719 5686 31728
rect 5540 31690 5592 31696
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5644 30802 5672 31719
rect 5736 31482 5764 31878
rect 5920 31804 5948 32422
rect 6000 32360 6052 32366
rect 6000 32302 6052 32308
rect 6012 31958 6040 32302
rect 6104 32298 6132 32846
rect 6092 32292 6144 32298
rect 6092 32234 6144 32240
rect 6104 32026 6132 32234
rect 6196 32230 6224 32982
rect 6184 32224 6236 32230
rect 6184 32166 6236 32172
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6092 32020 6144 32026
rect 6092 31962 6144 31968
rect 6000 31952 6052 31958
rect 6000 31894 6052 31900
rect 5895 31776 5948 31804
rect 5895 31736 5923 31776
rect 6552 31748 6604 31754
rect 5895 31708 5948 31736
rect 5724 31476 5776 31482
rect 5724 31418 5776 31424
rect 5632 30796 5684 30802
rect 5632 30738 5684 30744
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 5368 30258 5396 30670
rect 5448 30660 5500 30666
rect 5448 30602 5500 30608
rect 5356 30252 5408 30258
rect 5356 30194 5408 30200
rect 5356 29844 5408 29850
rect 5356 29786 5408 29792
rect 5368 29578 5396 29786
rect 5356 29572 5408 29578
rect 5356 29514 5408 29520
rect 5368 29170 5396 29514
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 5460 27606 5488 30602
rect 5540 28960 5592 28966
rect 5540 28902 5592 28908
rect 5552 27878 5580 28902
rect 5736 28762 5764 31418
rect 5816 30796 5868 30802
rect 5816 30738 5868 30744
rect 5724 28756 5776 28762
rect 5724 28698 5776 28704
rect 5540 27872 5592 27878
rect 5540 27814 5592 27820
rect 5448 27600 5500 27606
rect 5448 27542 5500 27548
rect 5264 27056 5316 27062
rect 5264 26998 5316 27004
rect 5552 26518 5580 27814
rect 5828 26897 5856 30738
rect 5920 30682 5948 31708
rect 6552 31690 6604 31696
rect 6564 31482 6592 31690
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 6092 31136 6144 31142
rect 6092 31078 6144 31084
rect 6104 30705 6132 31078
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6458 30832 6514 30841
rect 6184 30796 6236 30802
rect 6458 30767 6460 30776
rect 6184 30738 6236 30744
rect 6512 30767 6514 30776
rect 6460 30738 6512 30744
rect 6090 30696 6146 30705
rect 5920 30654 6040 30682
rect 5908 30592 5960 30598
rect 5908 30534 5960 30540
rect 5920 27130 5948 30534
rect 6012 29050 6040 30654
rect 6090 30631 6146 30640
rect 6196 29832 6224 30738
rect 6472 30394 6500 30738
rect 6460 30388 6512 30394
rect 6460 30330 6512 30336
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6196 29804 6408 29832
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6012 29022 6126 29050
rect 6098 29016 6126 29022
rect 6098 28988 6132 29016
rect 6000 27532 6052 27538
rect 6104 27520 6132 28988
rect 6196 28762 6224 29582
rect 6380 29510 6408 29804
rect 6552 29776 6604 29782
rect 6552 29718 6604 29724
rect 6368 29504 6420 29510
rect 6368 29446 6420 29452
rect 6380 29034 6408 29446
rect 6564 29238 6592 29718
rect 6552 29232 6604 29238
rect 6552 29174 6604 29180
rect 6368 29028 6420 29034
rect 6368 28970 6420 28976
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6564 28082 6592 28562
rect 6552 28076 6604 28082
rect 6552 28018 6604 28024
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6052 27492 6132 27520
rect 6000 27474 6052 27480
rect 5908 27124 5960 27130
rect 5908 27066 5960 27072
rect 5814 26888 5870 26897
rect 5814 26823 5870 26832
rect 5540 26512 5592 26518
rect 5540 26454 5592 26460
rect 5828 26330 5856 26823
rect 6012 26790 6040 27474
rect 6184 27464 6236 27470
rect 6184 27406 6236 27412
rect 6196 27130 6224 27406
rect 6184 27124 6236 27130
rect 6184 27066 6236 27072
rect 6092 26852 6144 26858
rect 6092 26794 6144 26800
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 5828 26302 5948 26330
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5172 25832 5224 25838
rect 5172 25774 5224 25780
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 5184 24682 5212 25094
rect 5172 24676 5224 24682
rect 5172 24618 5224 24624
rect 5184 23594 5212 24618
rect 5276 24614 5304 25638
rect 5552 25498 5580 26182
rect 5828 25838 5856 26182
rect 5816 25832 5868 25838
rect 5816 25774 5868 25780
rect 5828 25498 5856 25774
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5816 25492 5868 25498
rect 5816 25434 5868 25440
rect 5828 25362 5856 25434
rect 5816 25356 5868 25362
rect 5816 25298 5868 25304
rect 5448 25220 5500 25226
rect 5448 25162 5500 25168
rect 5460 24886 5488 25162
rect 5448 24880 5500 24886
rect 5446 24848 5448 24857
rect 5500 24848 5502 24857
rect 5446 24783 5502 24792
rect 5356 24744 5408 24750
rect 5356 24686 5408 24692
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5368 24410 5396 24686
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5724 24268 5776 24274
rect 5724 24210 5776 24216
rect 5736 24177 5764 24210
rect 5722 24168 5778 24177
rect 5540 24132 5592 24138
rect 5722 24103 5778 24112
rect 5540 24074 5592 24080
rect 5552 23730 5580 24074
rect 5828 24070 5856 25298
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 5724 23656 5776 23662
rect 5724 23598 5776 23604
rect 5172 23588 5224 23594
rect 5172 23530 5224 23536
rect 5092 23446 5212 23474
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 4710 22607 4766 22616
rect 4896 22636 4948 22642
rect 4724 21554 4752 22607
rect 4896 22578 4948 22584
rect 4908 22234 4936 22578
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4816 21418 4844 21830
rect 5000 21690 5028 21966
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4804 21412 4856 21418
rect 4804 21354 4856 21360
rect 4632 21100 4752 21128
rect 4448 20998 4660 21026
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4448 20602 4476 20878
rect 4436 20596 4488 20602
rect 4488 20556 4568 20584
rect 4436 20538 4488 20544
rect 4540 20330 4568 20556
rect 4528 20324 4580 20330
rect 4528 20266 4580 20272
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4356 18193 4384 19110
rect 4342 18184 4398 18193
rect 4342 18119 4398 18128
rect 4264 17462 4384 17490
rect 4250 17368 4306 17377
rect 4250 17303 4252 17312
rect 4304 17303 4306 17312
rect 4252 17274 4304 17280
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4264 17134 4292 17274
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3988 16250 4016 16934
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4080 16674 4108 16730
rect 4080 16646 4200 16674
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3988 16046 4016 16186
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3988 15473 4016 15982
rect 3974 15464 4030 15473
rect 3974 15399 4030 15408
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3422 15056 3478 15065
rect 3422 14991 3478 15000
rect 3436 14006 3464 14991
rect 4172 14958 4200 16646
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4066 14376 4122 14385
rect 4066 14311 4122 14320
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 4080 14074 4108 14311
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4068 13864 4120 13870
rect 4066 13832 4068 13841
rect 4120 13832 4122 13841
rect 4066 13767 4122 13776
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 4080 10810 4108 11154
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 4080 6769 4108 8774
rect 4066 6760 4122 6769
rect 4066 6695 4122 6704
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 4068 4072 4120 4078
rect 4172 4060 4200 13874
rect 4264 13462 4292 14214
rect 4356 13546 4384 17462
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4434 14512 4490 14521
rect 4434 14447 4490 14456
rect 4448 14074 4476 14447
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4356 13518 4476 13546
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4344 13456 4396 13462
rect 4448 13433 4476 13518
rect 4344 13398 4396 13404
rect 4434 13424 4490 13433
rect 4264 12986 4292 13398
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4356 12918 4384 13398
rect 4434 13359 4490 13368
rect 4540 13308 4568 14758
rect 4448 13280 4568 13308
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8634 4384 8978
rect 4448 8922 4476 13280
rect 4526 10160 4582 10169
rect 4526 10095 4528 10104
rect 4580 10095 4582 10104
rect 4528 10066 4580 10072
rect 4540 9722 4568 10066
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4528 8968 4580 8974
rect 4448 8916 4528 8922
rect 4448 8910 4580 8916
rect 4448 8894 4568 8910
rect 4448 8634 4476 8894
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4632 6866 4660 20998
rect 4724 20369 4752 21100
rect 4816 21010 4844 21354
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 4816 20602 4844 20946
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 5000 20534 5028 21490
rect 4988 20528 5040 20534
rect 4988 20470 5040 20476
rect 4710 20360 4766 20369
rect 4710 20295 4766 20304
rect 4724 12306 4752 20295
rect 5000 19990 5028 20470
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4908 19378 4936 19858
rect 4988 19848 5040 19854
rect 4986 19816 4988 19825
rect 5040 19816 5042 19825
rect 4986 19751 5042 19760
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 5000 18834 5028 19751
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4816 18358 4844 18634
rect 5000 18426 5028 18770
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5092 17746 5120 18022
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 16250 4844 16526
rect 4908 16454 4936 17478
rect 5092 17338 5120 17682
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 5078 14920 5134 14929
rect 5078 14855 5134 14864
rect 5092 14482 5120 14855
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5092 14074 5120 14418
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5000 12850 5028 13330
rect 5078 13288 5134 13297
rect 5078 13223 5134 13232
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5000 12442 5028 12786
rect 5092 12782 5120 13223
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4724 11830 4752 12242
rect 5184 11914 5212 23446
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 5264 22500 5316 22506
rect 5264 22442 5316 22448
rect 5276 22166 5304 22442
rect 5552 22166 5580 23258
rect 5632 23044 5684 23050
rect 5632 22986 5684 22992
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5276 21690 5304 22102
rect 5644 21962 5672 22986
rect 5736 22114 5764 23598
rect 5828 23225 5856 24006
rect 5920 23322 5948 26302
rect 6104 25906 6132 26794
rect 6092 25900 6144 25906
rect 6092 25842 6144 25848
rect 6092 25356 6144 25362
rect 6092 25298 6144 25304
rect 6000 24676 6052 24682
rect 6000 24618 6052 24624
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5814 23216 5870 23225
rect 5814 23151 5870 23160
rect 5908 23180 5960 23186
rect 5908 23122 5960 23128
rect 5814 22808 5870 22817
rect 5920 22778 5948 23122
rect 5814 22743 5816 22752
rect 5868 22743 5870 22752
rect 5908 22772 5960 22778
rect 5816 22714 5868 22720
rect 5908 22714 5960 22720
rect 5828 22234 5856 22714
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5736 22086 5856 22114
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5540 20324 5592 20330
rect 5540 20266 5592 20272
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 19446 5304 19654
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5276 18834 5304 19246
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5460 18766 5488 19110
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5276 17202 5304 17750
rect 5368 17338 5396 18090
rect 5460 17542 5488 18158
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5276 15638 5304 17138
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5446 16688 5502 16697
rect 5368 16046 5396 16662
rect 5446 16623 5448 16632
rect 5500 16623 5502 16632
rect 5448 16594 5500 16600
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5368 15706 5396 15982
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5262 15328 5318 15337
rect 5262 15263 5318 15272
rect 5276 14958 5304 15263
rect 5460 15162 5488 15574
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5276 14618 5304 14758
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5276 13938 5304 14554
rect 5552 13954 5580 20266
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5644 17134 5672 19110
rect 5828 18834 5856 22086
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 18358 5856 18566
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5920 17762 5948 21286
rect 6012 18465 6040 24618
rect 6104 23186 6132 25298
rect 6196 25294 6224 27066
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6460 26444 6512 26450
rect 6460 26386 6512 26392
rect 6472 26042 6500 26386
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6184 25288 6236 25294
rect 6184 25230 6236 25236
rect 6196 24138 6224 25230
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6184 24132 6236 24138
rect 6184 24074 6236 24080
rect 6196 23633 6224 24074
rect 6182 23624 6238 23633
rect 6182 23559 6238 23568
rect 6196 23304 6224 23559
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6196 23276 6316 23304
rect 6288 23186 6316 23276
rect 6092 23180 6144 23186
rect 6276 23180 6328 23186
rect 6144 23140 6224 23168
rect 6092 23122 6144 23128
rect 6092 22636 6144 22642
rect 6092 22578 6144 22584
rect 6104 21010 6132 22578
rect 6196 22166 6224 23140
rect 6276 23122 6328 23128
rect 6288 22778 6316 23122
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6196 20058 6224 22102
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6380 20330 6408 20946
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6564 20602 6592 20878
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6092 19712 6144 19718
rect 6092 19654 6144 19660
rect 6104 19378 6132 19654
rect 6288 19514 6316 19790
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6104 18970 6132 19314
rect 6656 19174 6684 37726
rect 6920 36304 6972 36310
rect 6920 36246 6972 36252
rect 6932 35850 6960 36246
rect 6748 35822 6960 35850
rect 6748 35494 6776 35822
rect 7024 35714 7052 39520
rect 7196 36576 7248 36582
rect 7196 36518 7248 36524
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 7208 36174 7236 36518
rect 7196 36168 7248 36174
rect 7196 36110 7248 36116
rect 7208 35834 7236 36110
rect 7196 35828 7248 35834
rect 7196 35770 7248 35776
rect 6920 35692 6972 35698
rect 7024 35686 7236 35714
rect 6920 35634 6972 35640
rect 6932 35601 6960 35634
rect 6918 35592 6974 35601
rect 6918 35527 6974 35536
rect 7012 35556 7064 35562
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 6748 34066 6776 35430
rect 6932 35290 6960 35527
rect 7012 35498 7064 35504
rect 6920 35284 6972 35290
rect 6920 35226 6972 35232
rect 7024 35222 7052 35498
rect 7012 35216 7064 35222
rect 7012 35158 7064 35164
rect 7024 34746 7052 35158
rect 7012 34740 7064 34746
rect 7012 34682 7064 34688
rect 6828 34536 6880 34542
rect 6880 34496 6960 34524
rect 6828 34478 6880 34484
rect 6932 34202 6960 34496
rect 6920 34196 6972 34202
rect 6920 34138 6972 34144
rect 7024 34134 7052 34682
rect 7012 34128 7064 34134
rect 7012 34070 7064 34076
rect 6736 34060 6788 34066
rect 6736 34002 6788 34008
rect 7012 33380 7064 33386
rect 7012 33322 7064 33328
rect 7024 32774 7052 33322
rect 7012 32768 7064 32774
rect 7012 32710 7064 32716
rect 7024 31958 7052 32710
rect 7104 32224 7156 32230
rect 7104 32166 7156 32172
rect 7012 31952 7064 31958
rect 7012 31894 7064 31900
rect 7024 31482 7052 31894
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6840 30025 6868 30126
rect 6826 30016 6882 30025
rect 6826 29951 6882 29960
rect 6736 28620 6788 28626
rect 6736 28562 6788 28568
rect 6748 27674 6776 28562
rect 6840 28558 6868 29951
rect 7024 29102 7052 30874
rect 7116 30598 7144 32166
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 7116 30122 7144 30534
rect 7104 30116 7156 30122
rect 7104 30058 7156 30064
rect 7116 29782 7144 30058
rect 7104 29776 7156 29782
rect 7104 29718 7156 29724
rect 7012 29096 7064 29102
rect 6932 29056 7012 29084
rect 6828 28552 6880 28558
rect 6828 28494 6880 28500
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6840 27878 6868 28018
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6736 27668 6788 27674
rect 6736 27610 6788 27616
rect 6748 27130 6776 27610
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6840 27010 6868 27814
rect 6748 26982 6868 27010
rect 6748 23497 6776 26982
rect 6828 26308 6880 26314
rect 6828 26250 6880 26256
rect 6840 25514 6868 26250
rect 6932 25838 6960 29056
rect 7012 29038 7064 29044
rect 7208 26874 7236 35686
rect 7300 35601 7328 36518
rect 7286 35592 7342 35601
rect 7286 35527 7342 35536
rect 7300 29209 7328 35527
rect 7472 35488 7524 35494
rect 7472 35430 7524 35436
rect 7484 34649 7512 35430
rect 7470 34640 7526 34649
rect 7470 34575 7526 34584
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7392 32366 7420 32710
rect 7380 32360 7432 32366
rect 7380 32302 7432 32308
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7286 29200 7342 29209
rect 7392 29170 7420 29582
rect 7286 29135 7342 29144
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7288 29096 7340 29102
rect 7288 29038 7340 29044
rect 7300 28694 7328 29038
rect 7288 28688 7340 28694
rect 7288 28630 7340 28636
rect 7288 28008 7340 28014
rect 7288 27950 7340 27956
rect 7300 27606 7328 27950
rect 7484 27946 7512 34575
rect 7576 33425 7604 36518
rect 7562 33416 7618 33425
rect 7562 33351 7618 33360
rect 7472 27940 7524 27946
rect 7472 27882 7524 27888
rect 7288 27600 7340 27606
rect 7288 27542 7340 27548
rect 7576 27538 7604 33351
rect 7668 27962 7696 39520
rect 8312 36666 8340 39520
rect 8576 37324 8628 37330
rect 8576 37266 8628 37272
rect 8588 36718 8616 37266
rect 8576 36712 8628 36718
rect 8312 36638 8524 36666
rect 8576 36654 8628 36660
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 7748 36100 7800 36106
rect 7748 36042 7800 36048
rect 7760 35766 7788 36042
rect 7748 35760 7800 35766
rect 7748 35702 7800 35708
rect 8298 35728 8354 35737
rect 7760 32910 7788 35702
rect 8298 35663 8354 35672
rect 8312 35154 8340 35663
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 7840 34128 7892 34134
rect 7840 34070 7892 34076
rect 7852 33658 7880 34070
rect 7944 33998 7972 35022
rect 8312 34746 8340 35090
rect 8300 34740 8352 34746
rect 8300 34682 8352 34688
rect 7932 33992 7984 33998
rect 7932 33934 7984 33940
rect 7840 33652 7892 33658
rect 7840 33594 7892 33600
rect 7944 33522 7972 33934
rect 8300 33924 8352 33930
rect 8300 33866 8352 33872
rect 8208 33856 8260 33862
rect 8208 33798 8260 33804
rect 7932 33516 7984 33522
rect 7932 33458 7984 33464
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 7760 32026 7788 32846
rect 7944 32026 7972 33458
rect 8024 33040 8076 33046
rect 8024 32982 8076 32988
rect 8036 32570 8064 32982
rect 8024 32564 8076 32570
rect 8024 32506 8076 32512
rect 8220 32298 8248 33798
rect 8312 33114 8340 33866
rect 8404 33658 8432 36518
rect 8496 35714 8524 36638
rect 8588 36038 8616 36654
rect 8576 36032 8628 36038
rect 8576 35974 8628 35980
rect 8864 35714 8892 39520
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9508 35714 9536 39520
rect 9772 36236 9824 36242
rect 9772 36178 9824 36184
rect 9588 36032 9640 36038
rect 9588 35974 9640 35980
rect 8496 35686 8616 35714
rect 8484 34740 8536 34746
rect 8484 34682 8536 34688
rect 8392 33652 8444 33658
rect 8392 33594 8444 33600
rect 8300 33108 8352 33114
rect 8300 33050 8352 33056
rect 8300 32904 8352 32910
rect 8300 32846 8352 32852
rect 8208 32292 8260 32298
rect 8208 32234 8260 32240
rect 7748 32020 7800 32026
rect 7748 31962 7800 31968
rect 7932 32020 7984 32026
rect 7932 31962 7984 31968
rect 7944 31346 7972 31962
rect 8312 31414 8340 32846
rect 8300 31408 8352 31414
rect 8300 31350 8352 31356
rect 7932 31340 7984 31346
rect 7932 31282 7984 31288
rect 7748 31204 7800 31210
rect 7748 31146 7800 31152
rect 7760 30598 7788 31146
rect 7840 30864 7892 30870
rect 7840 30806 7892 30812
rect 7748 30592 7800 30598
rect 7748 30534 7800 30540
rect 7760 30394 7788 30534
rect 7748 30388 7800 30394
rect 7748 30330 7800 30336
rect 7852 29850 7880 30806
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 8114 30696 8170 30705
rect 8036 30394 8064 30670
rect 8312 30666 8340 31350
rect 8114 30631 8170 30640
rect 8300 30660 8352 30666
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 8036 29850 8064 30330
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 8024 28620 8076 28626
rect 8024 28562 8076 28568
rect 8036 28082 8064 28562
rect 8024 28076 8076 28082
rect 8024 28018 8076 28024
rect 7668 27934 7880 27962
rect 7656 27872 7708 27878
rect 7656 27814 7708 27820
rect 7380 27532 7432 27538
rect 7380 27474 7432 27480
rect 7564 27532 7616 27538
rect 7564 27474 7616 27480
rect 7024 26846 7236 26874
rect 6920 25832 6972 25838
rect 6920 25774 6972 25780
rect 6840 25498 6960 25514
rect 6840 25492 6972 25498
rect 6840 25486 6920 25492
rect 6920 25434 6972 25440
rect 6932 24970 6960 25434
rect 6840 24954 6960 24970
rect 6840 24948 6972 24954
rect 6840 24942 6920 24948
rect 6840 24410 6868 24942
rect 6920 24890 6972 24896
rect 6918 24848 6974 24857
rect 6918 24783 6974 24792
rect 6932 24750 6960 24783
rect 6920 24744 6972 24750
rect 6920 24686 6972 24692
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 6828 24132 6880 24138
rect 6828 24074 6880 24080
rect 6840 23866 6868 24074
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6734 23488 6790 23497
rect 6734 23423 6790 23432
rect 6748 22642 6776 23423
rect 6840 23322 6868 23802
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6840 22522 6868 23122
rect 6748 22494 6868 22522
rect 6920 22500 6972 22506
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6196 18766 6224 19110
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 5998 18456 6054 18465
rect 5998 18391 6054 18400
rect 6196 17882 6224 18702
rect 6288 18426 6316 18770
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 5920 17734 6224 17762
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5644 16046 5672 16390
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5644 15638 5672 15982
rect 5632 15632 5684 15638
rect 5632 15574 5684 15580
rect 5644 14958 5672 15574
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5368 13926 5580 13954
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5276 13530 5304 13738
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5276 12442 5304 12650
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5092 11886 5212 11914
rect 5368 11898 5396 13926
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5552 13546 5580 13806
rect 5460 13518 5580 13546
rect 5460 13462 5488 13518
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5460 12714 5488 13398
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5644 12442 5672 13262
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5356 11892 5408 11898
rect 4712 11824 4764 11830
rect 5092 11801 5120 11886
rect 5356 11834 5408 11840
rect 5172 11824 5224 11830
rect 4712 11766 4764 11772
rect 5078 11792 5134 11801
rect 5172 11766 5224 11772
rect 5078 11727 5134 11736
rect 5092 11676 5120 11727
rect 5000 11648 5120 11676
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4816 10810 4844 11154
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9178 4752 9862
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 8634 4844 10746
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5000 7290 5028 11648
rect 5078 7984 5134 7993
rect 5078 7919 5080 7928
rect 5132 7919 5134 7928
rect 5080 7890 5132 7896
rect 5092 7478 5120 7890
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 5000 7262 5120 7290
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4632 6458 4660 6802
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4120 4032 4200 4060
rect 4068 4014 4120 4020
rect 2042 3088 2098 3097
rect 2042 3023 2098 3032
rect 388 2916 440 2922
rect 388 2858 440 2864
rect 400 480 428 2858
rect 1214 2816 1270 2825
rect 1214 2751 1270 2760
rect 1228 480 1256 2751
rect 2056 480 2084 3023
rect 2884 480 2912 4014
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3700 2984 3752 2990
rect 3698 2952 3700 2961
rect 3752 2952 3754 2961
rect 3698 2887 3754 2896
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 4250 2816 4306 2825
rect 3528 2553 3556 2790
rect 4250 2751 4306 2760
rect 3514 2544 3570 2553
rect 4264 2514 4292 2751
rect 3514 2479 3570 2488
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3700 740 3752 746
rect 3700 682 3752 688
rect 3712 480 3740 682
rect 4356 626 4384 6394
rect 5092 5012 5120 7262
rect 5184 5273 5212 11766
rect 5368 11082 5396 11834
rect 5644 11558 5672 12174
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5644 11014 5672 11494
rect 5736 11354 5764 17478
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 5828 17105 5856 17206
rect 5814 17096 5870 17105
rect 5814 17031 5870 17040
rect 6000 17060 6052 17066
rect 5828 16794 5856 17031
rect 6000 17002 6052 17008
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5920 16726 5948 16934
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5828 15502 5856 15914
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 14618 5856 15438
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5828 12918 5856 13262
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5920 12730 5948 16662
rect 5828 12702 5948 12730
rect 5828 11898 5856 12702
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5368 10674 5580 10690
rect 5368 10668 5592 10674
rect 5368 10662 5540 10668
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5276 10266 5304 10474
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5368 10146 5396 10662
rect 5540 10610 5592 10616
rect 5736 10554 5764 11290
rect 5828 11218 5856 11834
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5460 10538 5764 10554
rect 5448 10532 5764 10538
rect 5500 10526 5764 10532
rect 5448 10474 5500 10480
rect 5276 10118 5396 10146
rect 5276 9042 5304 10118
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5552 9178 5580 9998
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5632 9104 5684 9110
rect 5828 9058 5856 11018
rect 5632 9046 5684 9052
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5644 8430 5672 9046
rect 5736 9042 5856 9058
rect 5724 9036 5856 9042
rect 5776 9030 5856 9036
rect 5724 8978 5776 8984
rect 5828 8634 5856 9030
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5644 7954 5672 8366
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5446 7440 5502 7449
rect 5446 7375 5502 7384
rect 5460 7342 5488 7375
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5460 6934 5488 7278
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5552 6866 5580 7686
rect 5644 7546 5672 7890
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5644 7342 5672 7482
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 7002 5672 7278
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5644 6882 5672 6938
rect 5540 6860 5592 6866
rect 5644 6854 5764 6882
rect 5540 6802 5592 6808
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5170 5264 5226 5273
rect 5170 5199 5226 5208
rect 5262 5128 5318 5137
rect 5262 5063 5318 5072
rect 5092 4984 5212 5012
rect 4618 4312 4674 4321
rect 4618 4247 4674 4256
rect 4632 3602 4660 4247
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3602 4936 4082
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4632 3126 4660 3538
rect 4908 3126 4936 3538
rect 4986 3224 5042 3233
rect 4986 3159 5042 3168
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4448 2650 4476 2994
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 5000 746 5028 3159
rect 5092 2281 5120 3946
rect 5184 3890 5212 4984
rect 5276 4826 5304 5063
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5276 4078 5304 4762
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5552 3942 5580 6190
rect 5644 6118 5672 6734
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5914 5672 6054
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5736 5846 5764 6854
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5370 5672 5646
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5644 4758 5672 5170
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5644 3942 5672 4694
rect 5736 4146 5764 5782
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5540 3936 5592 3942
rect 5184 3862 5304 3890
rect 5540 3878 5592 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5276 2582 5304 3862
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5446 3360 5502 3369
rect 5368 2922 5396 3334
rect 5446 3295 5502 3304
rect 5460 3194 5488 3295
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5354 2816 5410 2825
rect 5354 2751 5410 2760
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 5078 2272 5134 2281
rect 5078 2207 5134 2216
rect 4988 740 5040 746
rect 4988 682 5040 688
rect 4356 598 4568 626
rect 4540 480 4568 598
rect 5368 480 5396 2751
rect 5552 2145 5580 3878
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5736 3058 5764 3334
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5538 2136 5594 2145
rect 5538 2071 5594 2080
rect 5828 1850 5856 8366
rect 5920 7562 5948 12582
rect 6012 12322 6040 17002
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 6104 13462 6132 15302
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6104 12986 6132 13398
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6104 12458 6132 12922
rect 6196 12646 6224 17734
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6564 15978 6592 16594
rect 6552 15972 6604 15978
rect 6552 15914 6604 15920
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6656 15609 6684 18702
rect 6642 15600 6698 15609
rect 6642 15535 6698 15544
rect 6642 15464 6698 15473
rect 6642 15399 6698 15408
rect 6656 14822 6684 15399
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6460 14408 6512 14414
rect 6458 14376 6460 14385
rect 6512 14376 6514 14385
rect 6514 14334 6592 14362
rect 6458 14311 6514 14320
rect 6564 13818 6592 14334
rect 6656 14074 6684 14486
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6564 13790 6684 13818
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6656 13530 6684 13790
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6748 12458 6776 22494
rect 6920 22442 6972 22448
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 6840 22234 6868 22374
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6932 22166 6960 22442
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6840 21350 6868 22034
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6840 19174 6868 19994
rect 7024 19854 7052 26846
rect 7392 26790 7420 27474
rect 7104 26784 7156 26790
rect 7104 26726 7156 26732
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7116 25430 7144 26726
rect 7196 26444 7248 26450
rect 7196 26386 7248 26392
rect 7104 25424 7156 25430
rect 7104 25366 7156 25372
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 7116 24177 7144 24618
rect 7208 24562 7236 26386
rect 7288 25356 7340 25362
rect 7288 25298 7340 25304
rect 7300 24954 7328 25298
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 7208 24534 7328 24562
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 7208 24313 7236 24346
rect 7194 24304 7250 24313
rect 7194 24239 7250 24248
rect 7102 24168 7158 24177
rect 7102 24103 7158 24112
rect 7300 23798 7328 24534
rect 7288 23792 7340 23798
rect 7286 23760 7288 23769
rect 7340 23760 7342 23769
rect 7286 23695 7342 23704
rect 7300 23322 7328 23695
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18902 6868 19110
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6932 18834 6960 19178
rect 7024 18970 7052 19790
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 7024 18698 7052 18906
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 6840 17882 6868 18634
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7024 17338 7052 17614
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7116 17105 7144 22714
rect 7288 22704 7340 22710
rect 7194 22672 7250 22681
rect 7288 22646 7340 22652
rect 7194 22607 7196 22616
rect 7248 22607 7250 22616
rect 7196 22578 7248 22584
rect 7300 22234 7328 22646
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7194 21992 7250 22001
rect 7194 21927 7250 21936
rect 7208 21078 7236 21927
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7300 20913 7328 21286
rect 7392 21078 7420 26726
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7576 24274 7604 24754
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 7576 23730 7604 24210
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7576 23322 7604 23666
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7576 21962 7604 23258
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7668 21486 7696 27814
rect 7852 26466 7880 27934
rect 7932 26920 7984 26926
rect 7932 26862 7984 26868
rect 7760 26450 7880 26466
rect 7748 26444 7880 26450
rect 7800 26438 7880 26444
rect 7748 26386 7800 26392
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 7746 24848 7802 24857
rect 7746 24783 7748 24792
rect 7800 24783 7802 24792
rect 7748 24754 7800 24760
rect 7852 24698 7880 25094
rect 7760 24670 7880 24698
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 21146 7696 21422
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7380 21072 7432 21078
rect 7380 21014 7432 21020
rect 7286 20904 7342 20913
rect 7286 20839 7342 20848
rect 7668 20074 7696 21082
rect 7760 20330 7788 24670
rect 7838 24304 7894 24313
rect 7838 24239 7840 24248
rect 7892 24239 7894 24248
rect 7840 24210 7892 24216
rect 7852 23662 7880 24210
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7668 20046 7788 20074
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7194 18320 7250 18329
rect 7194 18255 7250 18264
rect 7208 18222 7236 18255
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7208 17542 7236 18158
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7102 17096 7158 17105
rect 7102 17031 7158 17040
rect 6826 16824 6882 16833
rect 6826 16759 6828 16768
rect 6880 16759 6882 16768
rect 6828 16730 6880 16736
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6840 15026 6868 15642
rect 7116 15570 7144 15914
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6104 12430 6224 12458
rect 6196 12374 6224 12430
rect 6656 12430 6776 12458
rect 6840 13920 6868 14758
rect 7116 14618 7144 15506
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6920 13932 6972 13938
rect 6840 13892 6920 13920
rect 6184 12368 6236 12374
rect 6012 12294 6132 12322
rect 6184 12310 6236 12316
rect 6104 11778 6132 12294
rect 6196 11898 6224 12310
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6104 11750 6224 11778
rect 6092 11688 6144 11694
rect 6090 11656 6092 11665
rect 6144 11656 6146 11665
rect 6090 11591 6146 11600
rect 6104 11370 6132 11591
rect 6012 11342 6132 11370
rect 6196 11354 6224 11750
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6184 11348 6236 11354
rect 6012 8430 6040 11342
rect 6184 11290 6236 11296
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 11121 6592 11154
rect 6550 11112 6606 11121
rect 6550 11047 6606 11056
rect 6564 10810 6592 11047
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6288 9722 6316 10134
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6288 9450 6316 9658
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9042 6224 9318
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5920 7534 6040 7562
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5920 3534 5948 3946
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5920 2650 5948 3470
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6012 2582 6040 7534
rect 6104 7410 6132 7822
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6196 7206 6224 7958
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 6662 6224 7142
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6564 6458 6592 6870
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6274 5400 6330 5409
rect 6564 5370 6592 5714
rect 6274 5335 6276 5344
rect 6328 5335 6330 5344
rect 6552 5364 6604 5370
rect 6276 5306 6328 5312
rect 6552 5306 6604 5312
rect 6288 5166 6316 5306
rect 6656 5234 6684 12430
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10266 6776 11154
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6276 5160 6328 5166
rect 6748 5137 6776 10202
rect 6840 5710 6868 13892
rect 6920 13874 6972 13880
rect 6918 13832 6974 13841
rect 7024 13802 7052 14010
rect 6918 13767 6920 13776
rect 6972 13767 6974 13776
rect 7012 13796 7064 13802
rect 6920 13738 6972 13744
rect 7012 13738 7064 13744
rect 6932 13530 6960 13738
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7116 12442 7144 14350
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 11354 7144 12378
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7116 10674 7144 11290
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 10130 7052 10474
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9178 6960 9318
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7024 9042 7052 9454
rect 7208 9217 7236 17478
rect 7300 17270 7328 17682
rect 7392 17338 7420 18090
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7288 17264 7340 17270
rect 7288 17206 7340 17212
rect 7392 17134 7420 17274
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7392 16658 7420 17070
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7392 16250 7420 16594
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7484 14498 7512 19314
rect 7668 19310 7696 19858
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 18873 7604 19178
rect 7562 18864 7618 18873
rect 7562 18799 7618 18808
rect 7760 15978 7788 20046
rect 7852 19938 7880 23462
rect 7944 23186 7972 26862
rect 8128 26450 8156 30631
rect 8300 30602 8352 30608
rect 8312 30190 8340 30602
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8392 30048 8444 30054
rect 8390 30016 8392 30025
rect 8444 30016 8446 30025
rect 8390 29951 8446 29960
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8312 27470 8340 28970
rect 8392 28960 8444 28966
rect 8392 28902 8444 28908
rect 8404 27946 8432 28902
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8300 27464 8352 27470
rect 8300 27406 8352 27412
rect 8404 26926 8432 27474
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8116 26444 8168 26450
rect 8116 26386 8168 26392
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 7944 22778 7972 23122
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7944 22166 7972 22374
rect 7932 22160 7984 22166
rect 7932 22102 7984 22108
rect 7944 21690 7972 22102
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7852 19910 7972 19938
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7852 17377 7880 19790
rect 7944 19378 7972 19910
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7944 18426 7972 19178
rect 8036 19145 8064 25774
rect 8128 25158 8156 26386
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8220 23866 8248 24754
rect 8298 24712 8354 24721
rect 8298 24647 8354 24656
rect 8312 24274 8340 24647
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8312 23322 8340 24210
rect 8496 24154 8524 34682
rect 8588 24818 8616 35686
rect 8680 35686 8892 35714
rect 9324 35686 9536 35714
rect 8680 30841 8708 35686
rect 8760 35488 8812 35494
rect 8760 35430 8812 35436
rect 8772 34610 8800 35430
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8760 34604 8812 34610
rect 8760 34546 8812 34552
rect 9036 34468 9088 34474
rect 9036 34410 9088 34416
rect 9048 34134 9076 34410
rect 9036 34128 9088 34134
rect 9036 34070 9088 34076
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8758 33008 8814 33017
rect 8758 32943 8814 32952
rect 8772 31890 8800 32943
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8850 32328 8906 32337
rect 8850 32263 8906 32272
rect 8760 31884 8812 31890
rect 8760 31826 8812 31832
rect 8772 31142 8800 31826
rect 8760 31136 8812 31142
rect 8760 31078 8812 31084
rect 8666 30832 8722 30841
rect 8666 30767 8722 30776
rect 8680 28529 8708 30767
rect 8666 28520 8722 28529
rect 8666 28455 8722 28464
rect 8680 28150 8708 28455
rect 8668 28144 8720 28150
rect 8668 28086 8720 28092
rect 8772 26489 8800 31078
rect 8864 30326 8892 32263
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 9036 31272 9088 31278
rect 9036 31214 9088 31220
rect 9048 30938 9076 31214
rect 9036 30932 9088 30938
rect 9036 30874 9088 30880
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8852 30320 8904 30326
rect 8852 30262 8904 30268
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 9324 27962 9352 35686
rect 9496 35624 9548 35630
rect 9600 35578 9628 35974
rect 9548 35572 9628 35578
rect 9496 35566 9628 35572
rect 9508 35550 9628 35566
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9416 34202 9444 35022
rect 9404 34196 9456 34202
rect 9404 34138 9456 34144
rect 9508 33969 9536 35550
rect 9784 35494 9812 36178
rect 9772 35488 9824 35494
rect 9772 35430 9824 35436
rect 9784 35193 9812 35430
rect 9864 35216 9916 35222
rect 9770 35184 9826 35193
rect 9864 35158 9916 35164
rect 9770 35119 9826 35128
rect 9876 34542 9904 35158
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9680 33992 9732 33998
rect 9494 33960 9550 33969
rect 9680 33934 9732 33940
rect 9494 33895 9550 33904
rect 9508 31686 9536 33895
rect 9692 33114 9720 33934
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9588 32904 9640 32910
rect 9588 32846 9640 32852
rect 9600 32230 9628 32846
rect 9588 32224 9640 32230
rect 9588 32166 9640 32172
rect 9600 32026 9628 32166
rect 9692 32026 9720 33050
rect 9876 32298 9904 34478
rect 10152 34134 10180 39520
rect 10704 36378 10732 39520
rect 10966 36952 11022 36961
rect 10966 36887 10968 36896
rect 11020 36887 11022 36896
rect 10968 36858 11020 36864
rect 11152 36576 11204 36582
rect 11152 36518 11204 36524
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 10232 35624 10284 35630
rect 10230 35592 10232 35601
rect 10284 35592 10286 35601
rect 10230 35527 10286 35536
rect 11060 35080 11112 35086
rect 11060 35022 11112 35028
rect 10968 34944 11020 34950
rect 10968 34886 11020 34892
rect 10980 34678 11008 34886
rect 10968 34672 11020 34678
rect 10966 34640 10968 34649
rect 11020 34640 11022 34649
rect 10876 34604 10928 34610
rect 10966 34575 11022 34584
rect 10876 34546 10928 34552
rect 10980 34549 11008 34575
rect 10324 34400 10376 34406
rect 10324 34342 10376 34348
rect 10140 34128 10192 34134
rect 10140 34070 10192 34076
rect 10152 33658 10180 34070
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 10152 33386 10180 33594
rect 10336 33590 10364 34342
rect 10508 33856 10560 33862
rect 10508 33798 10560 33804
rect 10324 33584 10376 33590
rect 10520 33561 10548 33798
rect 10324 33526 10376 33532
rect 10506 33552 10562 33561
rect 10506 33487 10508 33496
rect 10560 33487 10562 33496
rect 10508 33458 10560 33464
rect 10140 33380 10192 33386
rect 10140 33322 10192 33328
rect 10046 32464 10102 32473
rect 10046 32399 10048 32408
rect 10100 32399 10102 32408
rect 10048 32370 10100 32376
rect 9864 32292 9916 32298
rect 9864 32234 9916 32240
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 10046 31920 10102 31929
rect 9956 31884 10008 31890
rect 10046 31855 10102 31864
rect 9956 31826 10008 31832
rect 9496 31680 9548 31686
rect 9496 31622 9548 31628
rect 9508 31278 9536 31622
rect 9588 31340 9640 31346
rect 9588 31282 9640 31288
rect 9496 31272 9548 31278
rect 9496 31214 9548 31220
rect 9600 30258 9628 31282
rect 9968 31210 9996 31826
rect 9956 31204 10008 31210
rect 9956 31146 10008 31152
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9680 30728 9732 30734
rect 9680 30670 9732 30676
rect 9588 30252 9640 30258
rect 9588 30194 9640 30200
rect 9600 29850 9628 30194
rect 9692 30054 9720 30670
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9588 29844 9640 29850
rect 9588 29786 9640 29792
rect 9692 29730 9720 29990
rect 9600 29702 9720 29730
rect 9600 28694 9628 29702
rect 9784 28966 9812 31078
rect 9968 30705 9996 31146
rect 10060 30716 10088 31855
rect 10152 30870 10180 33322
rect 10888 33046 10916 34546
rect 11072 34134 11100 35022
rect 11060 34128 11112 34134
rect 11060 34070 11112 34076
rect 10324 33040 10376 33046
rect 10324 32982 10376 32988
rect 10876 33040 10928 33046
rect 10876 32982 10928 32988
rect 10336 32570 10364 32982
rect 10324 32564 10376 32570
rect 10324 32506 10376 32512
rect 10888 32434 10916 32982
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 10888 32178 10916 32370
rect 10796 32150 10916 32178
rect 10600 31680 10652 31686
rect 10600 31622 10652 31628
rect 10612 31210 10640 31622
rect 10796 31346 10824 32150
rect 11164 31890 11192 36518
rect 11244 36236 11296 36242
rect 11244 36178 11296 36184
rect 11256 35578 11284 36178
rect 11348 35834 11376 39520
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11992 36961 12020 39520
rect 12070 37496 12126 37505
rect 12070 37431 12126 37440
rect 11978 36952 12034 36961
rect 11978 36887 12034 36896
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 12084 35834 12112 37431
rect 12544 36394 12572 39520
rect 12360 36378 12572 36394
rect 12348 36372 12572 36378
rect 12400 36366 12572 36372
rect 12348 36314 12400 36320
rect 11336 35828 11388 35834
rect 11336 35770 11388 35776
rect 12072 35828 12124 35834
rect 12072 35770 12124 35776
rect 11256 35550 11376 35578
rect 11348 35494 11376 35550
rect 11336 35488 11388 35494
rect 11336 35430 11388 35436
rect 11980 35488 12032 35494
rect 11980 35430 12032 35436
rect 12992 35488 13044 35494
rect 12992 35430 13044 35436
rect 11244 35148 11296 35154
rect 11244 35090 11296 35096
rect 11256 34542 11284 35090
rect 11244 34536 11296 34542
rect 11244 34478 11296 34484
rect 11152 31884 11204 31890
rect 11152 31826 11204 31832
rect 10784 31340 10836 31346
rect 10784 31282 10836 31288
rect 10600 31204 10652 31210
rect 10600 31146 10652 31152
rect 10612 30938 10640 31146
rect 10796 30938 10824 31282
rect 10600 30932 10652 30938
rect 10600 30874 10652 30880
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10140 30864 10192 30870
rect 10140 30806 10192 30812
rect 9954 30696 10010 30705
rect 10060 30688 10180 30716
rect 9954 30631 10010 30640
rect 10048 29776 10100 29782
rect 10048 29718 10100 29724
rect 9956 29640 10008 29646
rect 9956 29582 10008 29588
rect 9968 29073 9996 29582
rect 9954 29064 10010 29073
rect 10060 29034 10088 29718
rect 9954 28999 10010 29008
rect 10048 29028 10100 29034
rect 9772 28960 9824 28966
rect 9772 28902 9824 28908
rect 9588 28688 9640 28694
rect 9588 28630 9640 28636
rect 9784 28626 9812 28902
rect 9968 28762 9996 28999
rect 10048 28970 10100 28976
rect 9956 28756 10008 28762
rect 9956 28698 10008 28704
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9784 28218 9812 28562
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9680 28008 9732 28014
rect 8956 27674 8984 27950
rect 9324 27934 9536 27962
rect 9680 27950 9732 27956
rect 9404 27872 9456 27878
rect 9508 27849 9536 27934
rect 9404 27814 9456 27820
rect 9494 27840 9550 27849
rect 9416 27674 9444 27814
rect 9494 27775 9550 27784
rect 8944 27668 8996 27674
rect 8944 27610 8996 27616
rect 9404 27668 9456 27674
rect 9404 27610 9456 27616
rect 9508 27441 9536 27775
rect 9692 27674 9720 27950
rect 9772 27940 9824 27946
rect 9772 27882 9824 27888
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 9494 27432 9550 27441
rect 9494 27367 9550 27376
rect 9496 27328 9548 27334
rect 9494 27296 9496 27305
rect 9548 27296 9550 27305
rect 8956 27228 9252 27248
rect 9494 27231 9550 27240
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9692 26994 9720 27610
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 8758 26480 8814 26489
rect 8864 26450 8892 26726
rect 8758 26415 8814 26424
rect 8852 26444 8904 26450
rect 8852 26386 8904 26392
rect 8760 26376 8812 26382
rect 8760 26318 8812 26324
rect 8772 25498 8800 26318
rect 8864 25702 8892 26386
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 9600 25906 9628 26182
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 9600 25786 9628 25842
rect 9404 25764 9456 25770
rect 9600 25758 9720 25786
rect 9404 25706 9456 25712
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8772 24818 8800 25434
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 8576 24608 8628 24614
rect 8574 24576 8576 24585
rect 8628 24576 8630 24585
rect 8574 24511 8630 24520
rect 8404 24126 8524 24154
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8404 23202 8432 24126
rect 8588 23662 8616 24142
rect 8864 24138 8892 25638
rect 9416 25498 9444 25706
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 8852 24132 8904 24138
rect 8852 24074 8904 24080
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9324 23798 9352 24006
rect 8760 23792 8812 23798
rect 8758 23760 8760 23769
rect 9312 23792 9364 23798
rect 8812 23760 8814 23769
rect 9312 23734 9364 23740
rect 8758 23695 8814 23704
rect 8576 23656 8628 23662
rect 8574 23624 8576 23633
rect 8628 23624 8630 23633
rect 8574 23559 8630 23568
rect 9404 23588 9456 23594
rect 9404 23530 9456 23536
rect 8312 23174 8432 23202
rect 8484 23180 8536 23186
rect 8312 22098 8340 23174
rect 8484 23122 8536 23128
rect 8496 22710 8524 23122
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8484 22704 8536 22710
rect 8404 22664 8484 22692
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8128 21146 8156 21966
rect 8404 21486 8432 22664
rect 8484 22646 8536 22652
rect 8772 22642 8800 23054
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8772 22234 8800 22578
rect 8760 22228 8812 22234
rect 8760 22170 8812 22176
rect 8850 22128 8906 22137
rect 8576 22092 8628 22098
rect 8850 22063 8906 22072
rect 8576 22034 8628 22040
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8220 20584 8248 20946
rect 8404 20942 8432 21422
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8300 20596 8352 20602
rect 8128 20556 8300 20584
rect 8022 19136 8078 19145
rect 8022 19071 8078 19080
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 8036 18222 8064 19071
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 8128 17898 8156 20556
rect 8300 20538 8352 20544
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 8220 18834 8248 20266
rect 8404 19922 8432 20878
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8496 19446 8524 19722
rect 8484 19440 8536 19446
rect 8484 19382 8536 19388
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7944 17870 8156 17898
rect 8220 17882 8248 18770
rect 8312 18737 8340 19110
rect 8298 18728 8354 18737
rect 8298 18663 8354 18672
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8404 18222 8432 18634
rect 8392 18216 8444 18222
rect 8588 18170 8616 22034
rect 8760 21684 8812 21690
rect 8760 21626 8812 21632
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8680 21146 8708 21354
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8680 20466 8708 21082
rect 8772 20602 8800 21626
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8666 20224 8722 20233
rect 8666 20159 8722 20168
rect 8392 18158 8444 18164
rect 8496 18142 8616 18170
rect 8208 17876 8260 17882
rect 7838 17368 7894 17377
rect 7838 17303 7894 17312
rect 7944 17218 7972 17870
rect 8208 17818 8260 17824
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7852 17190 7972 17218
rect 7852 16046 7880 17190
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7944 16726 7972 17070
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 8036 16658 8064 17614
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7852 15706 7880 15982
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7852 15337 7880 15642
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7838 15328 7894 15337
rect 7838 15263 7894 15272
rect 8036 15162 8064 15506
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14550 7788 14758
rect 7392 14470 7512 14498
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 8022 14512 8078 14521
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7300 11898 7328 12310
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7194 9208 7250 9217
rect 7194 9143 7250 9152
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 7993 7052 8978
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8498 7144 8910
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7010 7984 7066 7993
rect 7010 7919 7066 7928
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6932 6866 6960 7210
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 7024 6798 7052 7346
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6186 7052 6598
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6932 5914 6960 6122
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 5846 7052 6122
rect 7116 5846 7144 7822
rect 7208 7449 7236 9143
rect 7392 9081 7420 14470
rect 8128 14482 8156 17682
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8220 16726 8248 17138
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8312 15706 8340 16594
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8404 15026 8432 15914
rect 8496 15722 8524 18142
rect 8574 18048 8630 18057
rect 8574 17983 8630 17992
rect 8588 17882 8616 17983
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8588 16250 8616 16662
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8680 16153 8708 20159
rect 8758 19816 8814 19825
rect 8758 19751 8814 19760
rect 8772 19718 8800 19751
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8772 19310 8800 19654
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8772 18465 8800 18838
rect 8758 18456 8814 18465
rect 8758 18391 8760 18400
rect 8812 18391 8814 18400
rect 8760 18362 8812 18368
rect 8864 16969 8892 22063
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9324 20330 9352 20538
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9324 18426 9352 20266
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9416 18306 9444 23530
rect 9508 22438 9536 24550
rect 9692 24410 9720 25758
rect 9784 25702 9812 27882
rect 10060 27606 10088 28970
rect 10152 27878 10180 30688
rect 10692 29776 10744 29782
rect 10692 29718 10744 29724
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10140 27872 10192 27878
rect 10140 27814 10192 27820
rect 10048 27600 10100 27606
rect 10048 27542 10100 27548
rect 10060 27130 10088 27542
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 10152 26586 10180 27406
rect 10244 27305 10272 28494
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 10230 27296 10286 27305
rect 10230 27231 10286 27240
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 9772 25696 9824 25702
rect 9772 25638 9824 25644
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 10060 25430 10088 25638
rect 10048 25424 10100 25430
rect 10048 25366 10100 25372
rect 10060 24682 10088 25366
rect 10048 24676 10100 24682
rect 10048 24618 10100 24624
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 9586 24032 9642 24041
rect 9586 23967 9642 23976
rect 9600 23866 9628 23967
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9692 23526 9720 24210
rect 10152 24138 10180 24210
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 10152 23866 10180 24074
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 9680 23520 9732 23526
rect 9678 23488 9680 23497
rect 9732 23488 9734 23497
rect 9678 23423 9734 23432
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9508 22234 9536 22374
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9692 22166 9720 22510
rect 9680 22160 9732 22166
rect 9680 22102 9732 22108
rect 9680 22024 9732 22030
rect 9678 21992 9680 22001
rect 9732 21992 9734 22001
rect 9678 21927 9734 21936
rect 9692 21622 9720 21927
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9600 20806 9628 21422
rect 9956 21412 10008 21418
rect 9956 21354 10008 21360
rect 9968 21078 9996 21354
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 10230 20904 10286 20913
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 19242 9628 20742
rect 9692 20398 9720 20878
rect 10230 20839 10286 20848
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9692 20058 9720 20334
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 10244 19990 10272 20839
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10060 19310 10088 19858
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9784 19174 9812 19246
rect 9772 19168 9824 19174
rect 9770 19136 9772 19145
rect 9824 19136 9826 19145
rect 9770 19071 9826 19080
rect 10244 18970 10272 19926
rect 10336 19394 10364 27814
rect 10704 27470 10732 29718
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 11058 29608 11114 29617
rect 10796 28490 10824 29582
rect 11058 29543 11114 29552
rect 10968 29504 11020 29510
rect 10968 29446 11020 29452
rect 10980 29238 11008 29446
rect 11072 29306 11100 29543
rect 11060 29300 11112 29306
rect 11060 29242 11112 29248
rect 10968 29232 11020 29238
rect 10968 29174 11020 29180
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 10888 28626 10916 29106
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10692 27464 10744 27470
rect 10692 27406 10744 27412
rect 10796 26874 10824 28426
rect 10888 27606 10916 28562
rect 10980 28150 11008 29174
rect 11060 29028 11112 29034
rect 11060 28970 11112 28976
rect 10968 28144 11020 28150
rect 10968 28086 11020 28092
rect 10876 27600 10928 27606
rect 10876 27542 10928 27548
rect 10888 26994 10916 27542
rect 11072 27538 11100 28970
rect 11256 28762 11284 34478
rect 11244 28756 11296 28762
rect 11244 28698 11296 28704
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 11164 28218 11192 28630
rect 11152 28212 11204 28218
rect 11152 28154 11204 28160
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 10876 26988 10928 26994
rect 11256 26976 11284 28698
rect 11348 27334 11376 35430
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11520 34128 11572 34134
rect 11520 34070 11572 34076
rect 11704 34128 11756 34134
rect 11704 34070 11756 34076
rect 11428 33312 11480 33318
rect 11428 33254 11480 33260
rect 11440 32570 11468 33254
rect 11532 33114 11560 34070
rect 11716 33658 11744 34070
rect 11992 33998 12020 35430
rect 12070 35320 12126 35329
rect 12070 35255 12072 35264
rect 12124 35255 12126 35264
rect 12072 35226 12124 35232
rect 12070 35184 12126 35193
rect 12070 35119 12126 35128
rect 12440 35148 12492 35154
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 11704 33652 11756 33658
rect 11704 33594 11756 33600
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11520 33108 11572 33114
rect 11520 33050 11572 33056
rect 11532 32910 11560 33050
rect 11888 33040 11940 33046
rect 11888 32982 11940 32988
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 11900 32570 11928 32982
rect 11428 32564 11480 32570
rect 11428 32506 11480 32512
rect 11888 32564 11940 32570
rect 11888 32506 11940 32512
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11992 31346 12020 33934
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11612 30864 11664 30870
rect 11612 30806 11664 30812
rect 11520 30728 11572 30734
rect 11520 30670 11572 30676
rect 11532 30394 11560 30670
rect 11520 30388 11572 30394
rect 11520 30330 11572 30336
rect 11532 29850 11560 30330
rect 11624 30326 11652 30806
rect 11992 30734 12020 31282
rect 11980 30728 12032 30734
rect 11980 30670 12032 30676
rect 11612 30320 11664 30326
rect 11612 30262 11664 30268
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11520 29844 11572 29850
rect 11520 29786 11572 29792
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11978 28520 12034 28529
rect 11978 28455 12034 28464
rect 11992 28082 12020 28455
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 11428 27872 11480 27878
rect 11426 27840 11428 27849
rect 11480 27840 11482 27849
rect 11426 27775 11482 27784
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11612 27600 11664 27606
rect 11612 27542 11664 27548
rect 11520 27396 11572 27402
rect 11520 27338 11572 27344
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 11256 26948 11376 26976
rect 10876 26930 10928 26936
rect 10600 26852 10652 26858
rect 10796 26846 10916 26874
rect 10600 26794 10652 26800
rect 10612 26586 10640 26794
rect 10600 26580 10652 26586
rect 10600 26522 10652 26528
rect 10612 26042 10640 26522
rect 10692 26512 10744 26518
rect 10692 26454 10744 26460
rect 10704 26042 10732 26454
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10704 25498 10732 25978
rect 10796 25702 10824 26318
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10796 25498 10824 25638
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10888 25430 10916 26846
rect 11244 26852 11296 26858
rect 11244 26794 11296 26800
rect 11256 26518 11284 26794
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 11256 25838 11284 26454
rect 11244 25832 11296 25838
rect 11244 25774 11296 25780
rect 11256 25430 11284 25774
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 11244 25424 11296 25430
rect 11244 25366 11296 25372
rect 10888 24818 10916 25366
rect 11256 24818 11284 25366
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 11242 24576 11298 24585
rect 11242 24511 11298 24520
rect 11256 24342 11284 24511
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 10520 23730 10548 24074
rect 10600 24064 10652 24070
rect 11072 24041 11100 24210
rect 10600 24006 10652 24012
rect 11058 24032 11114 24041
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10612 23610 10640 24006
rect 11058 23967 11114 23976
rect 11072 23866 11100 23967
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 10520 23594 10640 23610
rect 10508 23588 10640 23594
rect 10560 23582 10640 23588
rect 10508 23530 10560 23536
rect 10520 23254 10548 23530
rect 10508 23248 10560 23254
rect 10508 23190 10560 23196
rect 10416 23112 10468 23118
rect 10414 23080 10416 23089
rect 10468 23080 10470 23089
rect 10414 23015 10470 23024
rect 10520 22574 10548 23190
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10888 22234 10916 22442
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10980 21962 11008 22578
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10336 19366 10456 19394
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9324 18278 9444 18306
rect 9324 17785 9352 18278
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 17882 9444 18158
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9310 17776 9366 17785
rect 9600 17762 9628 18702
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10060 17814 10088 18090
rect 10048 17808 10100 17814
rect 9600 17746 9720 17762
rect 10048 17750 10100 17756
rect 9600 17740 9732 17746
rect 9600 17734 9680 17740
rect 9310 17711 9366 17720
rect 9680 17682 9732 17688
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 8850 16960 8906 16969
rect 8850 16895 8906 16904
rect 9140 16794 9168 17070
rect 9692 16794 9720 17682
rect 10060 17338 10088 17750
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9770 16824 9826 16833
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9680 16788 9732 16794
rect 9770 16759 9826 16768
rect 9680 16730 9732 16736
rect 8850 16688 8906 16697
rect 8850 16623 8906 16632
rect 9588 16652 9640 16658
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8666 16144 8722 16153
rect 8666 16079 8722 16088
rect 8666 16008 8722 16017
rect 8666 15943 8722 15952
rect 8496 15694 8616 15722
rect 8680 15706 8708 15943
rect 8482 15600 8538 15609
rect 8482 15535 8484 15544
rect 8536 15535 8538 15544
rect 8484 15506 8536 15512
rect 8496 15162 8524 15506
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8022 14447 8078 14456
rect 8116 14476 8168 14482
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 13326 7604 13806
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7484 9654 7512 10134
rect 7576 10062 7604 13262
rect 7668 12986 7696 13398
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7668 12714 7696 12922
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7668 12442 7696 12650
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7378 9072 7434 9081
rect 7378 9007 7434 9016
rect 7194 7440 7250 7449
rect 7194 7375 7250 7384
rect 7288 7200 7340 7206
rect 7208 7148 7288 7154
rect 7208 7142 7340 7148
rect 7208 7126 7328 7142
rect 7208 6322 7236 7126
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5166 6868 5646
rect 7010 5400 7066 5409
rect 7010 5335 7066 5344
rect 6828 5160 6880 5166
rect 6276 5102 6328 5108
rect 6734 5128 6790 5137
rect 6828 5102 6880 5108
rect 6734 5063 6790 5072
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4185 6132 4966
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6748 4842 6776 5063
rect 6748 4814 6960 4842
rect 6932 4758 6960 4814
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6196 4486 6224 4694
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6090 4176 6146 4185
rect 6090 4111 6146 4120
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3505 6132 3878
rect 6090 3496 6146 3505
rect 6196 3466 6224 4422
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6090 3431 6146 3440
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6288 3194 6316 3606
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6656 3058 6684 4082
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6748 2650 6776 3878
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6840 3058 6868 3538
rect 6932 3369 6960 3946
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 5920 2417 5948 2450
rect 5906 2408 5962 2417
rect 5906 2343 5962 2352
rect 7024 2258 7052 5335
rect 7116 5234 7144 5782
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7116 4554 7144 5170
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 2650 7144 4490
rect 7208 4146 7236 6258
rect 7668 5409 7696 12106
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7760 11286 7788 11630
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7852 11098 7880 12174
rect 7944 11830 7972 12378
rect 8036 12170 8064 14447
rect 8116 14418 8168 14424
rect 8128 14074 8156 14418
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8128 13870 8156 14010
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8312 12866 8340 14350
rect 8390 13424 8446 13433
rect 8390 13359 8446 13368
rect 8220 12850 8340 12866
rect 8208 12844 8340 12850
rect 8260 12838 8340 12844
rect 8208 12786 8260 12792
rect 8404 12753 8432 13359
rect 8390 12744 8446 12753
rect 8390 12679 8446 12688
rect 8208 12640 8260 12646
rect 8128 12600 8208 12628
rect 8128 12374 8156 12600
rect 8208 12582 8260 12588
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 11626 7972 11766
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7944 11286 7972 11562
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7760 11082 7880 11098
rect 7748 11076 7880 11082
rect 7800 11070 7880 11076
rect 7748 11018 7800 11024
rect 7760 10713 7788 11018
rect 7944 10810 7972 11222
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7746 10704 7802 10713
rect 7746 10639 7802 10648
rect 7944 9722 7972 10746
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10198 8064 10610
rect 8312 10266 8340 11086
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7944 9110 7972 9658
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7760 8566 7788 9046
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7760 7274 7788 8502
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7760 7002 7788 7210
rect 7852 7206 7880 7822
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7760 6458 7788 6938
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7654 5400 7710 5409
rect 7654 5335 7710 5344
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4146 7788 6394
rect 7944 5302 7972 8434
rect 8036 5846 8064 8774
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8128 8106 8156 8298
rect 8128 8078 8248 8106
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 7546 8156 7958
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8220 6474 8248 8078
rect 8220 6458 8340 6474
rect 8220 6452 8352 6458
rect 8220 6446 8300 6452
rect 8300 6394 8352 6400
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 8036 5370 8064 5782
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7932 5296 7984 5302
rect 8404 5250 8432 12679
rect 7932 5238 7984 5244
rect 7944 5166 7972 5238
rect 8312 5222 8432 5250
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7944 4282 7972 5102
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4593 8064 4626
rect 8022 4584 8078 4593
rect 8022 4519 8078 4528
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7196 4140 7248 4146
rect 7748 4140 7800 4146
rect 7196 4082 7248 4088
rect 7668 4100 7748 4128
rect 7286 3768 7342 3777
rect 7286 3703 7342 3712
rect 7300 2854 7328 3703
rect 7668 3670 7696 4100
rect 7748 4082 7800 4088
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7472 3392 7524 3398
rect 7470 3360 7472 3369
rect 7524 3360 7526 3369
rect 7470 3295 7526 3304
rect 7760 3194 7788 3878
rect 8024 3664 8076 3670
rect 7838 3632 7894 3641
rect 8024 3606 8076 3612
rect 7838 3567 7840 3576
rect 7892 3567 7894 3576
rect 7840 3538 7892 3544
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7852 2650 7880 3538
rect 8036 3194 8064 3606
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8312 2961 8340 5222
rect 8496 5166 8524 14554
rect 8588 13433 8616 15694
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8680 14618 8708 15642
rect 8772 15162 8800 16186
rect 8864 16114 8892 16623
rect 9588 16594 9640 16600
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8864 15706 8892 16050
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8772 14890 8800 15098
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8956 14618 8984 14962
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8574 13424 8630 13433
rect 8574 13359 8630 13368
rect 8680 13326 8708 13670
rect 8772 13530 8800 13806
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8772 13410 8800 13466
rect 8772 13382 8892 13410
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12374 8616 13126
rect 8680 12986 8708 13262
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8574 12200 8630 12209
rect 8574 12135 8630 12144
rect 8588 9518 8616 12135
rect 8772 11898 8800 12650
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8772 11234 8800 11834
rect 8680 11206 8800 11234
rect 8680 10538 8708 11206
rect 8864 11121 8892 13382
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9600 12866 9628 16594
rect 9784 15570 9812 16759
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9784 14618 9812 15506
rect 9876 14929 9904 17070
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16794 10088 16934
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9968 15638 9996 15914
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9968 15162 9996 15574
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9862 14920 9918 14929
rect 9862 14855 9918 14864
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9876 14550 9904 14758
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12986 9812 13262
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9600 12838 9720 12866
rect 9876 12850 9904 13398
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9140 11354 9168 11698
rect 9416 11354 9444 12174
rect 9508 11898 9536 12310
rect 9600 12102 9628 12650
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9600 11370 9628 12038
rect 9692 11558 9720 12838
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9968 12442 9996 15098
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10336 13802 10364 14010
rect 10232 13796 10284 13802
rect 10232 13738 10284 13744
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10244 13530 10272 13738
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 9956 12436 10008 12442
rect 10008 12396 10088 12424
rect 9956 12378 10008 12384
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9404 11348 9456 11354
rect 9600 11342 9812 11370
rect 9404 11290 9456 11296
rect 9140 11234 9168 11290
rect 9496 11280 9548 11286
rect 9140 11206 9352 11234
rect 9496 11222 9548 11228
rect 9586 11248 9642 11257
rect 8850 11112 8906 11121
rect 8850 11047 8906 11056
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10810 8800 10950
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 9324 10742 9352 11206
rect 9402 10840 9458 10849
rect 9508 10810 9536 11222
rect 9586 11183 9642 11192
rect 9402 10775 9458 10784
rect 9496 10804 9548 10810
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9416 10674 9444 10775
rect 9496 10746 9548 10752
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8772 10266 8800 10610
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 9600 9602 9628 11183
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9508 9574 9628 9602
rect 9692 9586 9720 9998
rect 9680 9580 9732 9586
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8588 9178 8616 9454
rect 8758 9208 8814 9217
rect 8576 9172 8628 9178
rect 8758 9143 8760 9152
rect 8576 9114 8628 9120
rect 8812 9143 8814 9152
rect 8760 9114 8812 9120
rect 8772 8514 8800 9114
rect 8680 8486 8800 8514
rect 8864 8498 8892 9454
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8852 8492 8904 8498
rect 8680 8430 8708 8486
rect 8852 8434 8904 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7290 8800 7822
rect 8864 7410 8892 8298
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 8850 7304 8906 7313
rect 8772 7262 8850 7290
rect 8850 7239 8906 7248
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6186 8800 6598
rect 8864 6338 8892 7239
rect 9232 7002 9260 7346
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8864 6322 8984 6338
rect 8864 6316 8996 6322
rect 8864 6310 8944 6316
rect 8944 6258 8996 6264
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 5914 8800 6122
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8956 5846 8984 6258
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8404 4078 8432 5034
rect 8496 4321 8524 5102
rect 8588 4690 8616 5238
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9232 4826 9260 5102
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8482 4312 8538 4321
rect 8482 4247 8538 4256
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8404 3670 8432 4014
rect 8666 3904 8722 3913
rect 8666 3839 8722 3848
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8680 3233 8708 3839
rect 8772 3738 8800 4558
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9508 4026 9536 9574
rect 9680 9522 9732 9528
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9600 8378 9628 9386
rect 9784 9178 9812 11342
rect 9862 11112 9918 11121
rect 9862 11047 9918 11056
rect 9876 9518 9904 11047
rect 10060 10198 10088 12396
rect 10244 12170 10272 12650
rect 10428 12594 10456 19366
rect 10690 18864 10746 18873
rect 10690 18799 10692 18808
rect 10744 18799 10746 18808
rect 10692 18770 10744 18776
rect 10704 18426 10732 18770
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10612 16250 10640 16526
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10704 15994 10732 16662
rect 10612 15966 10732 15994
rect 10612 15910 10640 15966
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10612 15162 10640 15302
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10612 14890 10640 15098
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10612 14074 10640 14826
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10336 12566 10456 12594
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10244 11150 10272 12106
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10152 10198 10180 10474
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10336 9738 10364 12566
rect 10520 12442 10548 13262
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10520 11762 10548 12378
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10428 11286 10456 11562
rect 10796 11558 10824 21422
rect 10968 20800 11020 20806
rect 10874 20768 10930 20777
rect 10968 20742 11020 20748
rect 10874 20703 10930 20712
rect 10888 19854 10916 20703
rect 10980 20534 11008 20742
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10980 20058 11008 20266
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10980 19514 11008 19994
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11072 19009 11100 22918
rect 11164 22642 11192 23054
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11164 20942 11192 22578
rect 11348 21486 11376 26948
rect 11428 26920 11480 26926
rect 11426 26888 11428 26897
rect 11480 26888 11482 26897
rect 11426 26823 11482 26832
rect 11532 26586 11560 27338
rect 11624 27130 11652 27542
rect 11978 27432 12034 27441
rect 11978 27367 12034 27376
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11992 26042 12020 27367
rect 12084 26450 12112 35119
rect 12440 35090 12492 35096
rect 12452 34921 12480 35090
rect 12438 34912 12494 34921
rect 12438 34847 12494 34856
rect 12348 34604 12400 34610
rect 12348 34546 12400 34552
rect 12176 33522 12296 33538
rect 12176 33516 12308 33522
rect 12176 33510 12256 33516
rect 12176 32910 12204 33510
rect 12256 33458 12308 33464
rect 12256 33380 12308 33386
rect 12256 33322 12308 33328
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 12268 32026 12296 33322
rect 12360 33114 12388 34546
rect 12452 34542 12480 34847
rect 12622 34640 12678 34649
rect 12622 34575 12678 34584
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 12544 33386 12572 33798
rect 12532 33380 12584 33386
rect 12532 33322 12584 33328
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 12360 32570 12388 33050
rect 12636 32570 12664 34575
rect 12900 32768 12952 32774
rect 12900 32710 12952 32716
rect 12348 32564 12400 32570
rect 12348 32506 12400 32512
rect 12624 32564 12676 32570
rect 12624 32506 12676 32512
rect 12912 32473 12940 32710
rect 12898 32464 12954 32473
rect 12898 32399 12954 32408
rect 12440 32360 12492 32366
rect 12440 32302 12492 32308
rect 12256 32020 12308 32026
rect 12256 31962 12308 31968
rect 12452 31929 12480 32302
rect 12438 31920 12494 31929
rect 12164 31884 12216 31890
rect 12438 31855 12494 31864
rect 12164 31826 12216 31832
rect 12176 31142 12204 31826
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 12176 27418 12204 31078
rect 12348 29708 12400 29714
rect 12348 29650 12400 29656
rect 12360 29306 12388 29650
rect 13004 29306 13032 35430
rect 13188 35329 13216 39520
rect 13728 35828 13780 35834
rect 13832 35816 13860 39520
rect 14384 37210 14412 39520
rect 13780 35788 13860 35816
rect 14200 37182 14412 37210
rect 13728 35770 13780 35776
rect 13174 35320 13230 35329
rect 14200 35290 14228 37182
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 13174 35255 13230 35264
rect 14188 35284 14240 35290
rect 14188 35226 14240 35232
rect 13634 35048 13690 35057
rect 13634 34983 13690 34992
rect 13648 34746 13676 34983
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 13912 34536 13964 34542
rect 13912 34478 13964 34484
rect 13542 34232 13598 34241
rect 13542 34167 13544 34176
rect 13596 34167 13598 34176
rect 13544 34138 13596 34144
rect 13544 34060 13596 34066
rect 13544 34002 13596 34008
rect 13556 33318 13584 34002
rect 13544 33312 13596 33318
rect 13544 33254 13596 33260
rect 13556 32978 13584 33254
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13556 32230 13584 32914
rect 13544 32224 13596 32230
rect 13544 32166 13596 32172
rect 12348 29300 12400 29306
rect 12348 29242 12400 29248
rect 12992 29300 13044 29306
rect 12992 29242 13044 29248
rect 13450 29200 13506 29209
rect 13450 29135 13506 29144
rect 13464 29102 13492 29135
rect 12440 29096 12492 29102
rect 13452 29096 13504 29102
rect 12440 29038 12492 29044
rect 12990 29064 13046 29073
rect 12348 28484 12400 28490
rect 12348 28426 12400 28432
rect 12360 27606 12388 28426
rect 12348 27600 12400 27606
rect 12348 27542 12400 27548
rect 12452 27554 12480 29038
rect 13452 29038 13504 29044
rect 12990 28999 12992 29008
rect 13044 28999 13046 29008
rect 12992 28970 13044 28976
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12544 27674 12572 28494
rect 13176 28144 13228 28150
rect 13176 28086 13228 28092
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12532 27668 12584 27674
rect 12532 27610 12584 27616
rect 12452 27526 12572 27554
rect 12176 27390 12296 27418
rect 12164 27328 12216 27334
rect 12164 27270 12216 27276
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12084 26042 12112 26386
rect 11980 26036 12032 26042
rect 11980 25978 12032 25984
rect 12072 26036 12124 26042
rect 12072 25978 12124 25984
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11532 22137 11560 25842
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 12070 24440 12126 24449
rect 12070 24375 12126 24384
rect 11978 23760 12034 23769
rect 11978 23695 12034 23704
rect 11992 23662 12020 23695
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11980 23248 12032 23254
rect 11978 23216 11980 23225
rect 12032 23216 12034 23225
rect 12084 23186 12112 24375
rect 11978 23151 12034 23160
rect 12072 23180 12124 23186
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11992 22166 12020 23151
rect 12072 23122 12124 23128
rect 12084 22778 12112 23122
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12176 22574 12204 27270
rect 12164 22568 12216 22574
rect 12084 22528 12164 22556
rect 11612 22160 11664 22166
rect 11518 22128 11574 22137
rect 11612 22102 11664 22108
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11518 22063 11574 22072
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11532 21078 11560 21830
rect 11624 21690 11652 22102
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11992 21690 12020 21966
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11164 20466 11192 20878
rect 11532 20602 11560 21014
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11992 20058 12020 21626
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12084 19990 12112 22528
rect 12164 22510 12216 22516
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12176 21554 12204 21966
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12176 20942 12204 21490
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11058 19000 11114 19009
rect 11058 18935 11114 18944
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 18329 10916 18566
rect 10874 18320 10930 18329
rect 10874 18255 10930 18264
rect 11060 18216 11112 18222
rect 11152 18216 11204 18222
rect 11060 18158 11112 18164
rect 11150 18184 11152 18193
rect 11204 18184 11206 18193
rect 11072 17882 11100 18158
rect 11150 18119 11206 18128
rect 11152 18080 11204 18086
rect 11150 18048 11152 18057
rect 11204 18048 11206 18057
rect 11440 18034 11468 19926
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11150 17983 11206 17992
rect 11348 18006 11468 18034
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11348 17338 11376 18006
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11348 17134 11376 17274
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10874 16144 10930 16153
rect 10874 16079 10930 16088
rect 10888 15910 10916 16079
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 13297 10916 15846
rect 11072 15638 11100 16934
rect 11440 16794 11468 17818
rect 11532 17814 11560 18702
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11532 17338 11560 17750
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17338 12204 17478
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12176 17066 12204 17274
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 11164 15450 11192 16458
rect 12176 16250 12204 16662
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11072 15422 11192 15450
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10980 15026 11008 15302
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 11072 14890 11100 15422
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 11072 14482 11100 14826
rect 11532 14618 11560 15574
rect 11716 15162 11744 15574
rect 12268 15570 12296 27390
rect 12438 27296 12494 27305
rect 12438 27231 12494 27240
rect 12452 27130 12480 27231
rect 12440 27124 12492 27130
rect 12440 27066 12492 27072
rect 12544 24857 12572 27526
rect 12530 24848 12586 24857
rect 12530 24783 12586 24792
rect 12728 24449 12756 27814
rect 13188 27674 13216 28086
rect 13176 27668 13228 27674
rect 13176 27610 13228 27616
rect 13082 27568 13138 27577
rect 13082 27503 13084 27512
rect 13136 27503 13138 27512
rect 13084 27474 13136 27480
rect 13096 27130 13124 27474
rect 13084 27124 13136 27130
rect 13136 27084 13216 27112
rect 13084 27066 13136 27072
rect 12714 24440 12770 24449
rect 12714 24375 12770 24384
rect 12530 24168 12586 24177
rect 12348 24132 12400 24138
rect 12400 24092 12480 24120
rect 12530 24103 12586 24112
rect 12348 24074 12400 24080
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12360 21978 12388 23530
rect 12452 22778 12480 24092
rect 12544 23662 12572 24103
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12728 23866 12756 24006
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12624 23792 12676 23798
rect 12622 23760 12624 23769
rect 12676 23760 12678 23769
rect 12622 23695 12678 23704
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12544 23322 12572 23598
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12898 23080 12954 23089
rect 12898 23015 12954 23024
rect 12912 22778 12940 23015
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 13096 22545 13124 23462
rect 13188 22574 13216 27084
rect 13176 22568 13228 22574
rect 13082 22536 13138 22545
rect 13176 22510 13228 22516
rect 13082 22471 13138 22480
rect 13188 22420 13216 22510
rect 12912 22392 13216 22420
rect 12360 21950 12480 21978
rect 12452 21944 12480 21950
rect 12532 21956 12584 21962
rect 12452 21916 12532 21944
rect 12532 21898 12584 21904
rect 12348 21888 12400 21894
rect 12400 21836 12480 21842
rect 12348 21830 12480 21836
rect 12360 21814 12480 21830
rect 12452 20602 12480 21814
rect 12544 21418 12572 21898
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12624 21412 12676 21418
rect 12624 21354 12676 21360
rect 12544 20942 12572 21354
rect 12636 21146 12664 21354
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12544 20777 12572 20878
rect 12530 20768 12586 20777
rect 12530 20703 12586 20712
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12532 20392 12584 20398
rect 12530 20360 12532 20369
rect 12584 20360 12586 20369
rect 12530 20295 12586 20304
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17202 12572 17478
rect 12714 17232 12770 17241
rect 12532 17196 12584 17202
rect 12820 17202 12848 17614
rect 12714 17167 12770 17176
rect 12808 17196 12860 17202
rect 12532 17138 12584 17144
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 15314 12388 15438
rect 12544 15314 12572 17138
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12636 16250 12664 16526
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12728 16114 12756 17167
rect 12808 17138 12860 17144
rect 12820 16726 12848 17138
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12820 16046 12848 16662
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12360 15286 12572 15314
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11164 14074 11192 14486
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11624 14074 11652 14350
rect 11992 14074 12020 14758
rect 12452 14550 12480 15286
rect 12714 15056 12770 15065
rect 12714 14991 12770 15000
rect 12728 14958 12756 14991
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12452 13938 12480 14486
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11150 13424 11206 13433
rect 11150 13359 11152 13368
rect 11204 13359 11206 13368
rect 11152 13330 11204 13336
rect 10874 13288 10930 13297
rect 10874 13223 10930 13232
rect 11164 12986 11192 13330
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 11072 11762 11100 12922
rect 11152 12776 11204 12782
rect 11150 12744 11152 12753
rect 11204 12744 11206 12753
rect 11150 12679 11206 12688
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11348 12238 11376 12582
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 12070 12472 12126 12481
rect 12070 12407 12126 12416
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11898 11376 12174
rect 11440 11898 11468 12310
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11242 11792 11298 11801
rect 11060 11756 11112 11762
rect 11242 11727 11298 11736
rect 11060 11698 11112 11704
rect 11256 11694 11284 11727
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10428 10674 10456 11222
rect 10968 11144 11020 11150
rect 11020 11092 11192 11098
rect 10968 11086 11192 11092
rect 10980 11070 11192 11086
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10713 11100 10950
rect 11164 10810 11192 11070
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11058 10704 11114 10713
rect 10416 10668 10468 10674
rect 11058 10639 11114 10648
rect 10416 10610 10468 10616
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10266 10640 10406
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10042 9716 10094 9722
rect 10244 9710 10364 9738
rect 10428 9722 10456 10066
rect 10416 9716 10468 9722
rect 10244 9704 10272 9710
rect 10042 9658 10094 9664
rect 10152 9676 10272 9704
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9600 8350 9720 8378
rect 9968 8362 9996 8978
rect 9692 7954 9720 8350
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7546 9720 7890
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9876 6866 9904 8230
rect 10060 8022 10088 9658
rect 10152 9042 10180 9676
rect 10416 9658 10468 9664
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 9110 10456 9454
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10690 9072 10746 9081
rect 10140 9036 10192 9042
rect 10690 9007 10692 9016
rect 10140 8978 10192 8984
rect 10744 9007 10746 9016
rect 10692 8978 10744 8984
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10244 8430 10272 8842
rect 10704 8634 10732 8978
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 7478 10088 7958
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10060 6934 10088 7414
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 7002 10180 7142
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 5914 9904 6802
rect 10060 6458 10088 6870
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10428 6186 10456 6938
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10612 5846 10640 7686
rect 11072 6338 11100 7822
rect 11152 7336 11204 7342
rect 11150 7304 11152 7313
rect 11204 7304 11206 7313
rect 11150 7239 11206 7248
rect 11256 6474 11284 11494
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 12084 11354 12112 12407
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12452 10849 12480 11494
rect 12544 11218 12572 12922
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12438 10840 12494 10849
rect 12544 10810 12572 11154
rect 12438 10775 12494 10784
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11704 7472 11756 7478
rect 11702 7440 11704 7449
rect 11756 7440 11758 7449
rect 11702 7375 11758 7384
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 10980 6322 11100 6338
rect 10968 6316 11100 6322
rect 11020 6310 11100 6316
rect 11164 6446 11284 6474
rect 11348 6458 11376 6802
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11532 6458 11560 6734
rect 11336 6452 11388 6458
rect 10968 6258 11020 6264
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5234 10180 5646
rect 10612 5370 10640 5782
rect 10980 5778 11008 6122
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9678 4584 9734 4593
rect 9678 4519 9734 4528
rect 9692 4146 9720 4519
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9508 3998 9628 4026
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8666 3224 8722 3233
rect 8666 3159 8722 3168
rect 8772 3058 8800 3674
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 8312 2553 8340 2887
rect 9508 2650 9536 3878
rect 9600 3777 9628 3998
rect 9586 3768 9642 3777
rect 9586 3703 9642 3712
rect 9784 3641 9812 5170
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9864 3664 9916 3670
rect 9770 3632 9826 3641
rect 9864 3606 9916 3612
rect 9770 3567 9826 3576
rect 9876 3194 9904 3606
rect 9968 3534 9996 4966
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10060 3942 10088 4694
rect 10152 4622 10180 5170
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10230 4176 10286 4185
rect 10230 4111 10232 4120
rect 10284 4111 10286 4120
rect 10232 4082 10284 4088
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10060 3466 10088 3878
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10060 2922 10088 3402
rect 10428 3058 10456 3674
rect 10520 3398 10548 4558
rect 10784 4480 10836 4486
rect 10782 4448 10784 4457
rect 10836 4448 10838 4457
rect 10782 4383 10838 4392
rect 10980 4146 11008 5510
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10704 3602 10732 3878
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10980 3466 11008 4082
rect 11164 4049 11192 6446
rect 11336 6394 11388 6400
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11532 5574 11560 6394
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11992 5778 12020 6734
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11992 5370 12020 5714
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11244 5296 11296 5302
rect 11242 5264 11244 5273
rect 11296 5264 11298 5273
rect 11242 5199 11298 5208
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11256 4690 11284 5102
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 4282 11284 4626
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11150 4040 11206 4049
rect 11150 3975 11206 3984
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 10520 2582 10548 3334
rect 10980 3126 11008 3402
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 11072 2650 11100 3470
rect 11440 3194 11468 3606
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11808 3194 11836 3470
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10508 2576 10560 2582
rect 7102 2544 7158 2553
rect 7102 2479 7158 2488
rect 8298 2544 8354 2553
rect 10508 2518 10560 2524
rect 11242 2544 11298 2553
rect 8298 2479 8354 2488
rect 8576 2508 8628 2514
rect 7116 2446 7144 2479
rect 11242 2479 11244 2488
rect 8576 2450 8628 2456
rect 11296 2479 11298 2488
rect 11244 2450 11296 2456
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7930 2408 7986 2417
rect 7930 2343 7986 2352
rect 7024 2230 7144 2258
rect 5828 1822 6316 1850
rect 6288 480 6316 1822
rect 7116 480 7144 2230
rect 7944 480 7972 2343
rect 8588 2145 8616 2450
rect 9864 2440 9916 2446
rect 9862 2408 9864 2417
rect 9916 2408 9918 2417
rect 9862 2343 9918 2352
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8574 2136 8630 2145
rect 8574 2071 8630 2080
rect 8772 480 8800 2246
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 10414 1592 10470 1601
rect 10414 1527 10470 1536
rect 9586 1456 9642 1465
rect 9586 1391 9642 1400
rect 9600 480 9628 1391
rect 10428 480 10456 1527
rect 11348 480 11376 3062
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 12084 2553 12112 5510
rect 12268 4690 12296 8298
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12070 2544 12126 2553
rect 12070 2479 12126 2488
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 1465 11560 2246
rect 11518 1456 11574 1465
rect 11518 1391 11574 1400
rect 12176 480 12204 4422
rect 12268 4282 12296 4626
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12452 3754 12480 4966
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12360 3738 12480 3754
rect 12348 3732 12480 3738
rect 12400 3726 12480 3732
rect 12348 3674 12400 3680
rect 12544 3505 12572 4014
rect 12530 3496 12586 3505
rect 12530 3431 12586 3440
rect 12636 3097 12664 11630
rect 12728 3194 12756 14894
rect 12820 14414 12848 15302
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 14074 12848 14350
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12806 12336 12862 12345
rect 12806 12271 12808 12280
rect 12860 12271 12862 12280
rect 12808 12242 12860 12248
rect 12820 11898 12848 12242
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12912 5370 12940 22392
rect 13174 22264 13230 22273
rect 13174 22199 13230 22208
rect 13188 21146 13216 22199
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 13464 21690 13492 22102
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 13096 20874 13124 20946
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 13096 20602 13124 20810
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13004 14822 13032 15506
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 11694 13032 14758
rect 12992 11688 13044 11694
rect 13280 11665 13308 14894
rect 13464 14521 13492 20334
rect 13556 15162 13584 32166
rect 13636 28620 13688 28626
rect 13636 28562 13688 28568
rect 13648 28218 13676 28562
rect 13636 28212 13688 28218
rect 13636 28154 13688 28160
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13832 21690 13860 21966
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13924 20398 13952 34478
rect 15028 34241 15056 39520
rect 15672 35057 15700 39520
rect 15658 35048 15714 35057
rect 15658 34983 15714 34992
rect 15014 34232 15070 34241
rect 15014 34167 15070 34176
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13450 14512 13506 14521
rect 13450 14447 13506 14456
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 13358 13288 13414 13297
rect 13358 13223 13414 13232
rect 12992 11630 13044 11636
rect 13266 11656 13322 11665
rect 13266 11591 13322 11600
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12912 5166 12940 5306
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12900 3936 12952 3942
rect 13084 3936 13136 3942
rect 12952 3896 13032 3924
rect 12900 3878 12952 3884
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12622 3088 12678 3097
rect 12622 3023 12678 3032
rect 12728 2990 12756 3130
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12820 1601 12848 2246
rect 12806 1592 12862 1601
rect 12806 1527 12862 1536
rect 13004 480 13032 3896
rect 13084 3878 13136 3884
rect 13096 3534 13124 3878
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13188 2650 13216 10746
rect 13372 4690 13400 13223
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13266 4448 13322 4457
rect 13266 4383 13322 4392
rect 13280 3194 13308 4383
rect 13372 4282 13400 4626
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13464 3602 13492 5238
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13544 4072 13596 4078
rect 13542 4040 13544 4049
rect 13596 4040 13598 4049
rect 13542 3975 13598 3984
rect 13542 3632 13598 3641
rect 13452 3596 13504 3602
rect 13542 3567 13598 3576
rect 13452 3538 13504 3544
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13464 3126 13492 3538
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13556 2990 13584 3567
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13648 2825 13676 3334
rect 13634 2816 13690 2825
rect 13634 2751 13690 2760
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13832 480 13860 4490
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14660 480 14688 4422
rect 15474 2816 15530 2825
rect 15474 2751 15530 2760
rect 15488 480 15516 2751
rect 386 0 442 480
rect 1214 0 1270 480
rect 2042 0 2098 480
rect 2870 0 2926 480
rect 3698 0 3754 480
rect 4526 0 4582 480
rect 5354 0 5410 480
rect 6274 0 6330 480
rect 7102 0 7158 480
rect 7930 0 7986 480
rect 8758 0 8814 480
rect 9586 0 9642 480
rect 10414 0 10470 480
rect 11334 0 11390 480
rect 12162 0 12218 480
rect 12990 0 13046 480
rect 13818 0 13874 480
rect 14646 0 14702 480
rect 15474 0 15530 480
<< via2 >>
rect 294 34720 350 34776
rect 1490 35536 1546 35592
rect 846 34584 902 34640
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3330 34992 3386 35048
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3146 34720 3202 34776
rect 3514 34584 3570 34640
rect 4158 34584 4214 34640
rect 3146 29144 3202 29200
rect 3054 29028 3110 29064
rect 3054 29008 3056 29028
rect 3056 29008 3108 29028
rect 3108 29008 3110 29028
rect 4066 33904 4122 33960
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3882 33496 3938 33552
rect 4250 33360 4306 33416
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 4526 34992 4582 35048
rect 4434 32952 4490 33008
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 4526 29552 4582 29608
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 2686 27512 2742 27568
rect 2962 24268 3018 24304
rect 2962 24248 2964 24268
rect 2964 24248 3016 24268
rect 3016 24248 3018 24268
rect 2870 20052 2926 20088
rect 2870 20032 2872 20052
rect 2872 20032 2924 20052
rect 2924 20032 2926 20052
rect 2870 18672 2926 18728
rect 2870 15952 2926 16008
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3974 24112 4030 24168
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3238 23704 3294 23760
rect 3146 22500 3202 22536
rect 3146 22480 3148 22500
rect 3148 22480 3200 22500
rect 3200 22480 3202 22500
rect 2962 10104 3018 10160
rect 3146 17740 3202 17776
rect 3146 17720 3148 17740
rect 3148 17720 3200 17740
rect 3200 17720 3202 17740
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3974 22652 3976 22672
rect 3976 22652 4028 22672
rect 4028 22652 4030 22672
rect 3974 22616 4030 22652
rect 4158 22752 4214 22808
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3974 18808 4030 18864
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 4342 24692 4344 24712
rect 4344 24692 4396 24712
rect 4396 24692 4398 24712
rect 4342 24656 4398 24692
rect 4526 22072 4582 22128
rect 5446 35536 5502 35592
rect 5170 34584 5226 34640
rect 5262 33396 5264 33416
rect 5264 33396 5316 33416
rect 5316 33396 5318 33416
rect 5262 33360 5318 33396
rect 4986 31864 5042 31920
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6274 34992 6330 35048
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 5354 31728 5410 31784
rect 5078 29008 5134 29064
rect 4894 27376 4950 27432
rect 4710 22616 4766 22672
rect 5630 31728 5686 31784
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6458 30796 6514 30832
rect 6458 30776 6460 30796
rect 6460 30776 6512 30796
rect 6512 30776 6514 30796
rect 6090 30640 6146 30696
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 5814 26832 5870 26888
rect 5446 24828 5448 24848
rect 5448 24828 5500 24848
rect 5500 24828 5502 24848
rect 5446 24792 5502 24828
rect 5722 24112 5778 24168
rect 4342 18128 4398 18184
rect 4250 17332 4306 17368
rect 4250 17312 4252 17332
rect 4252 17312 4304 17332
rect 4304 17312 4306 17332
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3974 15408 4030 15464
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3422 15000 3478 15056
rect 4066 14320 4122 14376
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 4066 13812 4068 13832
rect 4068 13812 4120 13832
rect 4120 13812 4122 13832
rect 4066 13776 4122 13812
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 4066 6704 4122 6760
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 4434 14456 4490 14512
rect 4434 13368 4490 13424
rect 4526 10124 4582 10160
rect 4526 10104 4528 10124
rect 4528 10104 4580 10124
rect 4580 10104 4582 10124
rect 4710 20304 4766 20360
rect 4986 19796 4988 19816
rect 4988 19796 5040 19816
rect 5040 19796 5042 19816
rect 4986 19760 5042 19796
rect 5078 14864 5134 14920
rect 5078 13232 5134 13288
rect 5814 23160 5870 23216
rect 5814 22772 5870 22808
rect 5814 22752 5816 22772
rect 5816 22752 5868 22772
rect 5868 22752 5870 22772
rect 5446 16652 5502 16688
rect 5446 16632 5448 16652
rect 5448 16632 5500 16652
rect 5500 16632 5502 16652
rect 5262 15272 5318 15328
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6182 23568 6238 23624
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6918 35536 6974 35592
rect 6826 29960 6882 30016
rect 7286 35536 7342 35592
rect 7470 34584 7526 34640
rect 7286 29144 7342 29200
rect 7562 33360 7618 33416
rect 8298 35672 8354 35728
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8114 30640 8170 30696
rect 6918 24792 6974 24848
rect 6734 23432 6790 23488
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 5998 18400 6054 18456
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 5078 11736 5134 11792
rect 5078 7948 5134 7984
rect 5078 7928 5080 7948
rect 5080 7928 5132 7948
rect 5132 7928 5134 7948
rect 2042 3032 2098 3088
rect 1214 2760 1270 2816
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3698 2932 3700 2952
rect 3700 2932 3752 2952
rect 3752 2932 3754 2952
rect 3698 2896 3754 2932
rect 4250 2760 4306 2816
rect 3514 2488 3570 2544
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 5814 17040 5870 17096
rect 5446 7384 5502 7440
rect 5170 5208 5226 5264
rect 5262 5072 5318 5128
rect 4618 4256 4674 4312
rect 4986 3168 5042 3224
rect 5446 3304 5502 3360
rect 5354 2760 5410 2816
rect 5078 2216 5134 2272
rect 5538 2080 5594 2136
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6642 15544 6698 15600
rect 6642 15408 6698 15464
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6458 14356 6460 14376
rect 6460 14356 6512 14376
rect 6512 14356 6514 14376
rect 6458 14320 6514 14356
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 7194 24248 7250 24304
rect 7102 24112 7158 24168
rect 7286 23740 7288 23760
rect 7288 23740 7340 23760
rect 7340 23740 7342 23760
rect 7286 23704 7342 23740
rect 7194 22636 7250 22672
rect 7194 22616 7196 22636
rect 7196 22616 7248 22636
rect 7248 22616 7250 22636
rect 7194 21936 7250 21992
rect 7746 24812 7802 24848
rect 7746 24792 7748 24812
rect 7748 24792 7800 24812
rect 7800 24792 7802 24812
rect 7286 20848 7342 20904
rect 7838 24268 7894 24304
rect 7838 24248 7840 24268
rect 7840 24248 7892 24268
rect 7892 24248 7894 24268
rect 7194 18264 7250 18320
rect 7102 17040 7158 17096
rect 6826 16788 6882 16824
rect 6826 16768 6828 16788
rect 6828 16768 6880 16788
rect 6880 16768 6882 16788
rect 6090 11636 6092 11656
rect 6092 11636 6144 11656
rect 6144 11636 6146 11656
rect 6090 11600 6146 11636
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6550 11056 6606 11112
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6274 5364 6330 5400
rect 6274 5344 6276 5364
rect 6276 5344 6328 5364
rect 6328 5344 6330 5364
rect 6918 13796 6974 13832
rect 6918 13776 6920 13796
rect 6920 13776 6972 13796
rect 6972 13776 6974 13796
rect 7562 18808 7618 18864
rect 8390 29996 8392 30016
rect 8392 29996 8444 30016
rect 8444 29996 8446 30016
rect 8390 29960 8446 29996
rect 8298 24656 8354 24712
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8758 32952 8814 33008
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8850 32272 8906 32328
rect 8666 30776 8722 30832
rect 8666 28464 8722 28520
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 9770 35128 9826 35184
rect 9494 33904 9550 33960
rect 10966 36916 11022 36952
rect 10966 36896 10968 36916
rect 10968 36896 11020 36916
rect 11020 36896 11022 36916
rect 10230 35572 10232 35592
rect 10232 35572 10284 35592
rect 10284 35572 10286 35592
rect 10230 35536 10286 35572
rect 10966 34620 10968 34640
rect 10968 34620 11020 34640
rect 11020 34620 11022 34640
rect 10966 34584 11022 34620
rect 10506 33516 10562 33552
rect 10506 33496 10508 33516
rect 10508 33496 10560 33516
rect 10560 33496 10562 33516
rect 10046 32428 10102 32464
rect 10046 32408 10048 32428
rect 10048 32408 10100 32428
rect 10100 32408 10102 32428
rect 10046 31864 10102 31920
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 12070 37440 12126 37496
rect 11978 36896 12034 36952
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 9954 30640 10010 30696
rect 9954 29008 10010 29064
rect 9494 27784 9550 27840
rect 9494 27376 9550 27432
rect 9494 27276 9496 27296
rect 9496 27276 9548 27296
rect 9548 27276 9550 27296
rect 9494 27240 9550 27276
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8758 26424 8814 26480
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8574 24556 8576 24576
rect 8576 24556 8628 24576
rect 8628 24556 8630 24576
rect 8574 24520 8630 24556
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8758 23740 8760 23760
rect 8760 23740 8812 23760
rect 8812 23740 8814 23760
rect 8758 23704 8814 23740
rect 8574 23604 8576 23624
rect 8576 23604 8628 23624
rect 8628 23604 8630 23624
rect 8574 23568 8630 23604
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8850 22072 8906 22128
rect 8022 19080 8078 19136
rect 8298 18672 8354 18728
rect 8666 20168 8722 20224
rect 7838 17312 7894 17368
rect 7838 15272 7894 15328
rect 7194 9152 7250 9208
rect 7010 7928 7066 7984
rect 8022 14456 8078 14512
rect 8574 17992 8630 18048
rect 8758 19760 8814 19816
rect 8758 18420 8814 18456
rect 8758 18400 8760 18420
rect 8760 18400 8812 18420
rect 8812 18400 8814 18420
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 10230 27240 10286 27296
rect 9586 23976 9642 24032
rect 9678 23468 9680 23488
rect 9680 23468 9732 23488
rect 9732 23468 9734 23488
rect 9678 23432 9734 23468
rect 9678 21972 9680 21992
rect 9680 21972 9732 21992
rect 9732 21972 9734 21992
rect 9678 21936 9734 21972
rect 10230 20848 10286 20904
rect 9770 19116 9772 19136
rect 9772 19116 9824 19136
rect 9824 19116 9826 19136
rect 9770 19080 9826 19116
rect 11058 29552 11114 29608
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 12070 35284 12126 35320
rect 12070 35264 12072 35284
rect 12072 35264 12124 35284
rect 12124 35264 12126 35284
rect 12070 35128 12126 35184
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11978 28464 12034 28520
rect 11426 27820 11428 27840
rect 11428 27820 11480 27840
rect 11480 27820 11482 27840
rect 11426 27784 11482 27820
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11242 24520 11298 24576
rect 11058 23976 11114 24032
rect 10414 23060 10416 23080
rect 10416 23060 10468 23080
rect 10468 23060 10470 23080
rect 10414 23024 10470 23060
rect 9310 17720 9366 17776
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8850 16904 8906 16960
rect 9770 16768 9826 16824
rect 8850 16632 8906 16688
rect 8666 16088 8722 16144
rect 8666 15952 8722 16008
rect 8482 15564 8538 15600
rect 8482 15544 8484 15564
rect 8484 15544 8536 15564
rect 8536 15544 8538 15564
rect 7378 9016 7434 9072
rect 7194 7384 7250 7440
rect 7010 5344 7066 5400
rect 6734 5072 6790 5128
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6090 4120 6146 4176
rect 6090 3440 6146 3496
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 6918 3304 6974 3360
rect 5906 2352 5962 2408
rect 8390 13368 8446 13424
rect 8390 12688 8446 12744
rect 7746 10648 7802 10704
rect 7654 5344 7710 5400
rect 8022 4528 8078 4584
rect 7286 3712 7342 3768
rect 7470 3340 7472 3360
rect 7472 3340 7524 3360
rect 7524 3340 7526 3360
rect 7470 3304 7526 3340
rect 7838 3596 7894 3632
rect 7838 3576 7840 3596
rect 7840 3576 7892 3596
rect 7892 3576 7894 3596
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8574 13368 8630 13424
rect 8574 12144 8630 12200
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 9862 14864 9918 14920
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8850 11056 8906 11112
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 9402 10784 9458 10840
rect 9586 11192 9642 11248
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8758 9172 8814 9208
rect 8758 9152 8760 9172
rect 8760 9152 8812 9172
rect 8812 9152 8814 9172
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8850 7248 8906 7304
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8482 4256 8538 4312
rect 8666 3848 8722 3904
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 9862 11056 9918 11112
rect 10690 18828 10746 18864
rect 10690 18808 10692 18828
rect 10692 18808 10744 18828
rect 10744 18808 10746 18828
rect 10874 20712 10930 20768
rect 11426 26868 11428 26888
rect 11428 26868 11480 26888
rect 11480 26868 11482 26888
rect 11426 26832 11482 26868
rect 11978 27376 12034 27432
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 12438 34856 12494 34912
rect 12622 34584 12678 34640
rect 12898 32408 12954 32464
rect 12438 31864 12494 31920
rect 13174 35264 13230 35320
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 13634 34992 13690 35048
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 13542 34196 13598 34232
rect 13542 34176 13544 34196
rect 13544 34176 13596 34196
rect 13596 34176 13598 34196
rect 13450 29144 13506 29200
rect 12990 29028 13046 29064
rect 12990 29008 12992 29028
rect 12992 29008 13044 29028
rect 13044 29008 13046 29028
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 12070 24384 12126 24440
rect 11978 23704 12034 23760
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11978 23196 11980 23216
rect 11980 23196 12032 23216
rect 12032 23196 12034 23216
rect 11978 23160 12034 23196
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11518 22072 11574 22128
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11058 18944 11114 19000
rect 10874 18264 10930 18320
rect 11150 18164 11152 18184
rect 11152 18164 11204 18184
rect 11204 18164 11206 18184
rect 11150 18128 11206 18164
rect 11150 18028 11152 18048
rect 11152 18028 11204 18048
rect 11204 18028 11206 18048
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11150 17992 11206 18028
rect 10874 16088 10930 16144
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 12438 27240 12494 27296
rect 12530 24792 12586 24848
rect 13082 27532 13138 27568
rect 13082 27512 13084 27532
rect 13084 27512 13136 27532
rect 13136 27512 13138 27532
rect 12714 24384 12770 24440
rect 12530 24112 12586 24168
rect 12622 23740 12624 23760
rect 12624 23740 12676 23760
rect 12676 23740 12678 23760
rect 12622 23704 12678 23740
rect 12898 23024 12954 23080
rect 13082 22480 13138 22536
rect 12530 20712 12586 20768
rect 12530 20340 12532 20360
rect 12532 20340 12584 20360
rect 12584 20340 12586 20360
rect 12530 20304 12586 20340
rect 12714 17176 12770 17232
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 12714 15000 12770 15056
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11150 13388 11206 13424
rect 11150 13368 11152 13388
rect 11152 13368 11204 13388
rect 11204 13368 11206 13388
rect 10874 13232 10930 13288
rect 11150 12724 11152 12744
rect 11152 12724 11204 12744
rect 11204 12724 11206 12744
rect 11150 12688 11206 12724
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 12070 12416 12126 12472
rect 11242 11736 11298 11792
rect 11058 10648 11114 10704
rect 10690 9036 10746 9072
rect 10690 9016 10692 9036
rect 10692 9016 10744 9036
rect 10744 9016 10746 9036
rect 11150 7284 11152 7304
rect 11152 7284 11204 7304
rect 11204 7284 11206 7304
rect 11150 7248 11206 7284
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 12438 10784 12494 10840
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11702 7420 11704 7440
rect 11704 7420 11756 7440
rect 11756 7420 11758 7440
rect 11702 7384 11758 7420
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 9678 4528 9734 4584
rect 8666 3168 8722 3224
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8298 2896 8354 2952
rect 9586 3712 9642 3768
rect 9770 3576 9826 3632
rect 10230 4140 10286 4176
rect 10230 4120 10232 4140
rect 10232 4120 10284 4140
rect 10284 4120 10286 4140
rect 10782 4428 10784 4448
rect 10784 4428 10836 4448
rect 10836 4428 10838 4448
rect 10782 4392 10838 4428
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11242 5244 11244 5264
rect 11244 5244 11296 5264
rect 11296 5244 11298 5264
rect 11242 5208 11298 5244
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11150 3984 11206 4040
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 7102 2488 7158 2544
rect 8298 2488 8354 2544
rect 11242 2508 11298 2544
rect 11242 2488 11244 2508
rect 11244 2488 11296 2508
rect 11296 2488 11298 2508
rect 7930 2352 7986 2408
rect 9862 2388 9864 2408
rect 9864 2388 9916 2408
rect 9916 2388 9918 2408
rect 9862 2352 9918 2388
rect 8574 2080 8630 2136
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 10414 1536 10470 1592
rect 9586 1400 9642 1456
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12070 2488 12126 2544
rect 11518 1400 11574 1456
rect 12530 3440 12586 3496
rect 12806 12300 12862 12336
rect 12806 12280 12808 12300
rect 12808 12280 12860 12300
rect 12860 12280 12862 12300
rect 13174 22208 13230 22264
rect 15658 34992 15714 35048
rect 15014 34176 15070 34232
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 13450 14456 13506 14512
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 13358 13232 13414 13288
rect 13266 11600 13322 11656
rect 12622 3032 12678 3088
rect 12806 1536 12862 1592
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 13266 4392 13322 4448
rect 13542 4020 13544 4040
rect 13544 4020 13596 4040
rect 13596 4020 13598 4040
rect 13542 3984 13598 4020
rect 13542 3576 13598 3632
rect 13634 2760 13690 2816
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 15474 2760 15530 2816
<< metal3 >>
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 12065 37498 12131 37501
rect 15520 37498 16000 37528
rect 12065 37496 16000 37498
rect 12065 37440 12070 37496
rect 12126 37440 16000 37496
rect 12065 37438 16000 37440
rect 12065 37435 12131 37438
rect 15520 37408 16000 37438
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 10961 36954 11027 36957
rect 11973 36954 12039 36957
rect 10961 36952 12039 36954
rect 10961 36896 10966 36952
rect 11022 36896 11978 36952
rect 12034 36896 12039 36952
rect 10961 36894 12039 36896
rect 10961 36891 11027 36894
rect 11973 36891 12039 36894
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 8293 35730 8359 35733
rect 5214 35728 8359 35730
rect 5214 35672 8298 35728
rect 8354 35672 8359 35728
rect 5214 35670 8359 35672
rect 1485 35594 1551 35597
rect 5214 35594 5274 35670
rect 8293 35667 8359 35670
rect 1485 35592 5274 35594
rect 1485 35536 1490 35592
rect 1546 35536 5274 35592
rect 1485 35534 5274 35536
rect 5441 35594 5507 35597
rect 6913 35594 6979 35597
rect 5441 35592 6979 35594
rect 5441 35536 5446 35592
rect 5502 35536 6918 35592
rect 6974 35536 6979 35592
rect 5441 35534 6979 35536
rect 1485 35531 1551 35534
rect 5441 35531 5507 35534
rect 6913 35531 6979 35534
rect 7281 35594 7347 35597
rect 10225 35594 10291 35597
rect 7281 35592 10291 35594
rect 7281 35536 7286 35592
rect 7342 35536 10230 35592
rect 10286 35536 10291 35592
rect 7281 35534 10291 35536
rect 7281 35531 7347 35534
rect 10225 35531 10291 35534
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 12065 35322 12131 35325
rect 13169 35322 13235 35325
rect 12065 35320 13235 35322
rect 12065 35264 12070 35320
rect 12126 35264 13174 35320
rect 13230 35264 13235 35320
rect 12065 35262 13235 35264
rect 12065 35259 12131 35262
rect 13169 35259 13235 35262
rect 9765 35186 9831 35189
rect 12065 35186 12131 35189
rect 9765 35184 12131 35186
rect 9765 35128 9770 35184
rect 9826 35128 12070 35184
rect 12126 35128 12131 35184
rect 9765 35126 12131 35128
rect 9765 35123 9831 35126
rect 12065 35123 12131 35126
rect 3325 35050 3391 35053
rect 4521 35050 4587 35053
rect 3325 35048 4587 35050
rect 3325 34992 3330 35048
rect 3386 34992 4526 35048
rect 4582 34992 4587 35048
rect 3325 34990 4587 34992
rect 3325 34987 3391 34990
rect 4521 34987 4587 34990
rect 6269 35050 6335 35053
rect 13629 35050 13695 35053
rect 15653 35050 15719 35053
rect 6269 35048 9506 35050
rect 6269 34992 6274 35048
rect 6330 34992 9506 35048
rect 6269 34990 9506 34992
rect 6269 34987 6335 34990
rect 9446 34916 9506 34990
rect 13629 35048 15719 35050
rect 13629 34992 13634 35048
rect 13690 34992 15658 35048
rect 15714 34992 15719 35048
rect 13629 34990 15719 34992
rect 13629 34987 13695 34990
rect 15653 34987 15719 34990
rect 9438 34852 9444 34916
rect 9508 34914 9514 34916
rect 12433 34914 12499 34917
rect 9508 34912 12499 34914
rect 9508 34856 12438 34912
rect 12494 34856 12499 34912
rect 9508 34854 12499 34856
rect 9508 34852 9514 34854
rect 12433 34851 12499 34854
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 289 34778 355 34781
rect 3141 34778 3207 34781
rect 289 34776 3207 34778
rect 289 34720 294 34776
rect 350 34720 3146 34776
rect 3202 34720 3207 34776
rect 289 34718 3207 34720
rect 289 34715 355 34718
rect 3141 34715 3207 34718
rect 841 34642 907 34645
rect 3509 34642 3575 34645
rect 4153 34642 4219 34645
rect 841 34640 4219 34642
rect 841 34584 846 34640
rect 902 34584 3514 34640
rect 3570 34584 4158 34640
rect 4214 34584 4219 34640
rect 841 34582 4219 34584
rect 841 34579 907 34582
rect 3509 34579 3575 34582
rect 4153 34579 4219 34582
rect 5165 34642 5231 34645
rect 7465 34642 7531 34645
rect 5165 34640 7531 34642
rect 5165 34584 5170 34640
rect 5226 34584 7470 34640
rect 7526 34584 7531 34640
rect 5165 34582 7531 34584
rect 5165 34579 5231 34582
rect 7465 34579 7531 34582
rect 10961 34642 11027 34645
rect 12617 34642 12683 34645
rect 10961 34640 12683 34642
rect 10961 34584 10966 34640
rect 11022 34584 12622 34640
rect 12678 34584 12683 34640
rect 10961 34582 12683 34584
rect 10961 34579 11027 34582
rect 12617 34579 12683 34582
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 13537 34234 13603 34237
rect 15009 34234 15075 34237
rect 13537 34232 15075 34234
rect 13537 34176 13542 34232
rect 13598 34176 15014 34232
rect 15070 34176 15075 34232
rect 13537 34174 15075 34176
rect 13537 34171 13603 34174
rect 15009 34171 15075 34174
rect 4061 33962 4127 33965
rect 9489 33962 9555 33965
rect 4061 33960 9555 33962
rect 4061 33904 4066 33960
rect 4122 33904 9494 33960
rect 9550 33904 9555 33960
rect 4061 33902 9555 33904
rect 4061 33899 4127 33902
rect 9489 33899 9555 33902
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 3877 33554 3943 33557
rect 10501 33554 10567 33557
rect 3877 33552 10567 33554
rect 3877 33496 3882 33552
rect 3938 33496 10506 33552
rect 10562 33496 10567 33552
rect 3877 33494 10567 33496
rect 3877 33491 3943 33494
rect 10501 33491 10567 33494
rect 0 33418 480 33448
rect 4245 33418 4311 33421
rect 0 33416 4311 33418
rect 0 33360 4250 33416
rect 4306 33360 4311 33416
rect 0 33358 4311 33360
rect 0 33328 480 33358
rect 4245 33355 4311 33358
rect 5257 33418 5323 33421
rect 7557 33418 7623 33421
rect 5257 33416 7623 33418
rect 5257 33360 5262 33416
rect 5318 33360 7562 33416
rect 7618 33360 7623 33416
rect 5257 33358 7623 33360
rect 5257 33355 5323 33358
rect 7557 33355 7623 33358
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 4429 33010 4495 33013
rect 8753 33010 8819 33013
rect 4429 33008 8819 33010
rect 4429 32952 4434 33008
rect 4490 32952 8758 33008
rect 8814 32952 8819 33008
rect 4429 32950 8819 32952
rect 4429 32947 4495 32950
rect 8753 32947 8819 32950
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 10041 32466 10107 32469
rect 12893 32466 12959 32469
rect 15520 32466 16000 32496
rect 10041 32464 12959 32466
rect 10041 32408 10046 32464
rect 10102 32408 12898 32464
rect 12954 32408 12959 32464
rect 10041 32406 12959 32408
rect 10041 32403 10107 32406
rect 12893 32403 12959 32406
rect 13126 32406 16000 32466
rect 8845 32330 8911 32333
rect 13126 32330 13186 32406
rect 15520 32376 16000 32406
rect 8845 32328 13186 32330
rect 8845 32272 8850 32328
rect 8906 32272 13186 32328
rect 8845 32270 13186 32272
rect 8845 32267 8911 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 4981 31922 5047 31925
rect 10041 31922 10107 31925
rect 12433 31922 12499 31925
rect 4981 31920 12499 31922
rect 4981 31864 4986 31920
rect 5042 31864 10046 31920
rect 10102 31864 12438 31920
rect 12494 31864 12499 31920
rect 4981 31862 12499 31864
rect 4981 31859 5047 31862
rect 10041 31859 10107 31862
rect 12433 31859 12499 31862
rect 5349 31786 5415 31789
rect 5625 31786 5691 31789
rect 5349 31784 5691 31786
rect 5349 31728 5354 31784
rect 5410 31728 5630 31784
rect 5686 31728 5691 31784
rect 5349 31726 5691 31728
rect 5349 31723 5415 31726
rect 5625 31723 5691 31726
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 6453 30834 6519 30837
rect 8661 30834 8727 30837
rect 6453 30832 8727 30834
rect 6453 30776 6458 30832
rect 6514 30776 8666 30832
rect 8722 30776 8727 30832
rect 6453 30774 8727 30776
rect 6453 30771 6519 30774
rect 8661 30771 8727 30774
rect 6085 30698 6151 30701
rect 8109 30698 8175 30701
rect 9949 30698 10015 30701
rect 6085 30696 10015 30698
rect 6085 30640 6090 30696
rect 6146 30640 8114 30696
rect 8170 30640 9954 30696
rect 10010 30640 10015 30696
rect 6085 30638 10015 30640
rect 6085 30635 6151 30638
rect 8109 30635 8175 30638
rect 9949 30635 10015 30638
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 6821 30018 6887 30021
rect 8385 30018 8451 30021
rect 6821 30016 8451 30018
rect 6821 29960 6826 30016
rect 6882 29960 8390 30016
rect 8446 29960 8451 30016
rect 6821 29958 8451 29960
rect 6821 29955 6887 29958
rect 8385 29955 8451 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 4521 29610 4587 29613
rect 11053 29610 11119 29613
rect 4521 29608 11119 29610
rect 4521 29552 4526 29608
rect 4582 29552 11058 29608
rect 11114 29552 11119 29608
rect 4521 29550 11119 29552
rect 4521 29547 4587 29550
rect 11053 29547 11119 29550
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 7054 29278 7482 29338
rect 3141 29202 3207 29205
rect 7054 29202 7114 29278
rect 7281 29202 7347 29205
rect 3141 29200 7114 29202
rect 3141 29144 3146 29200
rect 3202 29144 7114 29200
rect 3141 29142 7114 29144
rect 7238 29200 7347 29202
rect 7238 29144 7286 29200
rect 7342 29144 7347 29200
rect 3141 29139 3207 29142
rect 7238 29139 7347 29144
rect 7422 29202 7482 29278
rect 13445 29202 13511 29205
rect 7422 29200 13511 29202
rect 7422 29144 13450 29200
rect 13506 29144 13511 29200
rect 7422 29142 13511 29144
rect 13445 29139 13511 29142
rect 3049 29066 3115 29069
rect 5073 29066 5139 29069
rect 7238 29066 7298 29139
rect 3049 29064 7298 29066
rect 3049 29008 3054 29064
rect 3110 29008 5078 29064
rect 5134 29008 7298 29064
rect 3049 29006 7298 29008
rect 9949 29066 10015 29069
rect 12985 29066 13051 29069
rect 9949 29064 13051 29066
rect 9949 29008 9954 29064
rect 10010 29008 12990 29064
rect 13046 29008 13051 29064
rect 9949 29006 13051 29008
rect 3049 29003 3115 29006
rect 5073 29003 5139 29006
rect 9949 29003 10015 29006
rect 12985 29003 13051 29006
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 8661 28522 8727 28525
rect 11973 28522 12039 28525
rect 8661 28520 12039 28522
rect 8661 28464 8666 28520
rect 8722 28464 11978 28520
rect 12034 28464 12039 28520
rect 8661 28462 12039 28464
rect 8661 28459 8727 28462
rect 11973 28459 12039 28462
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 9489 27842 9555 27845
rect 11421 27842 11487 27845
rect 9489 27840 11487 27842
rect 9489 27784 9494 27840
rect 9550 27784 11426 27840
rect 11482 27784 11487 27840
rect 9489 27782 11487 27784
rect 9489 27779 9555 27782
rect 11421 27779 11487 27782
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 2681 27570 2747 27573
rect 13077 27570 13143 27573
rect 2681 27568 13143 27570
rect 2681 27512 2686 27568
rect 2742 27512 13082 27568
rect 13138 27512 13143 27568
rect 2681 27510 13143 27512
rect 2681 27507 2747 27510
rect 13077 27507 13143 27510
rect 4889 27434 4955 27437
rect 9489 27434 9555 27437
rect 4889 27432 9555 27434
rect 4889 27376 4894 27432
rect 4950 27376 9494 27432
rect 9550 27376 9555 27432
rect 4889 27374 9555 27376
rect 4889 27371 4955 27374
rect 9489 27371 9555 27374
rect 11973 27434 12039 27437
rect 15520 27434 16000 27464
rect 11973 27432 16000 27434
rect 11973 27376 11978 27432
rect 12034 27376 16000 27432
rect 11973 27374 16000 27376
rect 11973 27371 12039 27374
rect 15520 27344 16000 27374
rect 9489 27298 9555 27301
rect 10225 27298 10291 27301
rect 12433 27298 12499 27301
rect 9489 27296 12499 27298
rect 9489 27240 9494 27296
rect 9550 27240 10230 27296
rect 10286 27240 12438 27296
rect 12494 27240 12499 27296
rect 9489 27238 12499 27240
rect 9489 27235 9555 27238
rect 10225 27235 10291 27238
rect 12433 27235 12499 27238
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 5809 26890 5875 26893
rect 11421 26890 11487 26893
rect 5809 26888 11487 26890
rect 5809 26832 5814 26888
rect 5870 26832 11426 26888
rect 11482 26832 11487 26888
rect 5809 26830 11487 26832
rect 5809 26827 5875 26830
rect 11421 26827 11487 26830
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 8753 26484 8819 26485
rect 8702 26482 8708 26484
rect 8662 26422 8708 26482
rect 8772 26480 8819 26484
rect 8814 26424 8819 26480
rect 8702 26420 8708 26422
rect 8772 26420 8819 26424
rect 8753 26419 8819 26420
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 5441 24850 5507 24853
rect 6913 24850 6979 24853
rect 5441 24848 6979 24850
rect 5441 24792 5446 24848
rect 5502 24792 6918 24848
rect 6974 24792 6979 24848
rect 5441 24790 6979 24792
rect 5441 24787 5507 24790
rect 6913 24787 6979 24790
rect 7741 24850 7807 24853
rect 12525 24850 12591 24853
rect 7741 24848 12591 24850
rect 7741 24792 7746 24848
rect 7802 24792 12530 24848
rect 12586 24792 12591 24848
rect 7741 24790 12591 24792
rect 7741 24787 7807 24790
rect 12525 24787 12591 24790
rect 4337 24714 4403 24717
rect 8293 24714 8359 24717
rect 4337 24712 8359 24714
rect 4337 24656 4342 24712
rect 4398 24656 8298 24712
rect 8354 24656 8359 24712
rect 4337 24654 8359 24656
rect 4337 24651 4403 24654
rect 8293 24651 8359 24654
rect 8569 24578 8635 24581
rect 11237 24578 11303 24581
rect 8569 24576 11303 24578
rect 8569 24520 8574 24576
rect 8630 24520 11242 24576
rect 11298 24520 11303 24576
rect 8569 24518 11303 24520
rect 8569 24515 8635 24518
rect 11237 24515 11303 24518
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 12065 24442 12131 24445
rect 12709 24442 12775 24445
rect 12022 24440 12775 24442
rect 12022 24384 12070 24440
rect 12126 24384 12714 24440
rect 12770 24384 12775 24440
rect 12022 24382 12775 24384
rect 12022 24379 12131 24382
rect 12709 24379 12775 24382
rect 2957 24306 3023 24309
rect 7189 24306 7255 24309
rect 2957 24304 7255 24306
rect 2957 24248 2962 24304
rect 3018 24248 7194 24304
rect 7250 24248 7255 24304
rect 2957 24246 7255 24248
rect 2957 24243 3023 24246
rect 7189 24243 7255 24246
rect 7833 24306 7899 24309
rect 12022 24306 12082 24379
rect 7833 24304 12082 24306
rect 7833 24248 7838 24304
rect 7894 24248 12082 24304
rect 7833 24246 12082 24248
rect 7833 24243 7899 24246
rect 3969 24170 4035 24173
rect 5717 24170 5783 24173
rect 3969 24168 5783 24170
rect 3969 24112 3974 24168
rect 4030 24112 5722 24168
rect 5778 24112 5783 24168
rect 3969 24110 5783 24112
rect 3969 24107 4035 24110
rect 5717 24107 5783 24110
rect 7097 24170 7163 24173
rect 12525 24170 12591 24173
rect 7097 24168 12591 24170
rect 7097 24112 7102 24168
rect 7158 24112 12530 24168
rect 12586 24112 12591 24168
rect 7097 24110 12591 24112
rect 7097 24107 7163 24110
rect 12525 24107 12591 24110
rect 9581 24034 9647 24037
rect 11053 24034 11119 24037
rect 9581 24032 11119 24034
rect 9581 23976 9586 24032
rect 9642 23976 11058 24032
rect 11114 23976 11119 24032
rect 9581 23974 11119 23976
rect 9581 23971 9647 23974
rect 11053 23971 11119 23974
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 3233 23762 3299 23765
rect 7281 23762 7347 23765
rect 3233 23760 7347 23762
rect 3233 23704 3238 23760
rect 3294 23704 7286 23760
rect 7342 23704 7347 23760
rect 3233 23702 7347 23704
rect 3233 23699 3299 23702
rect 7281 23699 7347 23702
rect 8753 23762 8819 23765
rect 11973 23762 12039 23765
rect 12617 23762 12683 23765
rect 8753 23760 12683 23762
rect 8753 23704 8758 23760
rect 8814 23704 11978 23760
rect 12034 23704 12622 23760
rect 12678 23704 12683 23760
rect 8753 23702 12683 23704
rect 8753 23699 8819 23702
rect 11973 23699 12039 23702
rect 12617 23699 12683 23702
rect 6177 23626 6243 23629
rect 8569 23626 8635 23629
rect 6177 23624 8635 23626
rect 6177 23568 6182 23624
rect 6238 23568 8574 23624
rect 8630 23568 8635 23624
rect 6177 23566 8635 23568
rect 6177 23563 6243 23566
rect 8569 23563 8635 23566
rect 6729 23490 6795 23493
rect 9673 23490 9739 23493
rect 6729 23488 9739 23490
rect 6729 23432 6734 23488
rect 6790 23432 9678 23488
rect 9734 23432 9739 23488
rect 6729 23430 9739 23432
rect 6729 23427 6795 23430
rect 9673 23427 9739 23430
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 5809 23218 5875 23221
rect 11973 23218 12039 23221
rect 5809 23216 12039 23218
rect 5809 23160 5814 23216
rect 5870 23160 11978 23216
rect 12034 23160 12039 23216
rect 5809 23158 12039 23160
rect 5809 23155 5875 23158
rect 11973 23155 12039 23158
rect 10409 23082 10475 23085
rect 12893 23082 12959 23085
rect 10409 23080 12959 23082
rect 10409 23024 10414 23080
rect 10470 23024 12898 23080
rect 12954 23024 12959 23080
rect 10409 23022 12959 23024
rect 10409 23019 10475 23022
rect 12893 23019 12959 23022
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 4153 22810 4219 22813
rect 5809 22810 5875 22813
rect 4153 22808 5875 22810
rect 4153 22752 4158 22808
rect 4214 22752 5814 22808
rect 5870 22752 5875 22808
rect 4153 22750 5875 22752
rect 4153 22747 4219 22750
rect 5809 22747 5875 22750
rect 3969 22674 4035 22677
rect 4705 22674 4771 22677
rect 7189 22674 7255 22677
rect 3969 22672 7255 22674
rect 3969 22616 3974 22672
rect 4030 22616 4710 22672
rect 4766 22616 7194 22672
rect 7250 22616 7255 22672
rect 3969 22614 7255 22616
rect 3969 22611 4035 22614
rect 4705 22611 4771 22614
rect 7189 22611 7255 22614
rect 3141 22538 3207 22541
rect 13077 22538 13143 22541
rect 15520 22538 16000 22568
rect 3141 22536 13143 22538
rect 3141 22480 3146 22536
rect 3202 22480 13082 22536
rect 13138 22480 13143 22536
rect 3141 22478 13143 22480
rect 3141 22475 3207 22478
rect 13077 22475 13143 22478
rect 13310 22478 16000 22538
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 13169 22266 13235 22269
rect 13310 22266 13370 22478
rect 15520 22448 16000 22478
rect 13169 22264 13370 22266
rect 13169 22208 13174 22264
rect 13230 22208 13370 22264
rect 13169 22206 13370 22208
rect 13169 22203 13235 22206
rect 4521 22130 4587 22133
rect 8845 22130 8911 22133
rect 11513 22130 11579 22133
rect 4521 22128 11579 22130
rect 4521 22072 4526 22128
rect 4582 22072 8850 22128
rect 8906 22072 11518 22128
rect 11574 22072 11579 22128
rect 4521 22070 11579 22072
rect 4521 22067 4587 22070
rect 8845 22067 8911 22070
rect 11513 22067 11579 22070
rect 7189 21994 7255 21997
rect 9673 21994 9739 21997
rect 7189 21992 9739 21994
rect 7189 21936 7194 21992
rect 7250 21936 9678 21992
rect 9734 21936 9739 21992
rect 7189 21934 9739 21936
rect 7189 21931 7255 21934
rect 9673 21931 9739 21934
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 7281 20906 7347 20909
rect 10225 20906 10291 20909
rect 7281 20904 10291 20906
rect 7281 20848 7286 20904
rect 7342 20848 10230 20904
rect 10286 20848 10291 20904
rect 7281 20846 10291 20848
rect 7281 20843 7347 20846
rect 10225 20843 10291 20846
rect 10869 20770 10935 20773
rect 12525 20770 12591 20773
rect 10869 20768 12591 20770
rect 10869 20712 10874 20768
rect 10930 20712 12530 20768
rect 12586 20712 12591 20768
rect 10869 20710 12591 20712
rect 10869 20707 10935 20710
rect 12525 20707 12591 20710
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 4705 20362 4771 20365
rect 12525 20362 12591 20365
rect 4705 20360 12591 20362
rect 4705 20304 4710 20360
rect 4766 20304 12530 20360
rect 12586 20304 12591 20360
rect 4705 20302 12591 20304
rect 4705 20299 4771 20302
rect 12525 20299 12591 20302
rect 8661 20228 8727 20229
rect 8661 20226 8708 20228
rect 8616 20224 8708 20226
rect 8616 20168 8666 20224
rect 8616 20166 8708 20168
rect 8661 20164 8708 20166
rect 8772 20164 8778 20228
rect 8661 20163 8727 20164
rect 6277 20160 6597 20161
rect 0 20090 480 20120
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 2865 20090 2931 20093
rect 0 20088 2931 20090
rect 0 20032 2870 20088
rect 2926 20032 2931 20088
rect 0 20030 2931 20032
rect 0 20000 480 20030
rect 2865 20027 2931 20030
rect 4981 19818 5047 19821
rect 8753 19818 8819 19821
rect 4981 19816 8819 19818
rect 4981 19760 4986 19816
rect 5042 19760 8758 19816
rect 8814 19760 8819 19816
rect 4981 19758 8819 19760
rect 4981 19755 5047 19758
rect 8753 19755 8819 19758
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 8017 19138 8083 19141
rect 9765 19138 9831 19141
rect 8017 19136 9831 19138
rect 8017 19080 8022 19136
rect 8078 19080 9770 19136
rect 9826 19080 9831 19136
rect 8017 19078 9831 19080
rect 8017 19075 8083 19078
rect 9765 19075 9831 19078
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 11053 19002 11119 19005
rect 6686 19000 11119 19002
rect 6686 18944 11058 19000
rect 11114 18944 11119 19000
rect 6686 18942 11119 18944
rect 3969 18866 4035 18869
rect 6686 18866 6746 18942
rect 11053 18939 11119 18942
rect 3969 18864 6746 18866
rect 3969 18808 3974 18864
rect 4030 18808 6746 18864
rect 3969 18806 6746 18808
rect 7557 18866 7623 18869
rect 10685 18866 10751 18869
rect 7557 18864 10751 18866
rect 7557 18808 7562 18864
rect 7618 18808 10690 18864
rect 10746 18808 10751 18864
rect 7557 18806 10751 18808
rect 3969 18803 4035 18806
rect 7557 18803 7623 18806
rect 10685 18803 10751 18806
rect 2865 18730 2931 18733
rect 8293 18730 8359 18733
rect 2865 18728 8359 18730
rect 2865 18672 2870 18728
rect 2926 18672 8298 18728
rect 8354 18672 8359 18728
rect 2865 18670 8359 18672
rect 2865 18667 2931 18670
rect 8293 18667 8359 18670
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 5993 18458 6059 18461
rect 8753 18458 8819 18461
rect 5993 18456 8819 18458
rect 5993 18400 5998 18456
rect 6054 18400 8758 18456
rect 8814 18400 8819 18456
rect 5993 18398 8819 18400
rect 5993 18395 6059 18398
rect 8753 18395 8819 18398
rect 7189 18322 7255 18325
rect 10869 18322 10935 18325
rect 7189 18320 10935 18322
rect 7189 18264 7194 18320
rect 7250 18264 10874 18320
rect 10930 18264 10935 18320
rect 7189 18262 10935 18264
rect 7189 18259 7255 18262
rect 10869 18259 10935 18262
rect 4337 18186 4403 18189
rect 8518 18186 8524 18188
rect 4337 18184 8524 18186
rect 4337 18128 4342 18184
rect 4398 18128 8524 18184
rect 4337 18126 8524 18128
rect 4337 18123 4403 18126
rect 8518 18124 8524 18126
rect 8588 18186 8594 18188
rect 11145 18186 11211 18189
rect 8588 18184 11211 18186
rect 8588 18128 11150 18184
rect 11206 18128 11211 18184
rect 8588 18126 11211 18128
rect 8588 18124 8594 18126
rect 11145 18123 11211 18126
rect 8569 18050 8635 18053
rect 11145 18050 11211 18053
rect 8569 18048 11211 18050
rect 8569 17992 8574 18048
rect 8630 17992 11150 18048
rect 11206 17992 11211 18048
rect 8569 17990 11211 17992
rect 8569 17987 8635 17990
rect 11145 17987 11211 17990
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 3141 17778 3207 17781
rect 9305 17778 9371 17781
rect 3141 17776 9371 17778
rect 3141 17720 3146 17776
rect 3202 17720 9310 17776
rect 9366 17720 9371 17776
rect 3141 17718 9371 17720
rect 3141 17715 3207 17718
rect 9305 17715 9371 17718
rect 15520 17506 16000 17536
rect 14782 17446 16000 17506
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 4245 17370 4311 17373
rect 7833 17370 7899 17373
rect 4245 17368 7899 17370
rect 4245 17312 4250 17368
rect 4306 17312 7838 17368
rect 7894 17312 7899 17368
rect 4245 17310 7899 17312
rect 4245 17307 4311 17310
rect 7833 17307 7899 17310
rect 12709 17234 12775 17237
rect 14782 17234 14842 17446
rect 15520 17416 16000 17446
rect 12709 17232 14842 17234
rect 12709 17176 12714 17232
rect 12770 17176 14842 17232
rect 12709 17174 14842 17176
rect 12709 17171 12775 17174
rect 5809 17098 5875 17101
rect 7097 17098 7163 17101
rect 5809 17096 7163 17098
rect 5809 17040 5814 17096
rect 5870 17040 7102 17096
rect 7158 17040 7163 17096
rect 5809 17038 7163 17040
rect 5809 17035 5875 17038
rect 7097 17035 7163 17038
rect 8702 16900 8708 16964
rect 8772 16962 8778 16964
rect 8845 16962 8911 16965
rect 8772 16960 8911 16962
rect 8772 16904 8850 16960
rect 8906 16904 8911 16960
rect 8772 16902 8911 16904
rect 8772 16900 8778 16902
rect 8845 16899 8911 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 6821 16826 6887 16829
rect 9765 16826 9831 16829
rect 6821 16824 9831 16826
rect 6821 16768 6826 16824
rect 6882 16768 9770 16824
rect 9826 16768 9831 16824
rect 6821 16766 9831 16768
rect 6821 16763 6887 16766
rect 9765 16763 9831 16766
rect 5441 16690 5507 16693
rect 8845 16690 8911 16693
rect 5441 16688 8911 16690
rect 5441 16632 5446 16688
rect 5502 16632 8850 16688
rect 8906 16632 8911 16688
rect 5441 16630 8911 16632
rect 5441 16627 5507 16630
rect 8845 16627 8911 16630
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 8661 16146 8727 16149
rect 10869 16146 10935 16149
rect 8661 16144 10935 16146
rect 8661 16088 8666 16144
rect 8722 16088 10874 16144
rect 10930 16088 10935 16144
rect 8661 16086 10935 16088
rect 8661 16083 8727 16086
rect 10869 16083 10935 16086
rect 2865 16010 2931 16013
rect 8661 16010 8727 16013
rect 2865 16008 8727 16010
rect 2865 15952 2870 16008
rect 2926 15952 8666 16008
rect 8722 15952 8727 16008
rect 2865 15950 8727 15952
rect 2865 15947 2931 15950
rect 8661 15947 8727 15950
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 6637 15602 6703 15605
rect 8477 15602 8543 15605
rect 6637 15600 8543 15602
rect 6637 15544 6642 15600
rect 6698 15544 8482 15600
rect 8538 15544 8543 15600
rect 6637 15542 8543 15544
rect 6637 15539 6703 15542
rect 8477 15539 8543 15542
rect 3969 15466 4035 15469
rect 6637 15466 6703 15469
rect 3969 15464 6703 15466
rect 3969 15408 3974 15464
rect 4030 15408 6642 15464
rect 6698 15408 6703 15464
rect 3969 15406 6703 15408
rect 3969 15403 4035 15406
rect 6637 15403 6703 15406
rect 5257 15330 5323 15333
rect 7833 15330 7899 15333
rect 5257 15328 7899 15330
rect 5257 15272 5262 15328
rect 5318 15272 7838 15328
rect 7894 15272 7899 15328
rect 5257 15270 7899 15272
rect 5257 15267 5323 15270
rect 7833 15267 7899 15270
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 3417 15058 3483 15061
rect 12709 15058 12775 15061
rect 3417 15056 12775 15058
rect 3417 15000 3422 15056
rect 3478 15000 12714 15056
rect 12770 15000 12775 15056
rect 3417 14998 12775 15000
rect 3417 14995 3483 14998
rect 12709 14995 12775 14998
rect 5073 14922 5139 14925
rect 9857 14922 9923 14925
rect 5073 14920 9923 14922
rect 5073 14864 5078 14920
rect 5134 14864 9862 14920
rect 9918 14864 9923 14920
rect 5073 14862 9923 14864
rect 5073 14859 5139 14862
rect 9857 14859 9923 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 4429 14514 4495 14517
rect 8017 14514 8083 14517
rect 13445 14514 13511 14517
rect 4429 14512 13511 14514
rect 4429 14456 4434 14512
rect 4490 14456 8022 14512
rect 8078 14456 13450 14512
rect 13506 14456 13511 14512
rect 4429 14454 13511 14456
rect 4429 14451 4495 14454
rect 8017 14451 8083 14454
rect 13445 14451 13511 14454
rect 4061 14378 4127 14381
rect 6453 14378 6519 14381
rect 4061 14376 6519 14378
rect 4061 14320 4066 14376
rect 4122 14320 6458 14376
rect 6514 14320 6519 14376
rect 4061 14318 6519 14320
rect 4061 14315 4127 14318
rect 6453 14315 6519 14318
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 4061 13834 4127 13837
rect 6913 13834 6979 13837
rect 4061 13832 6979 13834
rect 4061 13776 4066 13832
rect 4122 13776 6918 13832
rect 6974 13776 6979 13832
rect 4061 13774 6979 13776
rect 4061 13771 4127 13774
rect 6913 13771 6979 13774
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 4429 13426 4495 13429
rect 8385 13426 8451 13429
rect 4429 13424 8451 13426
rect 4429 13368 4434 13424
rect 4490 13368 8390 13424
rect 8446 13368 8451 13424
rect 4429 13366 8451 13368
rect 4429 13363 4495 13366
rect 8385 13363 8451 13366
rect 8569 13426 8635 13429
rect 11145 13426 11211 13429
rect 8569 13424 11211 13426
rect 8569 13368 8574 13424
rect 8630 13368 11150 13424
rect 11206 13368 11211 13424
rect 8569 13366 11211 13368
rect 8569 13363 8635 13366
rect 11145 13363 11211 13366
rect 5073 13290 5139 13293
rect 10869 13290 10935 13293
rect 13353 13290 13419 13293
rect 5073 13288 13419 13290
rect 5073 13232 5078 13288
rect 5134 13232 10874 13288
rect 10930 13232 13358 13288
rect 13414 13232 13419 13288
rect 5073 13230 13419 13232
rect 5073 13227 5139 13230
rect 10869 13227 10935 13230
rect 13353 13227 13419 13230
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 8385 12746 8451 12749
rect 11145 12746 11211 12749
rect 8385 12744 11211 12746
rect 8385 12688 8390 12744
rect 8446 12688 11150 12744
rect 11206 12688 11211 12744
rect 8385 12686 11211 12688
rect 8385 12683 8451 12686
rect 11145 12683 11211 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 12065 12474 12131 12477
rect 15520 12474 16000 12504
rect 12065 12472 16000 12474
rect 12065 12416 12070 12472
rect 12126 12416 16000 12472
rect 12065 12414 16000 12416
rect 12065 12411 12131 12414
rect 15520 12384 16000 12414
rect 9438 12276 9444 12340
rect 9508 12338 9514 12340
rect 12801 12338 12867 12341
rect 9508 12336 12867 12338
rect 9508 12280 12806 12336
rect 12862 12280 12867 12336
rect 9508 12278 12867 12280
rect 9508 12276 9514 12278
rect 12801 12275 12867 12278
rect 8569 12204 8635 12205
rect 8518 12140 8524 12204
rect 8588 12202 8635 12204
rect 8588 12200 8680 12202
rect 8630 12144 8680 12200
rect 8588 12142 8680 12144
rect 8588 12140 8635 12142
rect 8569 12139 8635 12140
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 5073 11794 5139 11797
rect 11237 11794 11303 11797
rect 5073 11792 11303 11794
rect 5073 11736 5078 11792
rect 5134 11736 11242 11792
rect 11298 11736 11303 11792
rect 5073 11734 11303 11736
rect 5073 11731 5139 11734
rect 11237 11731 11303 11734
rect 6085 11658 6151 11661
rect 13261 11658 13327 11661
rect 6085 11656 13327 11658
rect 6085 11600 6090 11656
rect 6146 11600 13266 11656
rect 13322 11600 13327 11656
rect 6085 11598 13327 11600
rect 6085 11595 6151 11598
rect 13261 11595 13327 11598
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 8702 11188 8708 11252
rect 8772 11250 8778 11252
rect 9581 11250 9647 11253
rect 8772 11248 9647 11250
rect 8772 11192 9586 11248
rect 9642 11192 9647 11248
rect 8772 11190 9647 11192
rect 8772 11188 8778 11190
rect 9581 11187 9647 11190
rect 6545 11114 6611 11117
rect 8845 11114 8911 11117
rect 9857 11114 9923 11117
rect 6545 11112 9923 11114
rect 6545 11056 6550 11112
rect 6606 11056 8850 11112
rect 8906 11056 9862 11112
rect 9918 11056 9923 11112
rect 6545 11054 9923 11056
rect 6545 11051 6611 11054
rect 8845 11051 8911 11054
rect 9857 11051 9923 11054
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 9397 10842 9463 10845
rect 12433 10842 12499 10845
rect 9397 10840 12499 10842
rect 9397 10784 9402 10840
rect 9458 10784 12438 10840
rect 12494 10784 12499 10840
rect 9397 10782 12499 10784
rect 9397 10779 9463 10782
rect 12433 10779 12499 10782
rect 7741 10706 7807 10709
rect 11053 10706 11119 10709
rect 7741 10704 11119 10706
rect 7741 10648 7746 10704
rect 7802 10648 11058 10704
rect 11114 10648 11119 10704
rect 7741 10646 11119 10648
rect 7741 10643 7807 10646
rect 11053 10643 11119 10646
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 2957 10162 3023 10165
rect 4521 10162 4587 10165
rect 2957 10160 4587 10162
rect 2957 10104 2962 10160
rect 3018 10104 4526 10160
rect 4582 10104 4587 10160
rect 2957 10102 4587 10104
rect 2957 10099 3023 10102
rect 4521 10099 4587 10102
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 7189 9210 7255 9213
rect 8753 9210 8819 9213
rect 7189 9208 8819 9210
rect 7189 9152 7194 9208
rect 7250 9152 8758 9208
rect 8814 9152 8819 9208
rect 7189 9150 8819 9152
rect 7189 9147 7255 9150
rect 8753 9147 8819 9150
rect 7373 9074 7439 9077
rect 10685 9074 10751 9077
rect 7373 9072 10751 9074
rect 7373 9016 7378 9072
rect 7434 9016 10690 9072
rect 10746 9016 10751 9072
rect 7373 9014 10751 9016
rect 7373 9011 7439 9014
rect 10685 9011 10751 9014
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 5073 7986 5139 7989
rect 7005 7986 7071 7989
rect 5073 7984 7071 7986
rect 5073 7928 5078 7984
rect 5134 7928 7010 7984
rect 7066 7928 7071 7984
rect 5073 7926 7071 7928
rect 5073 7923 5139 7926
rect 7005 7923 7071 7926
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 5441 7442 5507 7445
rect 7189 7442 7255 7445
rect 5441 7440 7255 7442
rect 5441 7384 5446 7440
rect 5502 7384 7194 7440
rect 7250 7384 7255 7440
rect 5441 7382 7255 7384
rect 5441 7379 5507 7382
rect 7189 7379 7255 7382
rect 11697 7442 11763 7445
rect 15520 7442 16000 7472
rect 11697 7440 16000 7442
rect 11697 7384 11702 7440
rect 11758 7384 16000 7440
rect 11697 7382 16000 7384
rect 11697 7379 11763 7382
rect 15520 7352 16000 7382
rect 8845 7306 8911 7309
rect 11145 7306 11211 7309
rect 8845 7304 11211 7306
rect 8845 7248 8850 7304
rect 8906 7248 11150 7304
rect 11206 7248 11211 7304
rect 8845 7246 11211 7248
rect 8845 7243 8911 7246
rect 11145 7243 11211 7246
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 0 6762 480 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 480 6702
rect 4061 6699 4127 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 6269 5402 6335 5405
rect 7005 5402 7071 5405
rect 7649 5402 7715 5405
rect 6269 5400 7715 5402
rect 6269 5344 6274 5400
rect 6330 5344 7010 5400
rect 7066 5344 7654 5400
rect 7710 5344 7715 5400
rect 6269 5342 7715 5344
rect 6269 5339 6335 5342
rect 7005 5339 7071 5342
rect 7649 5339 7715 5342
rect 5165 5266 5231 5269
rect 11237 5266 11303 5269
rect 5165 5264 11303 5266
rect 5165 5208 5170 5264
rect 5226 5208 11242 5264
rect 11298 5208 11303 5264
rect 5165 5206 11303 5208
rect 5165 5203 5231 5206
rect 11237 5203 11303 5206
rect 5257 5130 5323 5133
rect 6729 5130 6795 5133
rect 5257 5128 6795 5130
rect 5257 5072 5262 5128
rect 5318 5072 6734 5128
rect 6790 5072 6795 5128
rect 5257 5070 6795 5072
rect 5257 5067 5323 5070
rect 6729 5067 6795 5070
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 8017 4586 8083 4589
rect 9673 4586 9739 4589
rect 8017 4584 9739 4586
rect 8017 4528 8022 4584
rect 8078 4528 9678 4584
rect 9734 4528 9739 4584
rect 8017 4526 9739 4528
rect 8017 4523 8083 4526
rect 9673 4523 9739 4526
rect 10777 4450 10843 4453
rect 13261 4450 13327 4453
rect 10777 4448 13327 4450
rect 10777 4392 10782 4448
rect 10838 4392 13266 4448
rect 13322 4392 13327 4448
rect 10777 4390 13327 4392
rect 10777 4387 10843 4390
rect 13261 4387 13327 4390
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 4613 4314 4679 4317
rect 8477 4314 8543 4317
rect 4613 4312 8543 4314
rect 4613 4256 4618 4312
rect 4674 4256 8482 4312
rect 8538 4256 8543 4312
rect 4613 4254 8543 4256
rect 4613 4251 4679 4254
rect 8477 4251 8543 4254
rect 6085 4178 6151 4181
rect 10225 4178 10291 4181
rect 6085 4176 10291 4178
rect 6085 4120 6090 4176
rect 6146 4120 10230 4176
rect 10286 4120 10291 4176
rect 6085 4118 10291 4120
rect 6085 4115 6151 4118
rect 10225 4115 10291 4118
rect 5390 3980 5396 4044
rect 5460 4042 5466 4044
rect 9438 4042 9444 4044
rect 5460 3982 9444 4042
rect 5460 3980 5466 3982
rect 9438 3980 9444 3982
rect 9508 3980 9514 4044
rect 11145 4042 11211 4045
rect 13537 4042 13603 4045
rect 9630 4040 13603 4042
rect 9630 3984 11150 4040
rect 11206 3984 13542 4040
rect 13598 3984 13603 4040
rect 9630 3982 13603 3984
rect 8661 3906 8727 3909
rect 9630 3906 9690 3982
rect 11145 3979 11211 3982
rect 13537 3979 13603 3982
rect 8661 3904 9690 3906
rect 8661 3848 8666 3904
rect 8722 3848 9690 3904
rect 8661 3846 9690 3848
rect 8661 3843 8727 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 7281 3770 7347 3773
rect 9581 3770 9647 3773
rect 7281 3768 10058 3770
rect 7281 3712 7286 3768
rect 7342 3712 9586 3768
rect 9642 3712 10058 3768
rect 7281 3710 10058 3712
rect 7281 3707 7347 3710
rect 9581 3707 9647 3710
rect 7833 3634 7899 3637
rect 9765 3634 9831 3637
rect 7833 3632 9831 3634
rect 7833 3576 7838 3632
rect 7894 3576 9770 3632
rect 9826 3576 9831 3632
rect 7833 3574 9831 3576
rect 9998 3634 10058 3710
rect 13537 3634 13603 3637
rect 9998 3632 13603 3634
rect 9998 3576 13542 3632
rect 13598 3576 13603 3632
rect 9998 3574 13603 3576
rect 7833 3571 7899 3574
rect 9765 3571 9831 3574
rect 13537 3571 13603 3574
rect 6085 3498 6151 3501
rect 12525 3498 12591 3501
rect 6085 3496 12591 3498
rect 6085 3440 6090 3496
rect 6146 3440 12530 3496
rect 12586 3440 12591 3496
rect 6085 3438 12591 3440
rect 6085 3435 6151 3438
rect 12525 3435 12591 3438
rect 5441 3362 5507 3365
rect 6913 3362 6979 3365
rect 7465 3362 7531 3365
rect 5441 3360 7531 3362
rect 5441 3304 5446 3360
rect 5502 3304 6918 3360
rect 6974 3304 7470 3360
rect 7526 3304 7531 3360
rect 5441 3302 7531 3304
rect 5441 3299 5507 3302
rect 6913 3299 6979 3302
rect 7465 3299 7531 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 4981 3226 5047 3229
rect 8661 3226 8727 3229
rect 4981 3224 8727 3226
rect 4981 3168 4986 3224
rect 5042 3168 8666 3224
rect 8722 3168 8727 3224
rect 4981 3166 8727 3168
rect 4981 3163 5047 3166
rect 8661 3163 8727 3166
rect 2037 3090 2103 3093
rect 12617 3090 12683 3093
rect 2037 3088 12683 3090
rect 2037 3032 2042 3088
rect 2098 3032 12622 3088
rect 12678 3032 12683 3088
rect 2037 3030 12683 3032
rect 2037 3027 2103 3030
rect 12617 3027 12683 3030
rect 3693 2954 3759 2957
rect 8293 2954 8359 2957
rect 3693 2952 8359 2954
rect 3693 2896 3698 2952
rect 3754 2896 8298 2952
rect 8354 2896 8359 2952
rect 3693 2894 8359 2896
rect 3693 2891 3759 2894
rect 8293 2891 8359 2894
rect 1209 2818 1275 2821
rect 4245 2818 4311 2821
rect 1209 2816 4311 2818
rect 1209 2760 1214 2816
rect 1270 2760 4250 2816
rect 4306 2760 4311 2816
rect 1209 2758 4311 2760
rect 1209 2755 1275 2758
rect 4245 2755 4311 2758
rect 5349 2820 5415 2821
rect 5349 2816 5396 2820
rect 5460 2818 5466 2820
rect 13629 2818 13695 2821
rect 15469 2818 15535 2821
rect 5349 2760 5354 2816
rect 5349 2756 5396 2760
rect 5460 2758 5506 2818
rect 13629 2816 15535 2818
rect 13629 2760 13634 2816
rect 13690 2760 15474 2816
rect 15530 2760 15535 2816
rect 13629 2758 15535 2760
rect 5460 2756 5466 2758
rect 5349 2755 5415 2756
rect 13629 2755 13695 2758
rect 15469 2755 15535 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 3509 2546 3575 2549
rect 7097 2546 7163 2549
rect 3509 2544 7163 2546
rect 3509 2488 3514 2544
rect 3570 2488 7102 2544
rect 7158 2488 7163 2544
rect 3509 2486 7163 2488
rect 3509 2483 3575 2486
rect 7097 2483 7163 2486
rect 8293 2546 8359 2549
rect 11237 2546 11303 2549
rect 8293 2544 11303 2546
rect 8293 2488 8298 2544
rect 8354 2488 11242 2544
rect 11298 2488 11303 2544
rect 8293 2486 11303 2488
rect 8293 2483 8359 2486
rect 11237 2483 11303 2486
rect 12065 2546 12131 2549
rect 15520 2546 16000 2576
rect 12065 2544 16000 2546
rect 12065 2488 12070 2544
rect 12126 2488 16000 2544
rect 12065 2486 16000 2488
rect 12065 2483 12131 2486
rect 15520 2456 16000 2486
rect 5901 2410 5967 2413
rect 7925 2410 7991 2413
rect 9857 2410 9923 2413
rect 5901 2408 7991 2410
rect 5901 2352 5906 2408
rect 5962 2352 7930 2408
rect 7986 2352 7991 2408
rect 5901 2350 7991 2352
rect 5901 2347 5967 2350
rect 7925 2347 7991 2350
rect 8710 2408 9923 2410
rect 8710 2352 9862 2408
rect 9918 2352 9923 2408
rect 8710 2350 9923 2352
rect 5073 2274 5139 2277
rect 8710 2274 8770 2350
rect 9857 2347 9923 2350
rect 5073 2272 8770 2274
rect 5073 2216 5078 2272
rect 5134 2216 8770 2272
rect 5073 2214 8770 2216
rect 5073 2211 5139 2214
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 5533 2138 5599 2141
rect 8569 2138 8635 2141
rect 5533 2136 8635 2138
rect 5533 2080 5538 2136
rect 5594 2080 8574 2136
rect 8630 2080 8635 2136
rect 5533 2078 8635 2080
rect 5533 2075 5599 2078
rect 8569 2075 8635 2078
rect 10409 1594 10475 1597
rect 12801 1594 12867 1597
rect 10409 1592 12867 1594
rect 10409 1536 10414 1592
rect 10470 1536 12806 1592
rect 12862 1536 12867 1592
rect 10409 1534 12867 1536
rect 10409 1531 10475 1534
rect 12801 1531 12867 1534
rect 9581 1458 9647 1461
rect 11513 1458 11579 1461
rect 9581 1456 11579 1458
rect 9581 1400 9586 1456
rect 9642 1400 11518 1456
rect 11574 1400 11579 1456
rect 9581 1398 11579 1400
rect 9581 1395 9647 1398
rect 11513 1395 11579 1398
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 9444 34852 9508 34916
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 8708 26480 8772 26484
rect 8708 26424 8758 26480
rect 8758 26424 8772 26480
rect 8708 26420 8772 26424
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 8708 20224 8772 20228
rect 8708 20168 8722 20224
rect 8722 20168 8772 20224
rect 8708 20164 8772 20168
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 8524 18124 8588 18188
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 8708 16900 8772 16964
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 9444 12276 9508 12340
rect 8524 12200 8588 12204
rect 8524 12144 8574 12200
rect 8574 12144 8588 12200
rect 8524 12140 8588 12144
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 8708 11188 8772 11252
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 5396 3980 5460 4044
rect 9444 3980 9508 4044
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 5396 2816 5460 2820
rect 5396 2760 5410 2816
rect 5410 2760 5460 2816
rect 5396 2756 5460 2760
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 9443 34916 9509 34917
rect 9443 34852 9444 34916
rect 9508 34852 9509 34916
rect 9443 34851 9509 34852
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8707 26484 8773 26485
rect 8707 26420 8708 26484
rect 8772 26420 8773 26484
rect 8707 26419 8773 26420
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 8710 20229 8770 26419
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8707 20228 8773 20229
rect 8707 20164 8708 20228
rect 8772 20164 8773 20228
rect 8707 20163 8773 20164
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8523 18188 8589 18189
rect 8523 18124 8524 18188
rect 8588 18124 8589 18188
rect 8523 18123 8589 18124
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 8526 12205 8586 18123
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8707 16964 8773 16965
rect 8707 16900 8708 16964
rect 8772 16900 8773 16964
rect 8707 16899 8773 16900
rect 8523 12204 8589 12205
rect 8523 12140 8524 12204
rect 8588 12140 8589 12204
rect 8523 12139 8589 12140
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 8710 11253 8770 16899
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 9446 12341 9506 34851
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 9443 12340 9509 12341
rect 9443 12276 9444 12340
rect 9508 12276 9509 12340
rect 9443 12275 9509 12276
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8707 11252 8773 11253
rect 8707 11188 8708 11252
rect 8772 11188 8773 11252
rect 8707 11187 8773 11188
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 5395 4044 5461 4045
rect 5395 3980 5396 4044
rect 5460 3980 5461 4044
rect 5395 3979 5461 3980
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 5398 2821 5458 3979
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 5395 2820 5461 2821
rect 5395 2756 5396 2820
rect 5460 2756 5461 2820
rect 5395 2755 5461 2756
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 9446 4045 9506 12275
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 9443 4044 9509 4045
rect 9443 3980 9444 4044
rect 9508 3980 9509 4044
rect 9443 3979 9509 3980
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_3_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_21 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_25 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _073_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_73
timestamp 1586364061
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_77
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _200_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_109
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_115
timestamp 1586364061
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _178_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_48
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_67
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_138 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_73
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_80
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_97
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_126
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_70
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_47
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_85
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _181_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_90
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_76
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 774 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_41
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_93
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_106
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_145
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_38
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_48
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_136
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_42
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_46
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_87
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_69
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_42
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_68
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_113
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_33
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_37
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_76
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_107
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_111
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_115
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_139
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_49
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_109
timestamp 1586364061
transform 1 0 11132 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_38
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_100
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_137
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_141
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_38
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_24_55
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_72
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 774 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 866 592
use scs8hd_decap_4  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_31
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 4692 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_46
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_42
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_48
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_52
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_65
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_102
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_115
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_111
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_decap_12  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_140
timestamp 1586364061
transform 1 0 13984 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_144
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_38
timestamp 1586364061
transform 1 0 4600 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_58
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_62
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_66
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_buf_1  _081_
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_41
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_106
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_or3_4  _069_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_48
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_52
timestamp 1586364061
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_65
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_4  FILLER_30_96
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 406 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_118
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_26
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 130 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_or3_4  _098_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_or3_4  _080_
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__C
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_19
timestamp 1586364061
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_8  _067_
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_43
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_47
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 406 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_60
timestamp 1586364061
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_77
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_81
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_85
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_32_98
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_109
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 774 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_120
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_132
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_144
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 3312 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_8  _159_
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_44
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_57
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_67
timestamp 1586364061
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_71
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_104
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_108
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_113
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_121
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_130
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_126
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_137
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_132
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_141
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_145
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_144
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_22
timestamp 1586364061
transform 1 0 3128 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_30
timestamp 1586364061
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_66
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_70
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_83
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_103
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_132
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_136
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_35_140
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_18
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_38
timestamp 1586364061
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_36_53
timestamp 1586364061
transform 1 0 5980 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_1  _093_
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_58
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_65
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_69
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_104
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 2300 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3312 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_16
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_20
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4876 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_33
timestamp 1586364061
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_37
timestamp 1586364061
transform 1 0 4508 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 6072 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_52
timestamp 1586364061
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_56
timestamp 1586364061
transform 1 0 6256 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_60
timestamp 1586364061
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_77
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_81
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8832 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_97
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_102
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 11868 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_137
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_141
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_145
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_or2_4  _171_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2576 0 -1 23392
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 4784 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_35
timestamp 1586364061
transform 1 0 4324 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_39
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 130 592
use scs8hd_nor3_4  _155_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 23392
box -38 -48 1234 592
use scs8hd_decap_3  FILLER_38_42
timestamp 1586364061
transform 1 0 4968 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_58
timestamp 1586364061
transform 1 0 6440 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_63
timestamp 1586364061
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_67
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_97
timestamp 1586364061
transform 1 0 10028 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_109
timestamp 1586364061
transform 1 0 11132 0 -1 23392
box -38 -48 774 592
use scs8hd_or2_4  _077_
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 682 592
use scs8hd_fill_2  FILLER_38_124
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_128
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _120_
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 866 592
use scs8hd_nor3_4  _156_
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 1234 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 4140 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__C
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_32
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_1  _076_
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 6164 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_42
timestamp 1586364061
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_46
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_53
timestamp 1586364061
transform 1 0 5980 0 -1 24480
box -38 -48 222 592
use scs8hd_or3_4  _119_
timestamp 1586364061
transform 1 0 6716 0 -1 24480
box -38 -48 866 592
use scs8hd_or4_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 6532 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_57
timestamp 1586364061
transform 1 0 6348 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_74
timestamp 1586364061
transform 1 0 7912 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_70
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 7728 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 8096 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_81
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_78
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 314 592
use scs8hd_or4_4  _147_
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__D
timestamp 1586364061
transform 1 0 9108 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_91
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_95
timestamp 1586364061
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_85
timestamp 1586364061
transform 1 0 8924 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_89
timestamp 1586364061
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 11224 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_99
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_119
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_144
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_36
timestamp 1586364061
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_or4_4  _095_
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_53
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_or4_4  _137_
timestamp 1586364061
transform 1 0 6992 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_73
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_77
timestamp 1586364061
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_81
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_97
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_101
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 774 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__D
timestamp 1586364061
transform 1 0 4692 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 4324 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_37
timestamp 1586364061
transform 1 0 4508 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_41
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 222 592
use scs8hd_nor3_4  _157_
timestamp 1586364061
transform 1 0 5244 0 -1 25568
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 5060 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 7176 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_58
timestamp 1586364061
transform 1 0 6440 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_62
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 8188 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_79
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_88
timestamp 1586364061
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_104
timestamp 1586364061
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_108
timestamp 1586364061
transform 1 0 11040 0 -1 25568
box -38 -48 406 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_115
timestamp 1586364061
transform 1 0 11684 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_119
timestamp 1586364061
transform 1 0 12052 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_131
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_42_143
timestamp 1586364061
transform 1 0 14260 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4784 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 4416 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_35
timestamp 1586364061
transform 1 0 4324 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_38
timestamp 1586364061
transform 1 0 4600 0 1 25568
box -38 -48 222 592
use scs8hd_or2_4  _129_
timestamp 1586364061
transform 1 0 5336 0 1 25568
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 5152 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_42
timestamp 1586364061
transform 1 0 4968 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_53
timestamp 1586364061
transform 1 0 5980 0 1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 774 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 7728 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 7544 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 8740 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_81
timestamp 1586364061
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_85
timestamp 1586364061
transform 1 0 8924 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_100
timestamp 1586364061
transform 1 0 10304 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_104
timestamp 1586364061
transform 1 0 10672 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_108
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_114
timestamp 1586364061
transform 1 0 11592 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_118
timestamp 1586364061
transform 1 0 11960 0 1 25568
box -38 -48 130 592
use scs8hd_fill_1  FILLER_43_121
timestamp 1586364061
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 4784 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 5796 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_49
timestamp 1586364061
transform 1 0 5612 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_53
timestamp 1586364061
transform 1 0 5980 0 -1 26656
box -38 -48 406 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 6348 0 -1 26656
box -38 -48 866 592
use scs8hd_decap_6  FILLER_44_66
timestamp 1586364061
transform 1 0 7176 0 -1 26656
box -38 -48 590 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 8004 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7728 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_74
timestamp 1586364061
transform 1 0 7912 0 -1 26656
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_84
timestamp 1586364061
transform 1 0 8832 0 -1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_44_88
timestamp 1586364061
transform 1 0 9200 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_44_91
timestamp 1586364061
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_98
timestamp 1586364061
transform 1 0 10120 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_111
timestamp 1586364061
transform 1 0 11316 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_115
timestamp 1586364061
transform 1 0 11684 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_122
timestamp 1586364061
transform 1 0 12328 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_134
timestamp 1586364061
transform 1 0 13432 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 4784 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 4140 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_35
timestamp 1586364061
transform 1 0 4324 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_53
timestamp 1586364061
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 7360 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_65
timestamp 1586364061
transform 1 0 7084 0 1 26656
box -38 -48 314 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 7728 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_70
timestamp 1586364061
transform 1 0 7544 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_83
timestamp 1586364061
transform 1 0 8740 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 8924 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 9292 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_87
timestamp 1586364061
transform 1 0 9108 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_91
timestamp 1586364061
transform 1 0 9476 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_95
timestamp 1586364061
transform 1 0 9844 0 1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 26656
box -38 -48 866 592
use scs8hd_decap_3  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_115
timestamp 1586364061
transform 1 0 11684 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_119
timestamp 1586364061
transform 1 0 12052 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_126
timestamp 1586364061
transform 1 0 12696 0 1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_45_132
timestamp 1586364061
transform 1 0 13248 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_144
timestamp 1586364061
transform 1 0 14352 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_nand2_4  _109_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 3220 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 3404 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_23
timestamp 1586364061
transform 1 0 3220 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_8  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_34
timestamp 1586364061
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 130 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 4140 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_38
timestamp 1586364061
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_36
timestamp 1586364061
transform 1 0 4416 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_40
timestamp 1586364061
transform 1 0 4784 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use scs8hd_nor3_4  _158_
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1234 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_53
timestamp 1586364061
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_57
timestamp 1586364061
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_61
timestamp 1586364061
transform 1 0 6716 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_57
timestamp 1586364061
transform 1 0 6348 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 6532 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 6900 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_65
timestamp 1586364061
transform 1 0 7084 0 -1 27744
box -38 -48 774 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 6900 0 1 27744
box -38 -48 866 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 7912 0 -1 27744
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_73
timestamp 1586364061
transform 1 0 7820 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_46_83
timestamp 1586364061
transform 1 0 8740 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_72
timestamp 1586364061
transform 1 0 7728 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_76
timestamp 1586364061
transform 1 0 8096 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 9660 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_87
timestamp 1586364061
transform 1 0 9108 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_91
timestamp 1586364061
transform 1 0 9476 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_95
timestamp 1586364061
transform 1 0 9844 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10212 0 1 27744
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_109
timestamp 1586364061
transform 1 0 11132 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_114
timestamp 1586364061
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_118
timestamp 1586364061
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_122
timestamp 1586364061
transform 1 0 12328 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 27744
box -38 -48 866 592
use scs8hd_or2_4  _072_
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 682 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 13248 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_126
timestamp 1586364061
transform 1 0 12696 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_133
timestamp 1586364061
transform 1 0 13340 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_130
timestamp 1586364061
transform 1 0 13064 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_134
timestamp 1586364061
transform 1 0 13432 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_47_138
timestamp 1586364061
transform 1 0 13800 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_8  _162_
timestamp 1586364061
transform 1 0 4692 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_36
timestamp 1586364061
transform 1 0 4416 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_48
timestamp 1586364061
transform 1 0 5520 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_52
timestamp 1586364061
transform 1 0 5888 0 -1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 7268 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_65
timestamp 1586364061
transform 1 0 7084 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_48_69
timestamp 1586364061
transform 1 0 7452 0 -1 28832
box -38 -48 590 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 8004 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_84
timestamp 1586364061
transform 1 0 8832 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 28832
box -38 -48 866 592
use scs8hd_fill_1  FILLER_48_97
timestamp 1586364061
transform 1 0 10028 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_107
timestamp 1586364061
transform 1 0 10948 0 -1 28832
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 28832
box -38 -48 866 592
use scs8hd_decap_8  FILLER_48_124
timestamp 1586364061
transform 1 0 12512 0 -1 28832
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_8  FILLER_48_135
timestamp 1586364061
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_143
timestamp 1586364061
transform 1 0 14260 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_19
timestamp 1586364061
transform 1 0 2852 0 1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_49_22
timestamp 1586364061
transform 1 0 3128 0 1 28832
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_33
timestamp 1586364061
transform 1 0 4140 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_37
timestamp 1586364061
transform 1 0 4508 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_50
timestamp 1586364061
transform 1 0 5704 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_54
timestamp 1586364061
transform 1 0 6072 0 1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8556 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_71
timestamp 1586364061
transform 1 0 7636 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_77
timestamp 1586364061
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_92
timestamp 1586364061
transform 1 0 9568 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_96
timestamp 1586364061
transform 1 0 9936 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_109
timestamp 1586364061
transform 1 0 11132 0 1 28832
box -38 -48 1142 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_fill_1  FILLER_49_121
timestamp 1586364061
transform 1 0 12236 0 1 28832
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 13248 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_126
timestamp 1586364061
transform 1 0 12696 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_130
timestamp 1586364061
transform 1 0 13064 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_137
timestamp 1586364061
transform 1 0 13708 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_141
timestamp 1586364061
transform 1 0 14076 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_145
timestamp 1586364061
transform 1 0 14444 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_19
timestamp 1586364061
transform 1 0 2852 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_23
timestamp 1586364061
transform 1 0 3220 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_36
timestamp 1586364061
transform 1 0 4416 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_48
timestamp 1586364061
transform 1 0 5520 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_52
timestamp 1586364061
transform 1 0 5888 0 -1 29920
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_58
timestamp 1586364061
transform 1 0 6440 0 -1 29920
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 8372 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_71
timestamp 1586364061
transform 1 0 7636 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_75
timestamp 1586364061
transform 1 0 8004 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_8  FILLER_50_82
timestamp 1586364061
transform 1 0 8648 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 29920
box -38 -48 222 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 11224 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_102
timestamp 1586364061
transform 1 0 10488 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_106
timestamp 1586364061
transform 1 0 10856 0 -1 29920
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_8  FILLER_50_113
timestamp 1586364061
transform 1 0 11500 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_12  FILLER_50_124
timestamp 1586364061
transform 1 0 12512 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_136
timestamp 1586364061
transform 1 0 13616 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_144
timestamp 1586364061
transform 1 0 14352 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 222 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 3956 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_34
timestamp 1586364061
transform 1 0 4232 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_40
timestamp 1586364061
transform 1 0 4784 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 29920
box -38 -48 866 592
use scs8hd_decap_4  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_55
timestamp 1586364061
transform 1 0 6164 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 6256 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_58
timestamp 1586364061
transform 1 0 6440 0 1 29920
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_73
timestamp 1586364061
transform 1 0 7820 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_77
timestamp 1586364061
transform 1 0 8188 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_81
timestamp 1586364061
transform 1 0 8556 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_85
timestamp 1586364061
transform 1 0 8924 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_89
timestamp 1586364061
transform 1 0 9292 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_104
timestamp 1586364061
transform 1 0 10672 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_108
timestamp 1586364061
transform 1 0 11040 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_114
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_118
timestamp 1586364061
transform 1 0 11960 0 1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 406 592
use scs8hd_inv_8  _161_
timestamp 1586364061
transform 1 0 4600 0 1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 4416 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_53_31
timestamp 1586364061
transform 1 0 3956 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_34
timestamp 1586364061
transform 1 0 4232 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 5612 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_47
timestamp 1586364061
transform 1 0 5428 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_51
timestamp 1586364061
transform 1 0 5796 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_55
timestamp 1586364061
transform 1 0 6164 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_47
timestamp 1586364061
transform 1 0 5428 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_55
timestamp 1586364061
transform 1 0 6164 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_66
timestamp 1586364061
transform 1 0 7176 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_52_67
timestamp 1586364061
transform 1 0 7268 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_63
timestamp 1586364061
transform 1 0 6900 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7084 0 -1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 31008
box -38 -48 866 592
use scs8hd_or2_4  _145_
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 682 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_78
timestamp 1586364061
transform 1 0 8280 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  FILLER_53_83
timestamp 1586364061
transform 1 0 8740 0 1 31008
box -38 -48 314 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 9016 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_84
timestamp 1586364061
transform 1 0 8832 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_88
timestamp 1586364061
transform 1 0 9200 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_95
timestamp 1586364061
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_104
timestamp 1586364061
transform 1 0 10672 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_108
timestamp 1586364061
transform 1 0 11040 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_99
timestamp 1586364061
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_103
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_121
timestamp 1586364061
transform 1 0 12236 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_113
timestamp 1586364061
transform 1 0 11500 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_117
timestamp 1586364061
transform 1 0 11868 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_121
timestamp 1586364061
transform 1 0 12236 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_133
timestamp 1586364061
transform 1 0 13340 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_35
timestamp 1586364061
transform 1 0 4324 0 -1 32096
box -38 -48 774 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 5244 0 -1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_54_43
timestamp 1586364061
transform 1 0 5060 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_54
timestamp 1586364061
transform 1 0 6072 0 -1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_58
timestamp 1586364061
transform 1 0 6440 0 -1 32096
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_71
timestamp 1586364061
transform 1 0 7636 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_75
timestamp 1586364061
transform 1 0 8004 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_79
timestamp 1586364061
transform 1 0 8372 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 9016 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_84
timestamp 1586364061
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_88
timestamp 1586364061
transform 1 0 9200 0 -1 32096
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_106
timestamp 1586364061
transform 1 0 10856 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_113
timestamp 1586364061
transform 1 0 11500 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_125
timestamp 1586364061
transform 1 0 12604 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_54_137
timestamp 1586364061
transform 1 0 13708 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_36
timestamp 1586364061
transform 1 0 4416 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_40
timestamp 1586364061
transform 1 0 4784 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7360 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_79
timestamp 1586364061
transform 1 0 8372 0 1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_55_83
timestamp 1586364061
transform 1 0 8740 0 1 32096
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_89
timestamp 1586364061
transform 1 0 9292 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_92
timestamp 1586364061
transform 1 0 9568 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_105
timestamp 1586364061
transform 1 0 10764 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_109
timestamp 1586364061
transform 1 0 11132 0 1 32096
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_113
timestamp 1586364061
transform 1 0 11500 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_117
timestamp 1586364061
transform 1 0 11868 0 1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_55_121
timestamp 1586364061
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_126
timestamp 1586364061
transform 1 0 12696 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_130
timestamp 1586364061
transform 1 0 13064 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_134
timestamp 1586364061
transform 1 0 13432 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_56_29
timestamp 1586364061
transform 1 0 3772 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_56_38
timestamp 1586364061
transform 1 0 4600 0 -1 33184
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 5520 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_42
timestamp 1586364061
transform 1 0 4968 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_46
timestamp 1586364061
transform 1 0 5336 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_61
timestamp 1586364061
transform 1 0 6716 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_65
timestamp 1586364061
transform 1 0 7084 0 -1 33184
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 33184
box -38 -48 866 592
use scs8hd_decap_3  FILLER_56_70
timestamp 1586364061
transform 1 0 7544 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_82
timestamp 1586364061
transform 1 0 8648 0 -1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_86
timestamp 1586364061
transform 1 0 9016 0 -1 33184
box -38 -48 590 592
use scs8hd_fill_2  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 33184
box -38 -48 866 592
use scs8hd_fill_1  FILLER_56_97
timestamp 1586364061
transform 1 0 10028 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_107
timestamp 1586364061
transform 1 0 10948 0 -1 33184
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_111
timestamp 1586364061
transform 1 0 11316 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_1  FILLER_56_114
timestamp 1586364061
transform 1 0 11592 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_124
timestamp 1586364061
transform 1 0 12512 0 -1 33184
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_135
timestamp 1586364061
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_143
timestamp 1586364061
transform 1 0 14260 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 3404 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_23
timestamp 1586364061
transform 1 0 3220 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_36
timestamp 1586364061
transform 1 0 4416 0 1 33184
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 5152 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_42
timestamp 1586364061
transform 1 0 4968 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_53
timestamp 1586364061
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8740 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_71
timestamp 1586364061
transform 1 0 7636 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_75
timestamp 1586364061
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_79
timestamp 1586364061
transform 1 0 8372 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_94
timestamp 1586364061
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_113
timestamp 1586364061
transform 1 0 11500 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_117
timestamp 1586364061
transform 1 0 11868 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_132
timestamp 1586364061
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_136
timestamp 1586364061
transform 1 0 13616 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_144
timestamp 1586364061
transform 1 0 14352 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 5244 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_43
timestamp 1586364061
transform 1 0 5060 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_47
timestamp 1586364061
transform 1 0 5428 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_62
timestamp 1586364061
transform 1 0 6808 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_66
timestamp 1586364061
transform 1 0 7176 0 -1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8648 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_79
timestamp 1586364061
transform 1 0 8372 0 -1 34272
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_84
timestamp 1586364061
transform 1 0 8832 0 -1 34272
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_104
timestamp 1586364061
transform 1 0 10672 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_108
timestamp 1586364061
transform 1 0 11040 0 -1 34272
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_121
timestamp 1586364061
transform 1 0 12236 0 -1 34272
box -38 -48 222 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 13340 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_58_125
timestamp 1586364061
transform 1 0 12604 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_8  FILLER_58_137
timestamp 1586364061
transform 1 0 13708 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 590 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_36
timestamp 1586364061
transform 1 0 4416 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_40
timestamp 1586364061
transform 1 0 4784 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 5152 0 1 34272
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 4968 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_53
timestamp 1586364061
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_46
timestamp 1586364061
transform 1 0 5336 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_50
timestamp 1586364061
transform 1 0 5704 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_6  FILLER_60_54
timestamp 1586364061
transform 1 0 6072 0 -1 35360
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_57
timestamp 1586364061
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8648 0 1 34272
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_73
timestamp 1586364061
transform 1 0 7820 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_78
timestamp 1586364061
transform 1 0 8280 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_71
timestamp 1586364061
transform 1 0 7636 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_60_75
timestamp 1586364061
transform 1 0 8004 0 -1 35360
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_93
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_84
timestamp 1586364061
transform 1 0 8832 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_1  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_97
timestamp 1586364061
transform 1 0 10028 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_110
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_103
timestamp 1586364061
transform 1 0 10580 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_60_107
timestamp 1586364061
transform 1 0 10948 0 -1 35360
box -38 -48 590 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 11500 0 -1 35360
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 11500 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_59_115
timestamp 1586364061
transform 1 0 11684 0 1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_59_121
timestamp 1586364061
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 13432 0 1 34272
box -38 -48 406 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 12696 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 13248 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_126
timestamp 1586364061
transform 1 0 12696 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_130
timestamp 1586364061
transform 1 0 13064 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_138
timestamp 1586364061
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_125
timestamp 1586364061
transform 1 0 12604 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_130
timestamp 1586364061
transform 1 0 13064 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_142
timestamp 1586364061
transform 1 0 14168 0 1 34272
box -38 -48 406 592
use scs8hd_decap_4  FILLER_60_142
timestamp 1586364061
transform 1 0 14168 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_57
timestamp 1586364061
transform 1 0 6348 0 1 35360
box -38 -48 222 592
use scs8hd_decap_3  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 8648 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 8464 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_78
timestamp 1586364061
transform 1 0 8280 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_91
timestamp 1586364061
transform 1 0 9476 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_95
timestamp 1586364061
transform 1 0 9844 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 10764 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_103
timestamp 1586364061
transform 1 0 10580 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_107
timestamp 1586364061
transform 1 0 10948 0 1 35360
box -38 -48 406 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 35360
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 11776 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_114
timestamp 1586364061
transform 1 0 11592 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_118
timestamp 1586364061
transform 1 0 11960 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 12972 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_127
timestamp 1586364061
transform 1 0 12788 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_131
timestamp 1586364061
transform 1 0 13156 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 36448
box -38 -48 866 592
use scs8hd_decap_8  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_62_64
timestamp 1586364061
transform 1 0 6992 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 8648 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_74
timestamp 1586364061
transform 1 0 7912 0 -1 36448
box -38 -48 774 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_84
timestamp 1586364061
transform 1 0 8832 0 -1 36448
box -38 -48 774 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 11224 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_97
timestamp 1586364061
transform 1 0 10028 0 -1 36448
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_62_109
timestamp 1586364061
transform 1 0 11132 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_114
timestamp 1586364061
transform 1 0 11592 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_126
timestamp 1586364061
transform 1 0 12696 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_62_138
timestamp 1586364061
transform 1 0 13800 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_66
timestamp 1586364061
transform 1 0 7176 0 1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 8004 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 7820 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_70
timestamp 1586364061
transform 1 0 7544 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_84
timestamp 1586364061
transform 1 0 8832 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_96
timestamp 1586364061
transform 1 0 9936 0 1 36448
box -38 -48 774 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 10764 0 1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_63_104
timestamp 1586364061
transform 1 0 10672 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_109
timestamp 1586364061
transform 1 0 11132 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 11316 0 1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_63_113
timestamp 1586364061
transform 1 0 11500 0 1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_63_121
timestamp 1586364061
transform 1 0 12236 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_64_77
timestamp 1586364061
transform 1 0 8188 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_89
timestamp 1586364061
transform 1 0 9292 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal2 s 5814 39520 5870 40000 6 address[0]
port 0 nsew default input
rlabel metal2 s 6366 39520 6422 40000 6 address[1]
port 1 nsew default input
rlabel metal2 s 7010 39520 7066 40000 6 address[2]
port 2 nsew default input
rlabel metal2 s 7654 39520 7710 40000 6 address[3]
port 3 nsew default input
rlabel metal2 s 8298 39520 8354 40000 6 address[4]
port 4 nsew default input
rlabel metal2 s 8850 39520 8906 40000 6 address[5]
port 5 nsew default input
rlabel metal2 s 9494 39520 9550 40000 6 address[6]
port 6 nsew default input
rlabel metal2 s 386 0 442 480 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 1214 0 1270 480 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 2042 0 2098 480 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 6274 0 6330 480 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal2 s 294 39520 350 40000 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 846 39520 902 40000 6 chany_top_in[1]
port 26 nsew default input
rlabel metal2 s 1490 39520 1546 40000 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_in[3]
port 28 nsew default input
rlabel metal2 s 2686 39520 2742 40000 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_in[5]
port 30 nsew default input
rlabel metal2 s 3974 39520 4030 40000 6 chany_top_in[6]
port 31 nsew default input
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_in[7]
port 32 nsew default input
rlabel metal2 s 5170 39520 5226 40000 6 chany_top_in[8]
port 33 nsew default input
rlabel metal2 s 10690 39520 10746 40000 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal2 s 11978 39520 12034 40000 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal2 s 13174 39520 13230 40000 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 13818 39520 13874 40000 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 14370 39520 14426 40000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal2 s 15014 39520 15070 40000 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal2 s 15658 39520 15714 40000 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal2 s 10138 39520 10194 40000 6 data_in
port 43 nsew default input
rlabel metal2 s 7930 0 7986 480 6 enable
port 44 nsew default input
rlabel metal3 s 0 6672 480 6792 6 left_grid_pin_1_
port 45 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 left_grid_pin_5_
port 46 nsew default tristate
rlabel metal3 s 0 33328 480 33448 6 left_grid_pin_9_
port 47 nsew default tristate
rlabel metal3 s 15520 2456 16000 2576 6 right_grid_pin_0_
port 48 nsew default tristate
rlabel metal3 s 15520 27344 16000 27464 6 right_grid_pin_10_
port 49 nsew default tristate
rlabel metal3 s 15520 32376 16000 32496 6 right_grid_pin_12_
port 50 nsew default tristate
rlabel metal3 s 15520 37408 16000 37528 6 right_grid_pin_14_
port 51 nsew default tristate
rlabel metal3 s 15520 7352 16000 7472 6 right_grid_pin_2_
port 52 nsew default tristate
rlabel metal3 s 15520 12384 16000 12504 6 right_grid_pin_4_
port 53 nsew default tristate
rlabel metal3 s 15520 17416 16000 17536 6 right_grid_pin_6_
port 54 nsew default tristate
rlabel metal3 s 15520 22448 16000 22568 6 right_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 56 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 57 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
