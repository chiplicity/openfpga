VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2223.700 BY 2027.600 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1364.040 51.880 1364.640 ;
    END
  END address[0]
  PIN address[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1710.840 2174.480 1711.440 ;
    END
  END address[10]
  PIN address[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1771.360 2174.480 1771.960 ;
    END
  END address[11]
  PIN address[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1471.480 51.880 1472.080 ;
    END
  END address[12]
  PIN address[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1525.200 51.880 1525.800 ;
    END
  END address[13]
  PIN address[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1842.190 1981.720 1842.470 1984.120 ;
    END
  END address[14]
  PIN address[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1579.600 51.880 1580.200 ;
    END
  END address[15]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1627.370 44.120 1627.650 46.520 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1528.600 2174.480 1529.200 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1691.770 44.120 1692.050 46.520 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.170 44.120 1756.450 46.520 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1709.710 1981.720 1709.990 1984.120 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1589.120 2174.480 1589.720 ;
    END
  END address[6]
  PIN address[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1417.760 51.880 1418.360 ;
    END
  END address[7]
  PIN address[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1650.320 2174.480 1650.920 ;
    END
  END address[8]
  PIN address[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1820.570 44.120 1820.850 46.520 ;
    END
  END address[9]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1975.130 1981.720 1975.410 1984.120 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1633.320 51.880 1633.920 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1884.970 44.120 1885.250 46.520 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 115.810 1981.720 116.090 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[10]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 647.110 1981.720 647.390 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[10]
  PIN gfpga_pad_GPIO_PAD[11]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 779.590 1981.720 779.870 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[11]
  PIN gfpga_pad_GPIO_PAD[12]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 912.530 1981.720 912.810 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[12]
  PIN gfpga_pad_GPIO_PAD[13]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1045.470 1981.720 1045.750 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[13]
  PIN gfpga_pad_GPIO_PAD[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1831.880 2174.480 1832.480 ;
    END
  END gfpga_pad_GPIO_PAD[14]
  PIN gfpga_pad_GPIO_PAD[15]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1902.600 51.880 1903.200 ;
    END
  END gfpga_pad_GPIO_PAD[15]
  PIN gfpga_pad_GPIO_PAD[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2108.070 1981.720 2108.350 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[16]
  PIN gfpga_pad_GPIO_PAD[17]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1892.400 2174.480 1893.000 ;
    END
  END gfpga_pad_GPIO_PAD[17]
  PIN gfpga_pad_GPIO_PAD[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2078.170 44.120 2078.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[18]
  PIN gfpga_pad_GPIO_PAD[19]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1952.920 2174.480 1953.520 ;
    END
  END gfpga_pad_GPIO_PAD[19]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 248.290 1981.720 248.570 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1178.410 1981.720 1178.690 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[20]
  PIN gfpga_pad_GPIO_PAD[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1310.890 1981.720 1311.170 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[21]
  PIN gfpga_pad_GPIO_PAD[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1443.830 1981.720 1444.110 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[22]
  PIN gfpga_pad_GPIO_PAD[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1576.770 1981.720 1577.050 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[23]
  PIN gfpga_pad_GPIO_PAD[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 74.080 2174.480 74.680 ;
    END
  END gfpga_pad_GPIO_PAD[24]
  PIN gfpga_pad_GPIO_PAD[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 134.600 2174.480 135.200 ;
    END
  END gfpga_pad_GPIO_PAD[25]
  PIN gfpga_pad_GPIO_PAD[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 195.120 2174.480 195.720 ;
    END
  END gfpga_pad_GPIO_PAD[26]
  PIN gfpga_pad_GPIO_PAD[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 255.640 2174.480 256.240 ;
    END
  END gfpga_pad_GPIO_PAD[27]
  PIN gfpga_pad_GPIO_PAD[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 316.160 2174.480 316.760 ;
    END
  END gfpga_pad_GPIO_PAD[28]
  PIN gfpga_pad_GPIO_PAD[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 376.680 2174.480 377.280 ;
    END
  END gfpga_pad_GPIO_PAD[29]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 381.230 1981.720 381.510 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 437.200 2174.480 437.800 ;
    END
  END gfpga_pad_GPIO_PAD[30]
  PIN gfpga_pad_GPIO_PAD[31]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 498.400 2174.480 499.000 ;
    END
  END gfpga_pad_GPIO_PAD[31]
  PIN gfpga_pad_GPIO_PAD[32]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 558.920 2174.480 559.520 ;
    END
  END gfpga_pad_GPIO_PAD[32]
  PIN gfpga_pad_GPIO_PAD[33]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 619.440 2174.480 620.040 ;
    END
  END gfpga_pad_GPIO_PAD[33]
  PIN gfpga_pad_GPIO_PAD[34]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 679.960 2174.480 680.560 ;
    END
  END gfpga_pad_GPIO_PAD[34]
  PIN gfpga_pad_GPIO_PAD[35]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 740.480 2174.480 741.080 ;
    END
  END gfpga_pad_GPIO_PAD[35]
  PIN gfpga_pad_GPIO_PAD[36]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 801.000 2174.480 801.600 ;
    END
  END gfpga_pad_GPIO_PAD[36]
  PIN gfpga_pad_GPIO_PAD[37]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 862.200 2174.480 862.800 ;
    END
  END gfpga_pad_GPIO_PAD[37]
  PIN gfpga_pad_GPIO_PAD[38]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 922.720 2174.480 923.320 ;
    END
  END gfpga_pad_GPIO_PAD[38]
  PIN gfpga_pad_GPIO_PAD[39]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 983.240 2174.480 983.840 ;
    END
  END gfpga_pad_GPIO_PAD[39]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 514.170 1981.720 514.450 1984.120 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[40]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1043.760 2174.480 1044.360 ;
    END
  END gfpga_pad_GPIO_PAD[40]
  PIN gfpga_pad_GPIO_PAD[41]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1104.280 2174.480 1104.880 ;
    END
  END gfpga_pad_GPIO_PAD[41]
  PIN gfpga_pad_GPIO_PAD[42]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1164.800 2174.480 1165.400 ;
    END
  END gfpga_pad_GPIO_PAD[42]
  PIN gfpga_pad_GPIO_PAD[43]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1225.320 2174.480 1225.920 ;
    END
  END gfpga_pad_GPIO_PAD[43]
  PIN gfpga_pad_GPIO_PAD[44]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1286.520 2174.480 1287.120 ;
    END
  END gfpga_pad_GPIO_PAD[44]
  PIN gfpga_pad_GPIO_PAD[45]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1347.040 2174.480 1347.640 ;
    END
  END gfpga_pad_GPIO_PAD[45]
  PIN gfpga_pad_GPIO_PAD[46]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1407.560 2174.480 1408.160 ;
    END
  END gfpga_pad_GPIO_PAD[46]
  PIN gfpga_pad_GPIO_PAD[47]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2172.080 1468.080 2174.480 1468.680 ;
    END
  END gfpga_pad_GPIO_PAD[47]
  PIN gfpga_pad_GPIO_PAD[48]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 81.770 44.120 82.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[48]
  PIN gfpga_pad_GPIO_PAD[49]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 146.170 44.120 146.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[49]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1687.040 51.880 1687.640 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[50]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 210.570 44.120 210.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[50]
  PIN gfpga_pad_GPIO_PAD[51]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 274.970 44.120 275.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[51]
  PIN gfpga_pad_GPIO_PAD[52]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 339.370 44.120 339.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[52]
  PIN gfpga_pad_GPIO_PAD[53]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 403.770 44.120 404.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[53]
  PIN gfpga_pad_GPIO_PAD[54]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 468.170 44.120 468.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[54]
  PIN gfpga_pad_GPIO_PAD[55]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 532.570 44.120 532.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[55]
  PIN gfpga_pad_GPIO_PAD[56]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 596.970 44.120 597.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[56]
  PIN gfpga_pad_GPIO_PAD[57]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 661.370 44.120 661.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[57]
  PIN gfpga_pad_GPIO_PAD[58]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 725.770 44.120 726.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[58]
  PIN gfpga_pad_GPIO_PAD[59]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 790.170 44.120 790.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[59]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1740.760 51.880 1741.360 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[60]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 854.570 44.120 854.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[60]
  PIN gfpga_pad_GPIO_PAD[61]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 918.970 44.120 919.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[61]
  PIN gfpga_pad_GPIO_PAD[62]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 983.370 44.120 983.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[62]
  PIN gfpga_pad_GPIO_PAD[63]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1047.770 44.120 1048.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[63]
  PIN gfpga_pad_GPIO_PAD[64]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1112.170 44.120 1112.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[64]
  PIN gfpga_pad_GPIO_PAD[65]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1176.570 44.120 1176.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[65]
  PIN gfpga_pad_GPIO_PAD[66]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1240.970 44.120 1241.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[66]
  PIN gfpga_pad_GPIO_PAD[67]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1305.370 44.120 1305.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[67]
  PIN gfpga_pad_GPIO_PAD[68]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1369.770 44.120 1370.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[68]
  PIN gfpga_pad_GPIO_PAD[69]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1434.170 44.120 1434.450 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[69]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1795.160 51.880 1795.760 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[70]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1498.570 44.120 1498.850 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[70]
  PIN gfpga_pad_GPIO_PAD[71]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1562.970 44.120 1563.250 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[71]
  PIN gfpga_pad_GPIO_PAD[72]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 70.680 51.880 71.280 ;
    END
  END gfpga_pad_GPIO_PAD[72]
  PIN gfpga_pad_GPIO_PAD[73]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 124.400 51.880 125.000 ;
    END
  END gfpga_pad_GPIO_PAD[73]
  PIN gfpga_pad_GPIO_PAD[74]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 178.120 51.880 178.720 ;
    END
  END gfpga_pad_GPIO_PAD[74]
  PIN gfpga_pad_GPIO_PAD[75]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 231.840 51.880 232.440 ;
    END
  END gfpga_pad_GPIO_PAD[75]
  PIN gfpga_pad_GPIO_PAD[76]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 286.240 51.880 286.840 ;
    END
  END gfpga_pad_GPIO_PAD[76]
  PIN gfpga_pad_GPIO_PAD[77]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 339.960 51.880 340.560 ;
    END
  END gfpga_pad_GPIO_PAD[77]
  PIN gfpga_pad_GPIO_PAD[78]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 393.680 51.880 394.280 ;
    END
  END gfpga_pad_GPIO_PAD[78]
  PIN gfpga_pad_GPIO_PAD[79]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 447.400 51.880 448.000 ;
    END
  END gfpga_pad_GPIO_PAD[79]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1949.370 44.120 1949.650 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN gfpga_pad_GPIO_PAD[80]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 501.800 51.880 502.400 ;
    END
  END gfpga_pad_GPIO_PAD[80]
  PIN gfpga_pad_GPIO_PAD[81]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 555.520 51.880 556.120 ;
    END
  END gfpga_pad_GPIO_PAD[81]
  PIN gfpga_pad_GPIO_PAD[82]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 609.240 51.880 609.840 ;
    END
  END gfpga_pad_GPIO_PAD[82]
  PIN gfpga_pad_GPIO_PAD[83]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 662.960 51.880 663.560 ;
    END
  END gfpga_pad_GPIO_PAD[83]
  PIN gfpga_pad_GPIO_PAD[84]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 717.360 51.880 717.960 ;
    END
  END gfpga_pad_GPIO_PAD[84]
  PIN gfpga_pad_GPIO_PAD[85]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 771.080 51.880 771.680 ;
    END
  END gfpga_pad_GPIO_PAD[85]
  PIN gfpga_pad_GPIO_PAD[86]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 824.800 51.880 825.400 ;
    END
  END gfpga_pad_GPIO_PAD[86]
  PIN gfpga_pad_GPIO_PAD[87]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 878.520 51.880 879.120 ;
    END
  END gfpga_pad_GPIO_PAD[87]
  PIN gfpga_pad_GPIO_PAD[88]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 932.920 51.880 933.520 ;
    END
  END gfpga_pad_GPIO_PAD[88]
  PIN gfpga_pad_GPIO_PAD[89]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 986.640 51.880 987.240 ;
    END
  END gfpga_pad_GPIO_PAD[89]
  PIN gfpga_pad_GPIO_PAD[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2013.770 44.120 2014.050 46.520 ;
    END
  END gfpga_pad_GPIO_PAD[8]
  PIN gfpga_pad_GPIO_PAD[90]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1040.360 51.880 1040.960 ;
    END
  END gfpga_pad_GPIO_PAD[90]
  PIN gfpga_pad_GPIO_PAD[91]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1094.080 51.880 1094.680 ;
    END
  END gfpga_pad_GPIO_PAD[91]
  PIN gfpga_pad_GPIO_PAD[92]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1148.480 51.880 1149.080 ;
    END
  END gfpga_pad_GPIO_PAD[92]
  PIN gfpga_pad_GPIO_PAD[93]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1202.200 51.880 1202.800 ;
    END
  END gfpga_pad_GPIO_PAD[93]
  PIN gfpga_pad_GPIO_PAD[94]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1255.920 51.880 1256.520 ;
    END
  END gfpga_pad_GPIO_PAD[94]
  PIN gfpga_pad_GPIO_PAD[95]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1309.640 51.880 1310.240 ;
    END
  END gfpga_pad_GPIO_PAD[95]
  PIN gfpga_pad_GPIO_PAD[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1848.880 51.880 1849.480 ;
    END
  END gfpga_pad_GPIO_PAD[9]
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2142.570 44.120 2142.850 46.520 ;
    END
  END reset
  PIN set
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1956.320 51.880 1956.920 ;
    END
  END set
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 2198.700 45.000 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 2223.700 20.000 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 97.925 104.915 2118.540 1975.915 ;
      LAYER met1 ;
        RECT 63.350 46.880 2151.150 1975.960 ;
      LAYER met2 ;
        RECT 63.370 1981.440 115.530 1981.720 ;
        RECT 116.370 1981.440 248.010 1981.720 ;
        RECT 248.850 1981.440 380.950 1981.720 ;
        RECT 381.790 1981.440 513.890 1981.720 ;
        RECT 514.730 1981.440 646.830 1981.720 ;
        RECT 647.670 1981.440 779.310 1981.720 ;
        RECT 780.150 1981.440 912.250 1981.720 ;
        RECT 913.090 1981.440 1045.190 1981.720 ;
        RECT 1046.030 1981.440 1178.130 1981.720 ;
        RECT 1178.970 1981.440 1310.610 1981.720 ;
        RECT 1311.450 1981.440 1443.550 1981.720 ;
        RECT 1444.390 1981.440 1576.490 1981.720 ;
        RECT 1577.330 1981.440 1709.430 1981.720 ;
        RECT 1710.270 1981.440 1841.910 1981.720 ;
        RECT 1842.750 1981.440 1974.850 1981.720 ;
        RECT 1975.690 1981.440 2107.790 1981.720 ;
        RECT 2108.630 1981.440 2151.130 1981.720 ;
        RECT 63.370 46.800 2151.130 1981.440 ;
        RECT 63.370 46.520 81.490 46.800 ;
        RECT 82.330 46.520 145.890 46.800 ;
        RECT 146.730 46.520 210.290 46.800 ;
        RECT 211.130 46.520 274.690 46.800 ;
        RECT 275.530 46.520 339.090 46.800 ;
        RECT 339.930 46.520 403.490 46.800 ;
        RECT 404.330 46.520 467.890 46.800 ;
        RECT 468.730 46.520 532.290 46.800 ;
        RECT 533.130 46.520 596.690 46.800 ;
        RECT 597.530 46.520 661.090 46.800 ;
        RECT 661.930 46.520 725.490 46.800 ;
        RECT 726.330 46.520 789.890 46.800 ;
        RECT 790.730 46.520 854.290 46.800 ;
        RECT 855.130 46.520 918.690 46.800 ;
        RECT 919.530 46.520 983.090 46.800 ;
        RECT 983.930 46.520 1047.490 46.800 ;
        RECT 1048.330 46.520 1111.890 46.800 ;
        RECT 1112.730 46.520 1176.290 46.800 ;
        RECT 1177.130 46.520 1240.690 46.800 ;
        RECT 1241.530 46.520 1305.090 46.800 ;
        RECT 1305.930 46.520 1369.490 46.800 ;
        RECT 1370.330 46.520 1433.890 46.800 ;
        RECT 1434.730 46.520 1498.290 46.800 ;
        RECT 1499.130 46.520 1562.690 46.800 ;
        RECT 1563.530 46.520 1627.090 46.800 ;
        RECT 1627.930 46.520 1691.490 46.800 ;
        RECT 1692.330 46.520 1755.890 46.800 ;
        RECT 1756.730 46.520 1820.290 46.800 ;
        RECT 1821.130 46.520 1884.690 46.800 ;
        RECT 1885.530 46.520 1949.090 46.800 ;
        RECT 1949.930 46.520 2013.490 46.800 ;
        RECT 2014.330 46.520 2077.890 46.800 ;
        RECT 2078.730 46.520 2142.290 46.800 ;
        RECT 2143.130 46.520 2151.130 46.800 ;
      LAYER met3 ;
        RECT 51.880 1957.320 2172.080 1969.025 ;
        RECT 52.280 1955.920 2172.080 1957.320 ;
        RECT 51.880 1953.920 2172.080 1955.920 ;
        RECT 51.880 1952.520 2171.680 1953.920 ;
        RECT 51.880 1903.600 2172.080 1952.520 ;
        RECT 52.280 1902.200 2172.080 1903.600 ;
        RECT 51.880 1893.400 2172.080 1902.200 ;
        RECT 51.880 1892.000 2171.680 1893.400 ;
        RECT 51.880 1849.880 2172.080 1892.000 ;
        RECT 52.280 1848.480 2172.080 1849.880 ;
        RECT 51.880 1832.880 2172.080 1848.480 ;
        RECT 51.880 1831.480 2171.680 1832.880 ;
        RECT 51.880 1796.160 2172.080 1831.480 ;
        RECT 52.280 1794.760 2172.080 1796.160 ;
        RECT 51.880 1772.360 2172.080 1794.760 ;
        RECT 51.880 1770.960 2171.680 1772.360 ;
        RECT 51.880 1741.760 2172.080 1770.960 ;
        RECT 52.280 1740.360 2172.080 1741.760 ;
        RECT 51.880 1711.840 2172.080 1740.360 ;
        RECT 51.880 1710.440 2171.680 1711.840 ;
        RECT 51.880 1688.040 2172.080 1710.440 ;
        RECT 52.280 1686.640 2172.080 1688.040 ;
        RECT 51.880 1651.320 2172.080 1686.640 ;
        RECT 51.880 1649.920 2171.680 1651.320 ;
        RECT 51.880 1634.320 2172.080 1649.920 ;
        RECT 52.280 1632.920 2172.080 1634.320 ;
        RECT 51.880 1590.120 2172.080 1632.920 ;
        RECT 51.880 1588.720 2171.680 1590.120 ;
        RECT 51.880 1580.600 2172.080 1588.720 ;
        RECT 52.280 1579.200 2172.080 1580.600 ;
        RECT 51.880 1529.600 2172.080 1579.200 ;
        RECT 51.880 1528.200 2171.680 1529.600 ;
        RECT 51.880 1526.200 2172.080 1528.200 ;
        RECT 52.280 1524.800 2172.080 1526.200 ;
        RECT 51.880 1472.480 2172.080 1524.800 ;
        RECT 52.280 1471.080 2172.080 1472.480 ;
        RECT 51.880 1469.080 2172.080 1471.080 ;
        RECT 51.880 1467.680 2171.680 1469.080 ;
        RECT 51.880 1418.760 2172.080 1467.680 ;
        RECT 52.280 1417.360 2172.080 1418.760 ;
        RECT 51.880 1408.560 2172.080 1417.360 ;
        RECT 51.880 1407.160 2171.680 1408.560 ;
        RECT 51.880 1365.040 2172.080 1407.160 ;
        RECT 52.280 1363.640 2172.080 1365.040 ;
        RECT 51.880 1348.040 2172.080 1363.640 ;
        RECT 51.880 1346.640 2171.680 1348.040 ;
        RECT 51.880 1310.640 2172.080 1346.640 ;
        RECT 52.280 1309.240 2172.080 1310.640 ;
        RECT 51.880 1287.520 2172.080 1309.240 ;
        RECT 51.880 1286.120 2171.680 1287.520 ;
        RECT 51.880 1256.920 2172.080 1286.120 ;
        RECT 52.280 1255.520 2172.080 1256.920 ;
        RECT 51.880 1226.320 2172.080 1255.520 ;
        RECT 51.880 1224.920 2171.680 1226.320 ;
        RECT 51.880 1203.200 2172.080 1224.920 ;
        RECT 52.280 1201.800 2172.080 1203.200 ;
        RECT 51.880 1165.800 2172.080 1201.800 ;
        RECT 51.880 1164.400 2171.680 1165.800 ;
        RECT 51.880 1149.480 2172.080 1164.400 ;
        RECT 52.280 1148.080 2172.080 1149.480 ;
        RECT 51.880 1105.280 2172.080 1148.080 ;
        RECT 51.880 1103.880 2171.680 1105.280 ;
        RECT 51.880 1095.080 2172.080 1103.880 ;
        RECT 52.280 1093.680 2172.080 1095.080 ;
        RECT 51.880 1044.760 2172.080 1093.680 ;
        RECT 51.880 1043.360 2171.680 1044.760 ;
        RECT 51.880 1041.360 2172.080 1043.360 ;
        RECT 52.280 1039.960 2172.080 1041.360 ;
        RECT 51.880 987.640 2172.080 1039.960 ;
        RECT 52.280 986.240 2172.080 987.640 ;
        RECT 51.880 984.240 2172.080 986.240 ;
        RECT 51.880 982.840 2171.680 984.240 ;
        RECT 51.880 933.920 2172.080 982.840 ;
        RECT 52.280 932.520 2172.080 933.920 ;
        RECT 51.880 923.720 2172.080 932.520 ;
        RECT 51.880 922.320 2171.680 923.720 ;
        RECT 51.880 879.520 2172.080 922.320 ;
        RECT 52.280 878.120 2172.080 879.520 ;
        RECT 51.880 863.200 2172.080 878.120 ;
        RECT 51.880 861.800 2171.680 863.200 ;
        RECT 51.880 825.800 2172.080 861.800 ;
        RECT 52.280 824.400 2172.080 825.800 ;
        RECT 51.880 802.000 2172.080 824.400 ;
        RECT 51.880 800.600 2171.680 802.000 ;
        RECT 51.880 772.080 2172.080 800.600 ;
        RECT 52.280 770.680 2172.080 772.080 ;
        RECT 51.880 741.480 2172.080 770.680 ;
        RECT 51.880 740.080 2171.680 741.480 ;
        RECT 51.880 718.360 2172.080 740.080 ;
        RECT 52.280 716.960 2172.080 718.360 ;
        RECT 51.880 680.960 2172.080 716.960 ;
        RECT 51.880 679.560 2171.680 680.960 ;
        RECT 51.880 663.960 2172.080 679.560 ;
        RECT 52.280 662.560 2172.080 663.960 ;
        RECT 51.880 620.440 2172.080 662.560 ;
        RECT 51.880 619.040 2171.680 620.440 ;
        RECT 51.880 610.240 2172.080 619.040 ;
        RECT 52.280 608.840 2172.080 610.240 ;
        RECT 51.880 559.920 2172.080 608.840 ;
        RECT 51.880 558.520 2171.680 559.920 ;
        RECT 51.880 556.520 2172.080 558.520 ;
        RECT 52.280 555.120 2172.080 556.520 ;
        RECT 51.880 502.800 2172.080 555.120 ;
        RECT 52.280 501.400 2172.080 502.800 ;
        RECT 51.880 499.400 2172.080 501.400 ;
        RECT 51.880 498.000 2171.680 499.400 ;
        RECT 51.880 448.400 2172.080 498.000 ;
        RECT 52.280 447.000 2172.080 448.400 ;
        RECT 51.880 438.200 2172.080 447.000 ;
        RECT 51.880 436.800 2171.680 438.200 ;
        RECT 51.880 394.680 2172.080 436.800 ;
        RECT 52.280 393.280 2172.080 394.680 ;
        RECT 51.880 377.680 2172.080 393.280 ;
        RECT 51.880 376.280 2171.680 377.680 ;
        RECT 51.880 340.960 2172.080 376.280 ;
        RECT 52.280 339.560 2172.080 340.960 ;
        RECT 51.880 317.160 2172.080 339.560 ;
        RECT 51.880 315.760 2171.680 317.160 ;
        RECT 51.880 287.240 2172.080 315.760 ;
        RECT 52.280 285.840 2172.080 287.240 ;
        RECT 51.880 256.640 2172.080 285.840 ;
        RECT 51.880 255.240 2171.680 256.640 ;
        RECT 51.880 232.840 2172.080 255.240 ;
        RECT 52.280 231.440 2172.080 232.840 ;
        RECT 51.880 196.120 2172.080 231.440 ;
        RECT 51.880 194.720 2171.680 196.120 ;
        RECT 51.880 179.120 2172.080 194.720 ;
        RECT 52.280 177.720 2172.080 179.120 ;
        RECT 51.880 135.600 2172.080 177.720 ;
        RECT 51.880 134.200 2171.680 135.600 ;
        RECT 51.880 125.400 2172.080 134.200 ;
        RECT 52.280 124.000 2172.080 125.400 ;
        RECT 51.880 75.080 2172.080 124.000 ;
        RECT 51.880 73.680 2171.680 75.080 ;
        RECT 51.880 71.680 2172.080 73.680 ;
        RECT 52.280 70.815 2172.080 71.680 ;
      LAYER met4 ;
        RECT 0.000 0.000 2223.700 2027.600 ;
      LAYER met5 ;
        RECT 0.000 70.850 2223.700 2027.600 ;
  END
END fpga_top
END LIBRARY

