* NGSPICE file created from sb_0__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt sb_0__2_ SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_left_grid_pin_1_
+ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] prog_clk right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ right_top_grid_pin_1_
+ VPWR VGND
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_20.mux_l1_in_0_/S
+ mux_right_track_20.mux_l2_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_18.mux_l1_in_0__S mux_right_track_18.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_83_ chanx_right_in[11] chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_66_ _66_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_36.mux_l2_in_0__A1 mux_right_track_36.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X _52_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_prog_clk_A clkbuf_1_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_49_ _49_/A SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__D mux_bottom_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A mux_right_track_22.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_38.mux_l1_in_0_ chany_bottom_in[19] right_bottom_grid_pin_40_ mux_right_track_38.mux_l1_in_0_/S
+ mux_right_track_38.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_18.mux_l2_in_0_/S
+ mux_right_track_20.mux_l1_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_82_ chanx_right_in[10] chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0__A0 _40_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_65_ _65_/A chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_6.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_48_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_25.mux_l1_in_0_/S
+ ccff_tail clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_1__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_81_ chanx_right_in[9] chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_20.mux_l2_in_0__S mux_right_track_20.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l2_in_0__A1 mux_right_track_10.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A mux_right_track_28.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_64_ _64_/A chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_6.mux_l2_in_0__A0 mux_right_track_6.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0__S mux_right_track_14.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_47_ _47_/HI _47_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_prog_clk clkbuf_1_0_0_prog_clk/X clkbuf_2_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_6.mux_l1_in_1__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_80_ chanx_right_in[8] chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0__S mux_right_track_6.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0__A1 mux_right_track_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ _63_/A chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_14.mux_l1_in_0__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_46_ _46_/HI _46_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_10.mux_l2_in_0_ _40_/HI mux_right_track_10.mux_l1_in_0_/X mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_29_ _29_/HI _29_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_5.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l1_in_0__A0 chany_bottom_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_62_ _62_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l2_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_45_ _45_/HI _45_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_10.mux_l1_in_0__S mux_right_track_10.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_38.mux_l2_in_0__S mux_right_track_38.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_28_ _28_/HI _28_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l2_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_10.mux_l1_in_0_ chany_bottom_in[13] right_bottom_grid_pin_34_ mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_30.mux_l1_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_22.mux_l2_in_0_ _47_/HI mux_right_track_22.mux_l1_in_0_/X mux_right_track_22.mux_l2_in_0_/S
+ mux_right_track_22.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_22.mux_l1_in_0__A1 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_1_ _34_/HI chany_bottom_in[14] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ _61_/A chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_44_ _44_/HI _44_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l2_in_0_/X _65_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27_ _27_/HI _27_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A mux_right_track_14.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_30.mux_l1_in_0__A1 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_8.mux_l1_in_0_ right_bottom_grid_pin_41_ right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l2_in_1__S mux_right_track_6.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_prog_clk clkbuf_1_0_0_prog_clk/X clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_22.mux_l1_in_0_ chany_bottom_in[7] right_bottom_grid_pin_40_ mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_60_ _60_/A chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_18.mux_l1_in_0_/S
+ mux_right_track_18.mux_l2_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 _38_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_34.mux_l2_in_0_ _29_/HI mux_right_track_34.mux_l1_in_0_/X mux_right_track_34.mux_l2_in_0_/S
+ mux_right_track_34.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 _43_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l2_in_0_/X _66_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_43_ _43_/HI _43_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_26_ _26_/HI _26_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_34.mux_l2_in_0__S mux_right_track_34.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 _24_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X _54_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_28.mux_l1_in_0__S mux_right_track_28.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X _57_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_18.mux_l1_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__53__A _53_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_0_ _36_/HI mux_bottom_track_25.mux_l1_in_0_/X ccff_tail
+ mux_bottom_track_25.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_42_ _42_/HI _42_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__48__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_34.mux_l1_in_0_ chany_bottom_in[1] right_bottom_grid_pin_38_ mux_right_track_34.mux_l1_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_25_ _25_/HI _25_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ _38_/HI mux_bottom_track_9.mux_l1_in_0_/X mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_2_0_prog_clk_A clkbuf_2_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_bottom_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 _28_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__61__A _61_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__56__A _56_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A mux_right_track_6.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_41_ _41_/HI _41_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA__64__A _64_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24_ _24_/HI _24_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[6] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__59__A _59_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_36.mux_l1_in_0_/S
+ mux_right_track_36.mux_l2_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_30.mux_l2_in_0__S mux_right_track_30.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[14] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__72__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l2_in_0_/X _86_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__67__A _67_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_28.mux_l1_in_0__A0 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_40_ _40_/HI _40_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__80__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__75__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_38.sky130_fd_sc_hd__buf_4_0__A mux_right_track_38.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_34.mux_l2_in_0_/S
+ mux_right_track_36.mux_l1_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_36.mux_l1_in_0__A0 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__83__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_28.mux_l1_in_0__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__78__A _78_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l3_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_1_ _32_/HI mux_right_track_4.mux_l1_in_2_/X mux_right_track_4.mux_l2_in_0_/S
+ mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_2_ chany_bottom_in[16] right_bottom_grid_pin_41_ mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__86__A _86_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_36.mux_l1_in_0__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_20.mux_l1_in_0__S mux_right_track_20.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l2_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l2_in_0_ _43_/HI mux_right_track_16.mux_l1_in_0_/X mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_0_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__89__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_12.mux_l2_in_0__S mux_right_track_12.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l2_in_0_/S clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_1_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l1_in_0_ chany_bottom_in[10] right_bottom_grid_pin_37_ mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ right_bottom_grid_pin_35_ right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_28.mux_l2_in_0_ _26_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _68_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_30.mux_l2_in_0_ _27_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_38.mux_l2_in_0__A0 _31_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_20.mux_l2_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__D mux_bottom_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 _32_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X _59_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_79_ chanx_right_in[7] chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_38.mux_l1_in_0__S mux_right_track_38.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X _62_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_38.mux_l2_in_0__A1 mux_right_track_38.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l1_in_0_ chany_bottom_in[4] right_bottom_grid_pin_35_ mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_30.mux_l1_in_0_ chany_bottom_in[3] right_bottom_grid_pin_36_ mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_0_ _37_/HI mux_bottom_track_5.mux_l1_in_0_/X mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_78_ _78_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 _37_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0__A0 _41_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_1.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_38.sky130_fd_sc_hd__buf_4_0_ mux_right_track_38.mux_l2_in_0_/X _51_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_2_3_0_prog_clk_A clkbuf_2_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_1__S mux_right_track_6.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l2_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l2_in_0_/X _88_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1__A0 _34_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_77_ chanx_right_in[5] chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_20.mux_l2_in_0__A0 _46_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[16] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_12.mux_l2_in_0__A1 mux_right_track_12.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 mux_right_track_8.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_34.mux_l1_in_0__S mux_right_track_34.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_76_ chanx_right_in[4] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_20.mux_l2_in_0__A1 mux_right_track_20.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_26.mux_l2_in_0__S mux_right_track_26.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A mux_right_track_10.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_59_ _59_/A chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_1_ _39_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l2_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[18] right_bottom_grid_pin_41_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_75_ chanx_right_in[3] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_58_ _58_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_30.mux_l1_in_0__S mux_right_track_30.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A mux_right_track_16.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.mux_l2_in_0_ _41_/HI mux_right_track_12.mux_l1_in_0_/X mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_12.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_74_ chanx_right_in[2] chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_57_ _57_/A chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__51__A _51_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_22.mux_l2_in_0__S mux_right_track_22.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A mux_right_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _70_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__D mux_bottom_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_90_ _90_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_12.mux_l1_in_0_ chany_bottom_in[12] right_bottom_grid_pin_35_ mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_35_ right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_1_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__54__A _54_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_14.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_73_ chanx_right_in[1] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_56_ _56_/A chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_24.mux_l1_in_1_ _24_/HI chany_bottom_in[6] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_18.mux_l2_in_0__A0 _44_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_39_ _39_/HI _39_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__62__A _62_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__57__A _57_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l2_in_0_/X _64_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__70__A _70_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_72_ chanx_right_in[0] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_26.mux_l2_in_0__A0 _25_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__65__A _65_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l3_in_0__S mux_right_track_6.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_55_ _55_/A chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_41_ right_top_grid_pin_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A mux_right_track_34.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_36.mux_l2_in_0_ _30_/HI mux_right_track_36.mux_l1_in_0_/X mux_right_track_36.mux_l2_in_0_/S
+ mux_right_track_36.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_18.mux_l2_in_0__A1 mux_right_track_18.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ _38_/HI _38_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_0_ _35_/HI mux_bottom_track_1.mux_l1_in_0_/X mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__73__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l1_in_0__S mux_right_track_12.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_38.mux_l1_in_0_/S
+ mux_right_track_38.mux_l2_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__68__A _68_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X _53_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_34.mux_l2_in_0__A0 _29_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_71_ chanx_right_in[19] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_26.mux_l2_in_0__A1 mux_right_track_26.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__81__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_54_ _54_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X _56_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__76__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ _37_/HI _37_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 _39_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l2_in_0_/X _90_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_36.mux_l1_in_0_ chany_bottom_in[0] right_bottom_grid_pin_39_ mux_right_track_36.mux_l1_in_0_/S
+ mux_right_track_36.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_36.mux_l2_in_0_/S
+ mux_right_track_38.mux_l1_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_1_ chanx_right_in[18] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__84__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_0.mux_l1_in_1_/S mux_right_track_0.mux_l2_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_18.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_34.mux_l2_in_0__A1 mux_right_track_34.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__79__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_70_ _70_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_53_ _53_/A chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l3_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_36_ _36_/HI _36_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__87__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 _35_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_right_track_0.mux_l1_in_1_/S
+ clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_36.mux_l2_in_0__S mux_right_track_36.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_38.mux_l1_in_0__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_52_ _52_/A chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l2_in_1_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35_ _35_/HI _35_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A mux_right_track_20.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_38.mux_l1_in_0__A1 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_51_ _51_/A chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/S clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_6.mux_l1_in_1_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S mux_right_track_6.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_34_ _34_/HI _34_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_1_ _33_/HI chany_bottom_in[15] mux_right_track_6.mux_l2_in_1_/S
+ mux_right_track_6.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_20.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0__A0 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A mux_right_track_26.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_50_ _50_/A SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_22.mux_l2_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_26.mux_l1_in_0__S mux_right_track_26.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33_ _33_/HI _33_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.mux_l2_in_0_ _44_/HI mux_right_track_18.mux_l1_in_0_/X mux_right_track_18.mux_l2_in_0_/S
+ mux_right_track_18.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_1_/S mux_right_track_6.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l2_in_0_ _46_/HI mux_right_track_20.mux_l1_in_0_/X mux_right_track_20.mux_l2_in_0_/S
+ mux_right_track_20.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_20.mux_l1_in_0__A0 chany_bottom_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_6.mux_l1_in_1_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l2_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__D mux_right_track_6.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_18.mux_l2_in_0__S mux_right_track_18.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ _32_/HI _32_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l2_in_1__A0 _33_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_20.mux_l1_in_0__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l3_in_0__A0 mux_right_track_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_18.mux_l1_in_0_ chany_bottom_in[9] right_bottom_grid_pin_38_ mux_right_track_18.mux_l1_in_0_/S
+ mux_right_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l1_in_0_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_38.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/S clkbuf_2_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l2_in_0_/X
+ _78_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_20.mux_l1_in_0_ chany_bottom_in[8] right_bottom_grid_pin_39_ mux_right_track_20.mux_l1_in_0_/S
+ mux_right_track_20.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.mux_l2_in_0_ _28_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X _67_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31_ _31_/HI _31_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X _55_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_6.mux_l2_in_1__A1 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l1_in_0__S mux_right_track_22.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l2_in_0_/X _58_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l2_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l3_in_0__A1 mux_right_track_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_14.mux_l2_in_0__A0 _42_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X _61_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_9.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l1_in_0_ chany_bottom_in[2] right_bottom_grid_pin_37_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_30_ _30_/HI _30_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0__S mux_right_track_14.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_0_0_prog_clk_A clkbuf_1_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A mux_right_track_12.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_10.mux_l1_in_0_/S
+ clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_22.mux_l2_in_0__A0 _47_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_14.mux_l2_in_0__A1 mux_right_track_14.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l2_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0__S mux_right_track_6.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_89_ chanx_right_in[17] chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_30.mux_l2_in_0__A0 _27_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l2_in_0__A1 mux_right_track_22.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A mux_right_track_18.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_18.mux_l1_in_0__A0 chany_bottom_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_14.mux_l2_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/S clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_88_ _88_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_30.mux_l2_in_0__A1 mux_right_track_30.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__52__A _52_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 _36_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0__S mux_right_track_10.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_26.mux_l1_in_0__A0 chany_bottom_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__D mux_bottom_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__60__A _60_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__55__A _55_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l2_in_1_ _45_/HI chany_bottom_in[17] mux_right_track_2.mux_l2_in_1_/S
+ mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A mux_right_track_30.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_87_ chanx_right_in[15] chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__63__A _63_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_34.mux_l1_in_0__A0 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__D mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_34.mux_l1_in_0_/S
+ mux_right_track_34.mux_l2_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__58__A _58_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_36.mux_l1_in_0__S mux_right_track_36.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__71__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_14.mux_l2_in_0_ _42_/HI mux_right_track_14.mux_l1_in_0_/X mux_right_track_14.mux_l2_in_0_/S
+ mux_right_track_14.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__66__A _66_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_86_ _86_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_69_ _69_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK clkbuf_2_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_34.mux_l1_in_0__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A mux_right_track_36.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/S clkbuf_2_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__74__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_28.mux_l2_in_0__S mux_right_track_28.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__69__A _69_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_2.mux_l2_in_1_/S mux_right_track_2.mux_l3_in_0_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__82__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_85_ chanx_right_in[13] chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK clkbuf_2_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _69_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_14.mux_l1_in_0_ chany_bottom_in[11] right_bottom_grid_pin_36_ mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__77__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_0_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_26.mux_l2_in_0_ _25_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_68_ _68_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_28.mux_l2_in_0__A0 _26_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__90__A _90_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__85__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X _60_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_1_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_1_/S
+ clkbuf_2_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_84_ chanx_right_in[12] chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l2_in_0_/X _63_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK clkbuf_2_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_67_ _67_/A chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_36.mux_l2_in_0__A0 _30_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__D mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__88__A _88_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_28.mux_l2_in_0__A1 mux_right_track_28.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_26.mux_l1_in_0_ chany_bottom_in[5] right_bottom_grid_pin_34_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_38.mux_l2_in_0_ _31_/HI mux_right_track_38.mux_l1_in_0_/X mux_right_track_38.mux_l2_in_0_/S
+ mux_right_track_38.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 _45_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_25.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

