VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2495.000 BY 2865.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END IO_ISOL_N
  PIN Test_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 2684.680 2495.000 2685.280 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 2861.000 46.370 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 536.560 2495.000 537.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 894.240 2495.000 894.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1252.600 2495.000 1253.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1610.960 2495.000 1611.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1968.640 2495.000 1969.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 2327.000 2495.000 2327.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.770 0.000 2189.050 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2200.270 0.000 2200.550 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2211.770 0.000 2212.050 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2223.270 0.000 2223.550 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 2861.000 138.370 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.770 0.000 2235.050 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.270 0.000 2246.550 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.770 0.000 2258.050 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2269.270 0.000 2269.550 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.770 0.000 2281.050 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.890 0.000 1877.170 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.390 0.000 1888.670 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.890 0.000 1900.170 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.390 0.000 1911.670 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.890 0.000 1923.170 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 2861.000 230.830 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.390 0.000 1934.670 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.890 0.000 1946.170 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.390 0.000 1957.670 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.890 0.000 1969.170 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.010 0.000 1565.290 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.510 0.000 1576.790 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.010 0.000 1588.290 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.510 0.000 1599.790 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.010 0.000 1611.290 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 0.000 1622.790 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 2861.000 323.290 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.010 0.000 1634.290 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.510 0.000 1645.790 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.010 0.000 1657.290 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 0.000 1253.410 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.630 0.000 1264.910 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.130 0.000 1276.410 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.630 0.000 1287.910 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 0.000 1322.410 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 2861.000 415.750 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 0.000 1333.910 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.130 0.000 1345.410 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 0.000 953.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 0.000 964.530 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 0.000 1010.530 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 0.000 1022.030 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 2861.000 508.210 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 0.000 710.150 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 2861.000 600.670 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 2861.000 693.130 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 2861.000 785.590 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1629.320 4.000 1629.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1925.800 4.000 1926.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2222.280 4.000 2222.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2518.080 4.000 2518.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 178.200 2495.000 178.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 2861.000 878.050 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 655.560 2495.000 656.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1013.920 2495.000 1014.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1371.600 2495.000 1372.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1729.960 2495.000 1730.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 2088.320 2495.000 2088.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 2446.000 2495.000 2446.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.730 0.000 2293.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.230 0.000 2304.510 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.730 0.000 2316.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2327.230 0.000 2327.510 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 2861.000 970.050 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.730 0.000 2339.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.230 0.000 2350.510 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.730 0.000 2362.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.230 0.000 2373.510 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.730 0.000 2385.010 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.850 0.000 1981.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.350 0.000 1992.630 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.850 0.000 2004.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.350 0.000 2015.630 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.850 0.000 2027.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 2861.000 1062.510 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.350 0.000 2038.630 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2049.850 0.000 2050.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2061.350 0.000 2061.630 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.850 0.000 2073.130 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.970 0.000 1669.250 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.470 0.000 1680.750 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 0.000 1692.250 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.470 0.000 1703.750 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.970 0.000 1715.250 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.470 0.000 1726.750 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 2861.000 1154.970 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.970 0.000 1738.250 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.470 0.000 1749.750 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 0.000 1761.250 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.090 0.000 1357.370 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 0.000 1380.370 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.590 0.000 1391.870 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.590 0.000 1414.870 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.090 0.000 1426.370 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 2861.000 1247.430 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 0.000 1437.870 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 0.000 1056.990 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 0.000 1068.490 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 2861.000 1339.890 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 0.000 768.110 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 0.000 791.110 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 0.000 825.610 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 2861.000 1432.350 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.530 2861.000 1524.810 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 2861.000 1617.270 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.920 4.000 1728.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2024.400 4.000 2025.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2320.880 4.000 2321.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2617.360 4.000 2617.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 297.880 2495.000 298.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.450 2861.000 1709.730 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 775.240 2495.000 775.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1132.920 2495.000 1133.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1491.280 2495.000 1491.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 1849.640 2495.000 1850.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 2207.320 2495.000 2207.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 2565.680 2495.000 2566.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.690 0.000 2396.970 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.190 0.000 2408.470 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.690 0.000 2419.970 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.190 0.000 2431.470 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.450 2861.000 1801.730 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2442.690 0.000 2442.970 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2454.190 0.000 2454.470 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2465.690 0.000 2465.970 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.190 0.000 2477.470 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.690 0.000 2488.970 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.810 0.000 2085.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.310 0.000 2096.590 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.810 0.000 2108.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.310 0.000 2119.590 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.810 0.000 2131.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.910 2861.000 1894.190 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.310 0.000 2142.590 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2153.810 0.000 2154.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.310 0.000 2165.590 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.810 0.000 2177.090 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.930 0.000 1773.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.430 0.000 1784.710 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.930 0.000 1796.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.430 0.000 1807.710 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.930 0.000 1819.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1830.430 0.000 1830.710 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.370 2861.000 1986.650 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 0.000 1842.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.430 0.000 1853.710 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.930 0.000 1865.210 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.050 0.000 1461.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 0.000 1472.830 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 0.000 1484.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.550 0.000 1495.830 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 0.000 1507.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.550 0.000 1518.830 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.050 0.000 1530.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.830 2861.000 2079.110 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.550 0.000 1541.830 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.050 0.000 1553.330 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.170 0.000 1149.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 0.000 1160.950 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 0.000 1172.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.670 0.000 1206.950 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.670 0.000 1229.950 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.290 2861.000 2171.570 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 0.000 883.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290 0.000 906.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.750 2861.000 2264.030 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.210 2861.000 2356.490 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.760 4.000 938.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2448.670 2861.000 2448.950 2865.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1530.720 4.000 1531.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1826.520 4.000 1827.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2123.000 4.000 2123.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2419.480 4.000 2420.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2715.960 4.000 2716.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 416.880 2495.000 417.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 59.200 2495.000 59.800 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2814.560 4.000 2815.160 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2491.000 2804.360 2495.000 2804.960 ;
    END
  END sc_tail
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2844.380 2489.060 2847.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2799.380 2489.060 2802.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2754.380 2489.060 2757.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2709.380 2489.060 2712.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2664.380 2489.060 2667.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2619.380 2489.060 2622.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2574.380 2489.060 2577.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2529.380 2489.060 2532.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2484.380 2489.060 2487.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2439.380 2489.060 2442.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2394.380 2489.060 2397.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2349.380 2489.060 2352.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2304.380 2489.060 2307.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2259.380 2489.060 2262.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2214.380 2489.060 2217.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2169.380 2489.060 2172.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2124.380 2489.060 2127.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2079.380 2489.060 2082.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 2034.380 2489.060 2037.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1989.380 2489.060 1992.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1944.380 2489.060 1947.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1899.380 2489.060 1902.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1854.380 2489.060 1857.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1809.380 2489.060 1812.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1764.380 2489.060 1767.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1719.380 2489.060 1722.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1674.380 2489.060 1677.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1629.380 2489.060 1632.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1584.380 2489.060 1587.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1539.380 2489.060 1542.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1494.380 2489.060 1497.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1449.380 2489.060 1452.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1404.380 2489.060 1407.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1359.380 2489.060 1362.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1314.380 2489.060 1317.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1269.380 2489.060 1272.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1224.380 2489.060 1227.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1179.380 2489.060 1182.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1134.380 2489.060 1137.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1089.380 2489.060 1092.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1044.380 2489.060 1047.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 999.380 2489.060 1002.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 954.380 2489.060 957.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 909.380 2489.060 912.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 864.380 2489.060 867.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 819.380 2489.060 822.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 774.380 2489.060 777.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 729.380 2489.060 732.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 684.380 2489.060 687.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 639.380 2489.060 642.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 594.380 2489.060 597.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 549.380 2489.060 552.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 504.380 2489.060 507.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 459.380 2489.060 462.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 414.380 2489.060 417.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 369.380 2489.060 372.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 324.380 2489.060 327.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 279.380 2489.060 282.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 234.380 2489.060 237.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 189.380 2489.060 192.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 144.380 2489.060 147.380 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 99.380 2489.060 102.380 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2821.880 2489.060 2824.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2776.880 2489.060 2779.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2731.880 2489.060 2734.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2686.880 2489.060 2689.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2641.880 2489.060 2644.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2596.880 2489.060 2599.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2551.880 2489.060 2554.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2506.880 2489.060 2509.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2461.880 2489.060 2464.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2416.880 2489.060 2419.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2371.880 2489.060 2374.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2326.880 2489.060 2329.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2281.880 2489.060 2284.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2236.880 2489.060 2239.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2191.880 2489.060 2194.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2146.880 2489.060 2149.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2101.880 2489.060 2104.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2056.880 2489.060 2059.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 2011.880 2489.060 2014.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1966.880 2489.060 1969.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1921.880 2489.060 1924.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1876.880 2489.060 1879.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1831.880 2489.060 1834.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1786.880 2489.060 1789.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1741.880 2489.060 1744.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1696.880 2489.060 1699.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1651.880 2489.060 1654.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1606.880 2489.060 1609.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1561.880 2489.060 1564.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1516.880 2489.060 1519.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1471.880 2489.060 1474.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1426.880 2489.060 1429.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1381.880 2489.060 1384.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1336.880 2489.060 1339.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1291.880 2489.060 1294.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1246.880 2489.060 1249.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1201.880 2489.060 1204.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1156.880 2489.060 1159.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1111.880 2489.060 1114.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1066.880 2489.060 1069.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1021.880 2489.060 1024.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 976.880 2489.060 979.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 931.880 2489.060 934.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 886.880 2489.060 889.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 841.880 2489.060 844.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 796.880 2489.060 799.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 751.880 2489.060 754.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 706.880 2489.060 709.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 661.880 2489.060 664.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 616.880 2489.060 619.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 571.880 2489.060 574.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 526.880 2489.060 529.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 481.880 2489.060 484.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 436.880 2489.060 439.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 391.880 2489.060 394.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 346.880 2489.060 349.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 301.880 2489.060 304.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.880 2489.060 259.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 211.880 2489.060 214.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 166.880 2489.060 169.880 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 121.880 2489.060 124.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 34.185 15.385 2440.255 2850.205 ;
      LAYER met1 ;
        RECT 5.590 13.980 2488.990 2850.360 ;
      LAYER met2 ;
        RECT 5.620 2860.720 45.810 2861.000 ;
        RECT 46.650 2860.720 137.810 2861.000 ;
        RECT 138.650 2860.720 230.270 2861.000 ;
        RECT 231.110 2860.720 322.730 2861.000 ;
        RECT 323.570 2860.720 415.190 2861.000 ;
        RECT 416.030 2860.720 507.650 2861.000 ;
        RECT 508.490 2860.720 600.110 2861.000 ;
        RECT 600.950 2860.720 692.570 2861.000 ;
        RECT 693.410 2860.720 785.030 2861.000 ;
        RECT 785.870 2860.720 877.490 2861.000 ;
        RECT 878.330 2860.720 969.490 2861.000 ;
        RECT 970.330 2860.720 1061.950 2861.000 ;
        RECT 1062.790 2860.720 1154.410 2861.000 ;
        RECT 1155.250 2860.720 1246.870 2861.000 ;
        RECT 1247.710 2860.720 1339.330 2861.000 ;
        RECT 1340.170 2860.720 1431.790 2861.000 ;
        RECT 1432.630 2860.720 1524.250 2861.000 ;
        RECT 1525.090 2860.720 1616.710 2861.000 ;
        RECT 1617.550 2860.720 1709.170 2861.000 ;
        RECT 1710.010 2860.720 1801.170 2861.000 ;
        RECT 1802.010 2860.720 1893.630 2861.000 ;
        RECT 1894.470 2860.720 1986.090 2861.000 ;
        RECT 1986.930 2860.720 2078.550 2861.000 ;
        RECT 2079.390 2860.720 2171.010 2861.000 ;
        RECT 2171.850 2860.720 2263.470 2861.000 ;
        RECT 2264.310 2860.720 2355.930 2861.000 ;
        RECT 2356.770 2860.720 2448.390 2861.000 ;
        RECT 2449.230 2860.720 2488.960 2861.000 ;
        RECT 5.620 4.280 2488.960 2860.720 ;
        RECT 6.170 4.000 16.830 4.280 ;
        RECT 17.670 4.000 28.330 4.280 ;
        RECT 29.170 4.000 39.830 4.280 ;
        RECT 40.670 4.000 51.330 4.280 ;
        RECT 52.170 4.000 62.830 4.280 ;
        RECT 63.670 4.000 74.330 4.280 ;
        RECT 75.170 4.000 85.830 4.280 ;
        RECT 86.670 4.000 97.330 4.280 ;
        RECT 98.170 4.000 109.290 4.280 ;
        RECT 110.130 4.000 120.790 4.280 ;
        RECT 121.630 4.000 132.290 4.280 ;
        RECT 133.130 4.000 143.790 4.280 ;
        RECT 144.630 4.000 155.290 4.280 ;
        RECT 156.130 4.000 166.790 4.280 ;
        RECT 167.630 4.000 178.290 4.280 ;
        RECT 179.130 4.000 189.790 4.280 ;
        RECT 190.630 4.000 201.290 4.280 ;
        RECT 202.130 4.000 213.250 4.280 ;
        RECT 214.090 4.000 224.750 4.280 ;
        RECT 225.590 4.000 236.250 4.280 ;
        RECT 237.090 4.000 247.750 4.280 ;
        RECT 248.590 4.000 259.250 4.280 ;
        RECT 260.090 4.000 270.750 4.280 ;
        RECT 271.590 4.000 282.250 4.280 ;
        RECT 283.090 4.000 293.750 4.280 ;
        RECT 294.590 4.000 305.250 4.280 ;
        RECT 306.090 4.000 317.210 4.280 ;
        RECT 318.050 4.000 328.710 4.280 ;
        RECT 329.550 4.000 340.210 4.280 ;
        RECT 341.050 4.000 351.710 4.280 ;
        RECT 352.550 4.000 363.210 4.280 ;
        RECT 364.050 4.000 374.710 4.280 ;
        RECT 375.550 4.000 386.210 4.280 ;
        RECT 387.050 4.000 397.710 4.280 ;
        RECT 398.550 4.000 409.210 4.280 ;
        RECT 410.050 4.000 421.170 4.280 ;
        RECT 422.010 4.000 432.670 4.280 ;
        RECT 433.510 4.000 444.170 4.280 ;
        RECT 445.010 4.000 455.670 4.280 ;
        RECT 456.510 4.000 467.170 4.280 ;
        RECT 468.010 4.000 478.670 4.280 ;
        RECT 479.510 4.000 490.170 4.280 ;
        RECT 491.010 4.000 501.670 4.280 ;
        RECT 502.510 4.000 513.170 4.280 ;
        RECT 514.010 4.000 525.130 4.280 ;
        RECT 525.970 4.000 536.630 4.280 ;
        RECT 537.470 4.000 548.130 4.280 ;
        RECT 548.970 4.000 559.630 4.280 ;
        RECT 560.470 4.000 571.130 4.280 ;
        RECT 571.970 4.000 582.630 4.280 ;
        RECT 583.470 4.000 594.130 4.280 ;
        RECT 594.970 4.000 605.630 4.280 ;
        RECT 606.470 4.000 617.130 4.280 ;
        RECT 617.970 4.000 629.090 4.280 ;
        RECT 629.930 4.000 640.590 4.280 ;
        RECT 641.430 4.000 652.090 4.280 ;
        RECT 652.930 4.000 663.590 4.280 ;
        RECT 664.430 4.000 675.090 4.280 ;
        RECT 675.930 4.000 686.590 4.280 ;
        RECT 687.430 4.000 698.090 4.280 ;
        RECT 698.930 4.000 709.590 4.280 ;
        RECT 710.430 4.000 721.090 4.280 ;
        RECT 721.930 4.000 733.050 4.280 ;
        RECT 733.890 4.000 744.550 4.280 ;
        RECT 745.390 4.000 756.050 4.280 ;
        RECT 756.890 4.000 767.550 4.280 ;
        RECT 768.390 4.000 779.050 4.280 ;
        RECT 779.890 4.000 790.550 4.280 ;
        RECT 791.390 4.000 802.050 4.280 ;
        RECT 802.890 4.000 813.550 4.280 ;
        RECT 814.390 4.000 825.050 4.280 ;
        RECT 825.890 4.000 837.010 4.280 ;
        RECT 837.850 4.000 848.510 4.280 ;
        RECT 849.350 4.000 860.010 4.280 ;
        RECT 860.850 4.000 871.510 4.280 ;
        RECT 872.350 4.000 883.010 4.280 ;
        RECT 883.850 4.000 894.510 4.280 ;
        RECT 895.350 4.000 906.010 4.280 ;
        RECT 906.850 4.000 917.510 4.280 ;
        RECT 918.350 4.000 929.010 4.280 ;
        RECT 929.850 4.000 940.970 4.280 ;
        RECT 941.810 4.000 952.470 4.280 ;
        RECT 953.310 4.000 963.970 4.280 ;
        RECT 964.810 4.000 975.470 4.280 ;
        RECT 976.310 4.000 986.970 4.280 ;
        RECT 987.810 4.000 998.470 4.280 ;
        RECT 999.310 4.000 1009.970 4.280 ;
        RECT 1010.810 4.000 1021.470 4.280 ;
        RECT 1022.310 4.000 1032.970 4.280 ;
        RECT 1033.810 4.000 1044.930 4.280 ;
        RECT 1045.770 4.000 1056.430 4.280 ;
        RECT 1057.270 4.000 1067.930 4.280 ;
        RECT 1068.770 4.000 1079.430 4.280 ;
        RECT 1080.270 4.000 1090.930 4.280 ;
        RECT 1091.770 4.000 1102.430 4.280 ;
        RECT 1103.270 4.000 1113.930 4.280 ;
        RECT 1114.770 4.000 1125.430 4.280 ;
        RECT 1126.270 4.000 1136.930 4.280 ;
        RECT 1137.770 4.000 1148.890 4.280 ;
        RECT 1149.730 4.000 1160.390 4.280 ;
        RECT 1161.230 4.000 1171.890 4.280 ;
        RECT 1172.730 4.000 1183.390 4.280 ;
        RECT 1184.230 4.000 1194.890 4.280 ;
        RECT 1195.730 4.000 1206.390 4.280 ;
        RECT 1207.230 4.000 1217.890 4.280 ;
        RECT 1218.730 4.000 1229.390 4.280 ;
        RECT 1230.230 4.000 1240.890 4.280 ;
        RECT 1241.730 4.000 1252.850 4.280 ;
        RECT 1253.690 4.000 1264.350 4.280 ;
        RECT 1265.190 4.000 1275.850 4.280 ;
        RECT 1276.690 4.000 1287.350 4.280 ;
        RECT 1288.190 4.000 1298.850 4.280 ;
        RECT 1299.690 4.000 1310.350 4.280 ;
        RECT 1311.190 4.000 1321.850 4.280 ;
        RECT 1322.690 4.000 1333.350 4.280 ;
        RECT 1334.190 4.000 1344.850 4.280 ;
        RECT 1345.690 4.000 1356.810 4.280 ;
        RECT 1357.650 4.000 1368.310 4.280 ;
        RECT 1369.150 4.000 1379.810 4.280 ;
        RECT 1380.650 4.000 1391.310 4.280 ;
        RECT 1392.150 4.000 1402.810 4.280 ;
        RECT 1403.650 4.000 1414.310 4.280 ;
        RECT 1415.150 4.000 1425.810 4.280 ;
        RECT 1426.650 4.000 1437.310 4.280 ;
        RECT 1438.150 4.000 1448.810 4.280 ;
        RECT 1449.650 4.000 1460.770 4.280 ;
        RECT 1461.610 4.000 1472.270 4.280 ;
        RECT 1473.110 4.000 1483.770 4.280 ;
        RECT 1484.610 4.000 1495.270 4.280 ;
        RECT 1496.110 4.000 1506.770 4.280 ;
        RECT 1507.610 4.000 1518.270 4.280 ;
        RECT 1519.110 4.000 1529.770 4.280 ;
        RECT 1530.610 4.000 1541.270 4.280 ;
        RECT 1542.110 4.000 1552.770 4.280 ;
        RECT 1553.610 4.000 1564.730 4.280 ;
        RECT 1565.570 4.000 1576.230 4.280 ;
        RECT 1577.070 4.000 1587.730 4.280 ;
        RECT 1588.570 4.000 1599.230 4.280 ;
        RECT 1600.070 4.000 1610.730 4.280 ;
        RECT 1611.570 4.000 1622.230 4.280 ;
        RECT 1623.070 4.000 1633.730 4.280 ;
        RECT 1634.570 4.000 1645.230 4.280 ;
        RECT 1646.070 4.000 1656.730 4.280 ;
        RECT 1657.570 4.000 1668.690 4.280 ;
        RECT 1669.530 4.000 1680.190 4.280 ;
        RECT 1681.030 4.000 1691.690 4.280 ;
        RECT 1692.530 4.000 1703.190 4.280 ;
        RECT 1704.030 4.000 1714.690 4.280 ;
        RECT 1715.530 4.000 1726.190 4.280 ;
        RECT 1727.030 4.000 1737.690 4.280 ;
        RECT 1738.530 4.000 1749.190 4.280 ;
        RECT 1750.030 4.000 1760.690 4.280 ;
        RECT 1761.530 4.000 1772.650 4.280 ;
        RECT 1773.490 4.000 1784.150 4.280 ;
        RECT 1784.990 4.000 1795.650 4.280 ;
        RECT 1796.490 4.000 1807.150 4.280 ;
        RECT 1807.990 4.000 1818.650 4.280 ;
        RECT 1819.490 4.000 1830.150 4.280 ;
        RECT 1830.990 4.000 1841.650 4.280 ;
        RECT 1842.490 4.000 1853.150 4.280 ;
        RECT 1853.990 4.000 1864.650 4.280 ;
        RECT 1865.490 4.000 1876.610 4.280 ;
        RECT 1877.450 4.000 1888.110 4.280 ;
        RECT 1888.950 4.000 1899.610 4.280 ;
        RECT 1900.450 4.000 1911.110 4.280 ;
        RECT 1911.950 4.000 1922.610 4.280 ;
        RECT 1923.450 4.000 1934.110 4.280 ;
        RECT 1934.950 4.000 1945.610 4.280 ;
        RECT 1946.450 4.000 1957.110 4.280 ;
        RECT 1957.950 4.000 1968.610 4.280 ;
        RECT 1969.450 4.000 1980.570 4.280 ;
        RECT 1981.410 4.000 1992.070 4.280 ;
        RECT 1992.910 4.000 2003.570 4.280 ;
        RECT 2004.410 4.000 2015.070 4.280 ;
        RECT 2015.910 4.000 2026.570 4.280 ;
        RECT 2027.410 4.000 2038.070 4.280 ;
        RECT 2038.910 4.000 2049.570 4.280 ;
        RECT 2050.410 4.000 2061.070 4.280 ;
        RECT 2061.910 4.000 2072.570 4.280 ;
        RECT 2073.410 4.000 2084.530 4.280 ;
        RECT 2085.370 4.000 2096.030 4.280 ;
        RECT 2096.870 4.000 2107.530 4.280 ;
        RECT 2108.370 4.000 2119.030 4.280 ;
        RECT 2119.870 4.000 2130.530 4.280 ;
        RECT 2131.370 4.000 2142.030 4.280 ;
        RECT 2142.870 4.000 2153.530 4.280 ;
        RECT 2154.370 4.000 2165.030 4.280 ;
        RECT 2165.870 4.000 2176.530 4.280 ;
        RECT 2177.370 4.000 2188.490 4.280 ;
        RECT 2189.330 4.000 2199.990 4.280 ;
        RECT 2200.830 4.000 2211.490 4.280 ;
        RECT 2212.330 4.000 2222.990 4.280 ;
        RECT 2223.830 4.000 2234.490 4.280 ;
        RECT 2235.330 4.000 2245.990 4.280 ;
        RECT 2246.830 4.000 2257.490 4.280 ;
        RECT 2258.330 4.000 2268.990 4.280 ;
        RECT 2269.830 4.000 2280.490 4.280 ;
        RECT 2281.330 4.000 2292.450 4.280 ;
        RECT 2293.290 4.000 2303.950 4.280 ;
        RECT 2304.790 4.000 2315.450 4.280 ;
        RECT 2316.290 4.000 2326.950 4.280 ;
        RECT 2327.790 4.000 2338.450 4.280 ;
        RECT 2339.290 4.000 2349.950 4.280 ;
        RECT 2350.790 4.000 2361.450 4.280 ;
        RECT 2362.290 4.000 2372.950 4.280 ;
        RECT 2373.790 4.000 2384.450 4.280 ;
        RECT 2385.290 4.000 2396.410 4.280 ;
        RECT 2397.250 4.000 2407.910 4.280 ;
        RECT 2408.750 4.000 2419.410 4.280 ;
        RECT 2420.250 4.000 2430.910 4.280 ;
        RECT 2431.750 4.000 2442.410 4.280 ;
        RECT 2443.250 4.000 2453.910 4.280 ;
        RECT 2454.750 4.000 2465.410 4.280 ;
        RECT 2466.250 4.000 2476.910 4.280 ;
        RECT 2477.750 4.000 2488.410 4.280 ;
      LAYER met3 ;
        RECT 4.000 2815.560 2491.000 2850.285 ;
        RECT 4.400 2814.160 2491.000 2815.560 ;
        RECT 4.000 2805.360 2491.000 2814.160 ;
        RECT 4.000 2803.960 2490.600 2805.360 ;
        RECT 4.000 2716.960 2491.000 2803.960 ;
        RECT 4.400 2715.560 2491.000 2716.960 ;
        RECT 4.000 2685.680 2491.000 2715.560 ;
        RECT 4.000 2684.280 2490.600 2685.680 ;
        RECT 4.000 2618.360 2491.000 2684.280 ;
        RECT 4.400 2616.960 2491.000 2618.360 ;
        RECT 4.000 2566.680 2491.000 2616.960 ;
        RECT 4.000 2565.280 2490.600 2566.680 ;
        RECT 4.000 2519.080 2491.000 2565.280 ;
        RECT 4.400 2517.680 2491.000 2519.080 ;
        RECT 4.000 2447.000 2491.000 2517.680 ;
        RECT 4.000 2445.600 2490.600 2447.000 ;
        RECT 4.000 2420.480 2491.000 2445.600 ;
        RECT 4.400 2419.080 2491.000 2420.480 ;
        RECT 4.000 2328.000 2491.000 2419.080 ;
        RECT 4.000 2326.600 2490.600 2328.000 ;
        RECT 4.000 2321.880 2491.000 2326.600 ;
        RECT 4.400 2320.480 2491.000 2321.880 ;
        RECT 4.000 2223.280 2491.000 2320.480 ;
        RECT 4.400 2221.880 2491.000 2223.280 ;
        RECT 4.000 2208.320 2491.000 2221.880 ;
        RECT 4.000 2206.920 2490.600 2208.320 ;
        RECT 4.000 2124.000 2491.000 2206.920 ;
        RECT 4.400 2122.600 2491.000 2124.000 ;
        RECT 4.000 2089.320 2491.000 2122.600 ;
        RECT 4.000 2087.920 2490.600 2089.320 ;
        RECT 4.000 2025.400 2491.000 2087.920 ;
        RECT 4.400 2024.000 2491.000 2025.400 ;
        RECT 4.000 1969.640 2491.000 2024.000 ;
        RECT 4.000 1968.240 2490.600 1969.640 ;
        RECT 4.000 1926.800 2491.000 1968.240 ;
        RECT 4.400 1925.400 2491.000 1926.800 ;
        RECT 4.000 1850.640 2491.000 1925.400 ;
        RECT 4.000 1849.240 2490.600 1850.640 ;
        RECT 4.000 1827.520 2491.000 1849.240 ;
        RECT 4.400 1826.120 2491.000 1827.520 ;
        RECT 4.000 1730.960 2491.000 1826.120 ;
        RECT 4.000 1729.560 2490.600 1730.960 ;
        RECT 4.000 1728.920 2491.000 1729.560 ;
        RECT 4.400 1727.520 2491.000 1728.920 ;
        RECT 4.000 1630.320 2491.000 1727.520 ;
        RECT 4.400 1628.920 2491.000 1630.320 ;
        RECT 4.000 1611.960 2491.000 1628.920 ;
        RECT 4.000 1610.560 2490.600 1611.960 ;
        RECT 4.000 1531.720 2491.000 1610.560 ;
        RECT 4.400 1530.320 2491.000 1531.720 ;
        RECT 4.000 1492.280 2491.000 1530.320 ;
        RECT 4.000 1490.880 2490.600 1492.280 ;
        RECT 4.000 1432.440 2491.000 1490.880 ;
        RECT 4.400 1431.040 2491.000 1432.440 ;
        RECT 4.000 1372.600 2491.000 1431.040 ;
        RECT 4.000 1371.200 2490.600 1372.600 ;
        RECT 4.000 1333.840 2491.000 1371.200 ;
        RECT 4.400 1332.440 2491.000 1333.840 ;
        RECT 4.000 1253.600 2491.000 1332.440 ;
        RECT 4.000 1252.200 2490.600 1253.600 ;
        RECT 4.000 1235.240 2491.000 1252.200 ;
        RECT 4.400 1233.840 2491.000 1235.240 ;
        RECT 4.000 1136.640 2491.000 1233.840 ;
        RECT 4.400 1135.240 2491.000 1136.640 ;
        RECT 4.000 1133.920 2491.000 1135.240 ;
        RECT 4.000 1132.520 2490.600 1133.920 ;
        RECT 4.000 1037.360 2491.000 1132.520 ;
        RECT 4.400 1035.960 2491.000 1037.360 ;
        RECT 4.000 1014.920 2491.000 1035.960 ;
        RECT 4.000 1013.520 2490.600 1014.920 ;
        RECT 4.000 938.760 2491.000 1013.520 ;
        RECT 4.400 937.360 2491.000 938.760 ;
        RECT 4.000 895.240 2491.000 937.360 ;
        RECT 4.000 893.840 2490.600 895.240 ;
        RECT 4.000 840.160 2491.000 893.840 ;
        RECT 4.400 838.760 2491.000 840.160 ;
        RECT 4.000 776.240 2491.000 838.760 ;
        RECT 4.000 774.840 2490.600 776.240 ;
        RECT 4.000 740.880 2491.000 774.840 ;
        RECT 4.400 739.480 2491.000 740.880 ;
        RECT 4.000 656.560 2491.000 739.480 ;
        RECT 4.000 655.160 2490.600 656.560 ;
        RECT 4.000 642.280 2491.000 655.160 ;
        RECT 4.400 640.880 2491.000 642.280 ;
        RECT 4.000 543.680 2491.000 640.880 ;
        RECT 4.400 542.280 2491.000 543.680 ;
        RECT 4.000 537.560 2491.000 542.280 ;
        RECT 4.000 536.160 2490.600 537.560 ;
        RECT 4.000 445.080 2491.000 536.160 ;
        RECT 4.400 443.680 2491.000 445.080 ;
        RECT 4.000 417.880 2491.000 443.680 ;
        RECT 4.000 416.480 2490.600 417.880 ;
        RECT 4.000 345.800 2491.000 416.480 ;
        RECT 4.400 344.400 2491.000 345.800 ;
        RECT 4.000 298.880 2491.000 344.400 ;
        RECT 4.000 297.480 2490.600 298.880 ;
        RECT 4.000 247.200 2491.000 297.480 ;
        RECT 4.400 245.800 2491.000 247.200 ;
        RECT 4.000 179.200 2491.000 245.800 ;
        RECT 4.000 177.800 2490.600 179.200 ;
        RECT 4.000 148.600 2491.000 177.800 ;
        RECT 4.400 147.200 2491.000 148.600 ;
        RECT 4.000 60.200 2491.000 147.200 ;
        RECT 4.000 58.800 2490.600 60.200 ;
        RECT 4.000 50.000 2491.000 58.800 ;
        RECT 4.400 48.600 2491.000 50.000 ;
        RECT 4.000 4.255 2491.000 48.600 ;
      LAYER met4 ;
        RECT 61.935 17.175 2443.225 2850.360 ;
      LAYER met5 ;
        RECT 72.045 2826.480 2422.955 2842.780 ;
        RECT 72.045 2803.980 2422.955 2820.280 ;
        RECT 72.045 2781.480 2422.955 2797.780 ;
        RECT 72.045 2758.980 2422.955 2775.280 ;
        RECT 72.045 2736.480 2422.955 2752.780 ;
        RECT 72.045 2713.980 2422.955 2730.280 ;
        RECT 72.045 2691.480 2422.955 2707.780 ;
        RECT 72.045 2668.980 2422.955 2685.280 ;
        RECT 72.045 2646.480 2422.955 2662.780 ;
        RECT 72.045 2623.980 2422.955 2640.280 ;
        RECT 72.045 2601.480 2422.955 2617.780 ;
        RECT 72.045 2578.980 2422.955 2595.280 ;
        RECT 72.045 2556.480 2422.955 2572.780 ;
        RECT 72.045 2533.980 2422.955 2550.280 ;
        RECT 72.045 2511.480 2422.955 2527.780 ;
        RECT 72.045 2488.980 2422.955 2505.280 ;
        RECT 72.045 2466.480 2422.955 2482.780 ;
        RECT 72.045 2443.980 2422.955 2460.280 ;
        RECT 72.045 2421.480 2422.955 2437.780 ;
        RECT 72.045 2398.980 2422.955 2415.280 ;
        RECT 72.045 2376.480 2422.955 2392.780 ;
        RECT 72.045 2353.980 2422.955 2370.280 ;
        RECT 72.045 2331.480 2422.955 2347.780 ;
        RECT 72.045 2308.980 2422.955 2325.280 ;
        RECT 72.045 2286.480 2422.955 2302.780 ;
        RECT 72.045 2263.980 2422.955 2280.280 ;
        RECT 72.045 2241.480 2422.955 2257.780 ;
        RECT 72.045 2218.980 2422.955 2235.280 ;
        RECT 72.045 2196.480 2422.955 2212.780 ;
        RECT 72.045 2173.980 2422.955 2190.280 ;
        RECT 72.045 2151.480 2422.955 2167.780 ;
        RECT 72.045 2128.980 2422.955 2145.280 ;
        RECT 72.045 2106.480 2422.955 2122.780 ;
        RECT 72.045 2083.980 2422.955 2100.280 ;
        RECT 72.045 2061.480 2422.955 2077.780 ;
        RECT 72.045 2038.980 2422.955 2055.280 ;
        RECT 72.045 2016.480 2422.955 2032.780 ;
        RECT 72.045 1993.980 2422.955 2010.280 ;
        RECT 72.045 1971.480 2422.955 1987.780 ;
        RECT 72.045 1948.980 2422.955 1965.280 ;
        RECT 72.045 1926.480 2422.955 1942.780 ;
        RECT 72.045 1903.980 2422.955 1920.280 ;
        RECT 72.045 1881.480 2422.955 1897.780 ;
        RECT 72.045 1858.980 2422.955 1875.280 ;
        RECT 72.045 1836.480 2422.955 1852.780 ;
        RECT 72.045 1813.980 2422.955 1830.280 ;
        RECT 72.045 1791.480 2422.955 1807.780 ;
        RECT 72.045 1768.980 2422.955 1785.280 ;
        RECT 72.045 1746.480 2422.955 1762.780 ;
        RECT 72.045 1723.980 2422.955 1740.280 ;
        RECT 72.045 1701.480 2422.955 1717.780 ;
        RECT 72.045 1678.980 2422.955 1695.280 ;
        RECT 72.045 1656.480 2422.955 1672.780 ;
        RECT 72.045 1633.980 2422.955 1650.280 ;
        RECT 72.045 1611.480 2422.955 1627.780 ;
        RECT 72.045 1588.980 2422.955 1605.280 ;
        RECT 72.045 1566.480 2422.955 1582.780 ;
        RECT 72.045 1543.980 2422.955 1560.280 ;
        RECT 72.045 1521.480 2422.955 1537.780 ;
        RECT 72.045 1498.980 2422.955 1515.280 ;
        RECT 72.045 1476.480 2422.955 1492.780 ;
        RECT 72.045 1453.980 2422.955 1470.280 ;
        RECT 72.045 1431.480 2422.955 1447.780 ;
        RECT 72.045 1408.980 2422.955 1425.280 ;
        RECT 72.045 1386.480 2422.955 1402.780 ;
        RECT 72.045 1363.980 2422.955 1380.280 ;
        RECT 72.045 1341.480 2422.955 1357.780 ;
        RECT 72.045 1318.980 2422.955 1335.280 ;
        RECT 72.045 1296.480 2422.955 1312.780 ;
        RECT 72.045 1273.980 2422.955 1290.280 ;
        RECT 72.045 1251.480 2422.955 1267.780 ;
        RECT 72.045 1228.980 2422.955 1245.280 ;
        RECT 72.045 1206.480 2422.955 1222.780 ;
        RECT 72.045 1183.980 2422.955 1200.280 ;
        RECT 72.045 1161.480 2422.955 1177.780 ;
        RECT 72.045 1138.980 2422.955 1155.280 ;
        RECT 72.045 1116.480 2422.955 1132.780 ;
        RECT 72.045 1093.980 2422.955 1110.280 ;
        RECT 72.045 1071.480 2422.955 1087.780 ;
        RECT 72.045 1048.980 2422.955 1065.280 ;
        RECT 72.045 1026.480 2422.955 1042.780 ;
        RECT 72.045 1003.980 2422.955 1020.280 ;
        RECT 72.045 981.480 2422.955 997.780 ;
        RECT 72.045 958.980 2422.955 975.280 ;
        RECT 72.045 936.480 2422.955 952.780 ;
        RECT 72.045 913.980 2422.955 930.280 ;
        RECT 72.045 891.480 2422.955 907.780 ;
        RECT 72.045 868.980 2422.955 885.280 ;
        RECT 72.045 846.480 2422.955 862.780 ;
        RECT 72.045 823.980 2422.955 840.280 ;
        RECT 72.045 801.480 2422.955 817.780 ;
        RECT 72.045 778.980 2422.955 795.280 ;
        RECT 72.045 756.480 2422.955 772.780 ;
        RECT 72.045 733.980 2422.955 750.280 ;
        RECT 72.045 711.480 2422.955 727.780 ;
        RECT 72.045 688.980 2422.955 705.280 ;
        RECT 72.045 666.480 2422.955 682.780 ;
        RECT 72.045 643.980 2422.955 660.280 ;
        RECT 72.045 621.480 2422.955 637.780 ;
        RECT 72.045 598.980 2422.955 615.280 ;
        RECT 72.045 576.480 2422.955 592.780 ;
        RECT 72.045 553.980 2422.955 570.280 ;
        RECT 72.045 531.480 2422.955 547.780 ;
        RECT 72.045 508.980 2422.955 525.280 ;
        RECT 72.045 486.480 2422.955 502.780 ;
        RECT 72.045 463.980 2422.955 480.280 ;
        RECT 72.045 441.480 2422.955 457.780 ;
        RECT 72.045 418.980 2422.955 435.280 ;
        RECT 72.045 396.480 2422.955 412.780 ;
        RECT 72.045 373.980 2422.955 390.280 ;
        RECT 72.045 351.480 2422.955 367.780 ;
        RECT 72.045 328.980 2422.955 345.280 ;
        RECT 72.045 306.480 2422.955 322.780 ;
        RECT 72.045 283.980 2422.955 300.280 ;
        RECT 72.045 261.480 2422.955 277.780 ;
        RECT 72.045 238.980 2422.955 255.280 ;
        RECT 72.045 216.480 2422.955 232.780 ;
        RECT 72.045 193.980 2422.955 210.280 ;
        RECT 72.045 171.480 2422.955 187.780 ;
        RECT 72.045 148.980 2422.955 165.280 ;
        RECT 72.045 126.480 2422.955 142.780 ;
        RECT 72.045 103.980 2422.955 120.280 ;
  END
END fpga_core
END LIBRARY

