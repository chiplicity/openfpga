magic
tech sky130A
magscale 1 2
timestamp 1609023970
<< locali >>
rect 8309 14331 8343 14501
rect 6561 13243 6595 13481
rect 9505 13175 9539 13481
rect 9505 10115 9539 10217
rect 16129 10115 16163 10965
rect 9505 5559 9539 5797
rect 12909 2839 12943 3077
<< viali >>
rect 1777 17289 1811 17323
rect 7297 17289 7331 17323
rect 8125 17289 8159 17323
rect 8401 17289 8435 17323
rect 14381 17289 14415 17323
rect 14565 17221 14599 17255
rect 9505 17153 9539 17187
rect 10609 17153 10643 17187
rect 11437 17153 11471 17187
rect 1593 17085 1627 17119
rect 2053 17085 2087 17119
rect 7113 17085 7147 17119
rect 7941 17085 7975 17119
rect 12633 17085 12667 17119
rect 14933 17085 14967 17119
rect 3617 17017 3651 17051
rect 7481 17017 7515 17051
rect 10425 17017 10459 17051
rect 11253 17017 11287 17051
rect 12900 17017 12934 17051
rect 3157 16949 3191 16983
rect 6009 16949 6043 16983
rect 6929 16949 6963 16983
rect 7665 16949 7699 16983
rect 9229 16949 9263 16983
rect 9873 16949 9907 16983
rect 10057 16949 10091 16983
rect 10517 16949 10551 16983
rect 10885 16949 10919 16983
rect 11345 16949 11379 16983
rect 14013 16949 14047 16983
rect 15025 16949 15059 16983
rect 2605 16745 2639 16779
rect 2973 16745 3007 16779
rect 3709 16745 3743 16779
rect 4721 16745 4755 16779
rect 5457 16745 5491 16779
rect 6193 16745 6227 16779
rect 6561 16745 6595 16779
rect 6929 16745 6963 16779
rect 9413 16745 9447 16779
rect 10149 16745 10183 16779
rect 10885 16745 10919 16779
rect 12449 16745 12483 16779
rect 12817 16745 12851 16779
rect 1777 16677 1811 16711
rect 7205 16677 7239 16711
rect 10057 16677 10091 16711
rect 10701 16677 10735 16711
rect 11314 16677 11348 16711
rect 13185 16677 13219 16711
rect 13912 16677 13946 16711
rect 1501 16609 1535 16643
rect 2053 16609 2087 16643
rect 2421 16609 2455 16643
rect 2789 16609 2823 16643
rect 3157 16609 3191 16643
rect 3525 16609 3559 16643
rect 4077 16609 4111 16643
rect 4537 16609 4571 16643
rect 4905 16609 4939 16643
rect 5273 16609 5307 16643
rect 5641 16609 5675 16643
rect 6009 16609 6043 16643
rect 6377 16609 6411 16643
rect 6745 16609 6779 16643
rect 7656 16609 7690 16643
rect 8861 16609 8895 16643
rect 9229 16609 9263 16643
rect 11069 16609 11103 16643
rect 13277 16609 13311 16643
rect 7389 16541 7423 16575
rect 10241 16541 10275 16575
rect 13461 16541 13495 16575
rect 13645 16541 13679 16575
rect 2237 16473 2271 16507
rect 3341 16473 3375 16507
rect 4261 16473 4295 16507
rect 5089 16473 5123 16507
rect 5825 16473 5859 16507
rect 8769 16473 8803 16507
rect 9045 16405 9079 16439
rect 9689 16405 9723 16439
rect 10517 16405 10551 16439
rect 15025 16405 15059 16439
rect 3433 16201 3467 16235
rect 8217 16201 8251 16235
rect 10149 16201 10183 16235
rect 12173 16201 12207 16235
rect 12449 16201 12483 16235
rect 13737 16201 13771 16235
rect 5733 16133 5767 16167
rect 13553 16133 13587 16167
rect 1685 16065 1719 16099
rect 6561 16065 6595 16099
rect 8677 16065 8711 16099
rect 10701 16065 10735 16099
rect 10793 16065 10827 16099
rect 11621 16065 11655 16099
rect 13001 16065 13035 16099
rect 14289 16065 14323 16099
rect 14657 16065 14691 16099
rect 15669 16065 15703 16099
rect 1501 15997 1535 16031
rect 3249 15997 3283 16031
rect 3617 15997 3651 16031
rect 6837 15997 6871 16031
rect 8769 15997 8803 16031
rect 7104 15929 7138 15963
rect 8493 15929 8527 15963
rect 9014 15929 9048 15963
rect 11437 15929 11471 15963
rect 11897 15929 11931 15963
rect 12817 15929 12851 15963
rect 12909 15929 12943 15963
rect 13369 15929 13403 15963
rect 14749 15929 14783 15963
rect 2513 15861 2547 15895
rect 2881 15861 2915 15895
rect 3893 15861 3927 15895
rect 4537 15861 4571 15895
rect 4905 15861 4939 15895
rect 5365 15861 5399 15895
rect 5917 15861 5951 15895
rect 6285 15861 6319 15895
rect 6377 15861 6411 15895
rect 10241 15861 10275 15895
rect 10609 15861 10643 15895
rect 11069 15861 11103 15895
rect 11529 15861 11563 15895
rect 14105 15861 14139 15895
rect 14197 15861 14231 15895
rect 7205 15657 7239 15691
rect 8033 15657 8067 15691
rect 8493 15657 8527 15691
rect 10149 15657 10183 15691
rect 10517 15657 10551 15691
rect 10885 15657 10919 15691
rect 11345 15657 11379 15691
rect 11805 15657 11839 15691
rect 12449 15657 12483 15691
rect 14381 15657 14415 15691
rect 15301 15657 15335 15691
rect 1777 15589 1811 15623
rect 3525 15589 3559 15623
rect 8401 15589 8435 15623
rect 10977 15589 11011 15623
rect 1501 15521 1535 15555
rect 3617 15521 3651 15555
rect 5540 15521 5574 15555
rect 7573 15521 7607 15555
rect 7665 15521 7699 15555
rect 10057 15521 10091 15555
rect 11713 15521 11747 15555
rect 12909 15521 12943 15555
rect 13176 15521 13210 15555
rect 14749 15521 14783 15555
rect 3801 15453 3835 15487
rect 5273 15453 5307 15487
rect 7849 15453 7883 15487
rect 8585 15453 8619 15487
rect 8861 15453 8895 15487
rect 10241 15453 10275 15487
rect 11069 15453 11103 15487
rect 11897 15453 11931 15487
rect 12265 15453 12299 15487
rect 14841 15453 14875 15487
rect 14933 15453 14967 15487
rect 6653 15385 6687 15419
rect 9689 15385 9723 15419
rect 14289 15385 14323 15419
rect 3157 15317 3191 15351
rect 9137 15317 9171 15351
rect 9413 15317 9447 15351
rect 2145 15113 2179 15147
rect 4169 15113 4203 15147
rect 6929 15113 6963 15147
rect 11621 15113 11655 15147
rect 13277 15113 13311 15147
rect 14197 15113 14231 15147
rect 1777 15045 1811 15079
rect 5273 15045 5307 15079
rect 7573 15045 7607 15079
rect 2329 14977 2363 15011
rect 4721 14977 4755 15011
rect 5549 14977 5583 15011
rect 8125 14977 8159 15011
rect 8953 14977 8987 15011
rect 9781 14977 9815 15011
rect 13093 14977 13127 15011
rect 13829 14977 13863 15011
rect 14841 14977 14875 15011
rect 15025 14977 15059 15011
rect 1593 14909 1627 14943
rect 1961 14909 1995 14943
rect 2697 14909 2731 14943
rect 4537 14909 4571 14943
rect 5457 14909 5491 14943
rect 7941 14909 7975 14943
rect 9597 14909 9631 14943
rect 10241 14909 10275 14943
rect 10508 14909 10542 14943
rect 11897 14909 11931 14943
rect 12909 14909 12943 14943
rect 2605 14841 2639 14875
rect 2964 14841 2998 14875
rect 4629 14841 4663 14875
rect 5733 14841 5767 14875
rect 7205 14841 7239 14875
rect 8033 14841 8067 14875
rect 9689 14841 9723 14875
rect 12173 14841 12207 14875
rect 13645 14841 13679 14875
rect 14565 14841 14599 14875
rect 15301 14841 15335 14875
rect 4077 14773 4111 14807
rect 4997 14773 5031 14807
rect 7389 14773 7423 14807
rect 8401 14773 8435 14807
rect 8769 14773 8803 14807
rect 8861 14773 8895 14807
rect 9229 14773 9263 14807
rect 10149 14773 10183 14807
rect 11713 14773 11747 14807
rect 12449 14773 12483 14807
rect 12817 14773 12851 14807
rect 13737 14773 13771 14807
rect 14657 14773 14691 14807
rect 15485 14773 15519 14807
rect 3065 14569 3099 14603
rect 6009 14569 6043 14603
rect 6929 14569 6963 14603
rect 7481 14569 7515 14603
rect 7849 14569 7883 14603
rect 13553 14569 13587 14603
rect 8309 14501 8343 14535
rect 11406 14501 11440 14535
rect 13093 14501 13127 14535
rect 14197 14501 14231 14535
rect 1685 14433 1719 14467
rect 1952 14433 1986 14467
rect 3525 14433 3559 14467
rect 4436 14433 4470 14467
rect 6101 14433 6135 14467
rect 6837 14433 6871 14467
rect 7941 14433 7975 14467
rect 3617 14365 3651 14399
rect 3801 14365 3835 14399
rect 4169 14365 4203 14399
rect 6193 14365 6227 14399
rect 7021 14365 7055 14399
rect 8125 14365 8159 14399
rect 8769 14433 8803 14467
rect 9689 14433 9723 14467
rect 9956 14433 9990 14467
rect 11161 14433 11195 14467
rect 13185 14433 13219 14467
rect 13737 14433 13771 14467
rect 8861 14365 8895 14399
rect 9045 14365 9079 14399
rect 13277 14365 13311 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 3157 14297 3191 14331
rect 5549 14297 5583 14331
rect 8309 14297 8343 14331
rect 8401 14297 8435 14331
rect 9321 14297 9355 14331
rect 9505 14297 9539 14331
rect 12541 14297 12575 14331
rect 5641 14229 5675 14263
rect 6469 14229 6503 14263
rect 7297 14229 7331 14263
rect 11069 14229 11103 14263
rect 12725 14229 12759 14263
rect 15393 14229 15427 14263
rect 3157 14025 3191 14059
rect 3985 14025 4019 14059
rect 4813 14025 4847 14059
rect 9781 14025 9815 14059
rect 15071 14025 15105 14059
rect 14749 13957 14783 13991
rect 1685 13889 1719 13923
rect 2789 13889 2823 13923
rect 2973 13889 3007 13923
rect 3801 13889 3835 13923
rect 4629 13889 4663 13923
rect 5273 13889 5307 13923
rect 5457 13889 5491 13923
rect 6193 13889 6227 13923
rect 11989 13889 12023 13923
rect 13093 13889 13127 13923
rect 1501 13821 1535 13855
rect 3617 13821 3651 13855
rect 4353 13821 4387 13855
rect 6101 13821 6135 13855
rect 6469 13821 6503 13855
rect 6837 13821 6871 13855
rect 7093 13821 7127 13855
rect 8401 13821 8435 13855
rect 8668 13821 8702 13855
rect 12265 13821 12299 13855
rect 13001 13821 13035 13855
rect 13369 13821 13403 13855
rect 13625 13821 13659 13855
rect 15000 13821 15034 13855
rect 2697 13753 2731 13787
rect 5181 13753 5215 13787
rect 12909 13753 12943 13787
rect 2329 13685 2363 13719
rect 3525 13685 3559 13719
rect 4445 13685 4479 13719
rect 5641 13685 5675 13719
rect 6009 13685 6043 13719
rect 8217 13685 8251 13719
rect 12541 13685 12575 13719
rect 2881 13481 2915 13515
rect 5641 13481 5675 13515
rect 6561 13481 6595 13515
rect 8953 13481 8987 13515
rect 9505 13481 9539 13515
rect 11437 13481 11471 13515
rect 13277 13481 13311 13515
rect 13369 13481 13403 13515
rect 3249 13413 3283 13447
rect 3801 13413 3835 13447
rect 4905 13413 4939 13447
rect 1501 13345 1535 13379
rect 5549 13345 5583 13379
rect 1685 13277 1719 13311
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 4353 13277 4387 13311
rect 5825 13277 5859 13311
rect 6745 13413 6779 13447
rect 7840 13345 7874 13379
rect 7573 13277 7607 13311
rect 9229 13277 9263 13311
rect 4077 13209 4111 13243
rect 6561 13209 6595 13243
rect 11713 13413 11747 13447
rect 12449 13413 12483 13447
rect 12541 13413 12575 13447
rect 9873 13345 9907 13379
rect 10057 13345 10091 13379
rect 10324 13345 10358 13379
rect 11897 13277 11931 13311
rect 12725 13277 12759 13311
rect 13553 13277 13587 13311
rect 12081 13209 12115 13243
rect 12909 13209 12943 13243
rect 5181 13141 5215 13175
rect 7297 13141 7331 13175
rect 7481 13141 7515 13175
rect 9045 13141 9079 13175
rect 9505 13141 9539 13175
rect 9689 13141 9723 13175
rect 2421 12937 2455 12971
rect 5365 12937 5399 12971
rect 6561 12937 6595 12971
rect 8585 12937 8619 12971
rect 11069 12937 11103 12971
rect 13553 12937 13587 12971
rect 6193 12869 6227 12903
rect 1685 12801 1719 12835
rect 3065 12801 3099 12835
rect 5825 12801 5859 12835
rect 6009 12801 6043 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 8217 12801 8251 12835
rect 9137 12801 9171 12835
rect 10057 12801 10091 12835
rect 10885 12801 10919 12835
rect 11621 12801 11655 12835
rect 13001 12801 13035 12835
rect 15301 12801 15335 12835
rect 1501 12733 1535 12767
rect 2789 12733 2823 12767
rect 3249 12733 3283 12767
rect 6377 12733 6411 12767
rect 9781 12733 9815 12767
rect 11437 12733 11471 12767
rect 12909 12733 12943 12767
rect 15025 12733 15059 12767
rect 3516 12665 3550 12699
rect 8953 12665 8987 12699
rect 11529 12665 11563 12699
rect 12817 12665 12851 12699
rect 13277 12665 13311 12699
rect 2881 12597 2915 12631
rect 4629 12597 4663 12631
rect 5733 12597 5767 12631
rect 6837 12597 6871 12631
rect 7205 12597 7239 12631
rect 7665 12597 7699 12631
rect 8033 12597 8067 12631
rect 8125 12597 8159 12631
rect 9045 12597 9079 12631
rect 9413 12597 9447 12631
rect 9873 12597 9907 12631
rect 10241 12597 10275 12631
rect 10609 12597 10643 12631
rect 10701 12597 10735 12631
rect 11897 12597 11931 12631
rect 12449 12597 12483 12631
rect 14841 12597 14875 12631
rect 3617 12393 3651 12427
rect 9873 12393 9907 12427
rect 12081 12393 12115 12427
rect 5080 12325 5114 12359
rect 10241 12325 10275 12359
rect 12633 12325 12667 12359
rect 1501 12257 1535 12291
rect 2145 12257 2179 12291
rect 2412 12257 2446 12291
rect 4629 12257 4663 12291
rect 6552 12257 6586 12291
rect 7757 12257 7791 12291
rect 8013 12257 8047 12291
rect 10701 12257 10735 12291
rect 10968 12257 11002 12291
rect 13093 12257 13127 12291
rect 1685 12189 1719 12223
rect 4813 12189 4847 12223
rect 6285 12189 6319 12223
rect 10333 12189 10367 12223
rect 10517 12189 10551 12223
rect 12173 12189 12207 12223
rect 13277 12189 13311 12223
rect 3525 12121 3559 12155
rect 6193 12121 6227 12155
rect 9137 12121 9171 12155
rect 3893 12053 3927 12087
rect 4445 12053 4479 12087
rect 7665 12053 7699 12087
rect 9505 12053 9539 12087
rect 12449 12053 12483 12087
rect 2789 11849 2823 11883
rect 4077 11849 4111 11883
rect 4997 11849 5031 11883
rect 7941 11849 7975 11883
rect 9689 11849 9723 11883
rect 10609 11849 10643 11883
rect 11713 11849 11747 11883
rect 12449 11849 12483 11883
rect 13553 11849 13587 11883
rect 9781 11781 9815 11815
rect 4721 11713 4755 11747
rect 5457 11713 5491 11747
rect 5641 11713 5675 11747
rect 6377 11713 6411 11747
rect 7297 11713 7331 11747
rect 7389 11713 7423 11747
rect 7665 11713 7699 11747
rect 9229 11713 9263 11747
rect 10241 11713 10275 11747
rect 10425 11713 10459 11747
rect 11161 11713 11195 11747
rect 13001 11713 13035 11747
rect 1409 11645 1443 11679
rect 5365 11645 5399 11679
rect 7205 11645 7239 11679
rect 8125 11645 8159 11679
rect 11069 11645 11103 11679
rect 11621 11645 11655 11679
rect 12817 11645 12851 11679
rect 1676 11577 1710 11611
rect 4537 11577 4571 11611
rect 6193 11577 6227 11611
rect 9045 11577 9079 11611
rect 10977 11577 11011 11611
rect 4169 11509 4203 11543
rect 4629 11509 4663 11543
rect 5825 11509 5859 11543
rect 6285 11509 6319 11543
rect 6837 11509 6871 11543
rect 8677 11509 8711 11543
rect 9137 11509 9171 11543
rect 10149 11509 10183 11543
rect 11437 11509 11471 11543
rect 12909 11509 12943 11543
rect 13369 11509 13403 11543
rect 2053 11305 2087 11339
rect 2421 11305 2455 11339
rect 5457 11305 5491 11339
rect 5641 11305 5675 11339
rect 7573 11305 7607 11339
rect 8309 11305 8343 11339
rect 10517 11305 10551 11339
rect 11437 11305 11471 11339
rect 3525 11237 3559 11271
rect 8401 11237 8435 11271
rect 11253 11237 11287 11271
rect 4344 11169 4378 11203
rect 6009 11169 6043 11203
rect 6276 11169 6310 11203
rect 9137 11169 9171 11203
rect 9229 11169 9263 11203
rect 10609 11169 10643 11203
rect 11713 11169 11747 11203
rect 11980 11169 12014 11203
rect 2513 11101 2547 11135
rect 2697 11101 2731 11135
rect 3617 11101 3651 11135
rect 3801 11101 3835 11135
rect 4077 11101 4111 11135
rect 8493 11101 8527 11135
rect 9413 11101 9447 11135
rect 9965 11101 9999 11135
rect 10701 11101 10735 11135
rect 7389 11033 7423 11067
rect 9689 11033 9723 11067
rect 10149 11033 10183 11067
rect 10977 11033 11011 11067
rect 3157 10965 3191 10999
rect 7941 10965 7975 10999
rect 8769 10965 8803 10999
rect 13093 10965 13127 10999
rect 16129 10965 16163 10999
rect 3433 10761 3467 10795
rect 5917 10761 5951 10795
rect 11529 10761 11563 10795
rect 14105 10761 14139 10795
rect 5641 10693 5675 10727
rect 9229 10693 9263 10727
rect 1685 10625 1719 10659
rect 3249 10625 3283 10659
rect 3893 10625 3927 10659
rect 4077 10625 4111 10659
rect 4261 10625 4295 10659
rect 6561 10625 6595 10659
rect 7573 10625 7607 10659
rect 9321 10625 9355 10659
rect 12173 10625 12207 10659
rect 1501 10557 1535 10591
rect 6377 10557 6411 10591
rect 7481 10557 7515 10591
rect 7849 10557 7883 10591
rect 9689 10557 9723 10591
rect 10057 10557 10091 10591
rect 12725 10557 12759 10591
rect 2973 10489 3007 10523
rect 4528 10489 4562 10523
rect 6285 10489 6319 10523
rect 8116 10489 8150 10523
rect 10324 10489 10358 10523
rect 11897 10489 11931 10523
rect 12992 10489 13026 10523
rect 2605 10421 2639 10455
rect 3065 10421 3099 10455
rect 3801 10421 3835 10455
rect 7021 10421 7055 10455
rect 7389 10421 7423 10455
rect 11437 10421 11471 10455
rect 11989 10421 12023 10455
rect 14197 10421 14231 10455
rect 2973 10217 3007 10251
rect 3065 10217 3099 10251
rect 3617 10217 3651 10251
rect 5089 10217 5123 10251
rect 7297 10217 7331 10251
rect 7389 10217 7423 10251
rect 9505 10217 9539 10251
rect 14013 10217 14047 10251
rect 14749 10217 14783 10251
rect 6184 10149 6218 10183
rect 7665 10149 7699 10183
rect 11704 10149 11738 10183
rect 15301 10149 15335 10183
rect 1511 10081 1545 10115
rect 4261 10081 4295 10115
rect 4537 10081 4571 10115
rect 5457 10081 5491 10115
rect 5917 10081 5951 10115
rect 9505 10081 9539 10115
rect 10333 10081 10367 10115
rect 13921 10081 13955 10115
rect 14841 10081 14875 10115
rect 15485 10081 15519 10115
rect 16129 10081 16163 10115
rect 1685 10013 1719 10047
rect 3157 10013 3191 10047
rect 5549 10013 5583 10047
rect 5733 10013 5767 10047
rect 10425 10013 10459 10047
rect 10609 10013 10643 10047
rect 11437 10013 11471 10047
rect 14105 10013 14139 10047
rect 14933 10013 14967 10047
rect 2605 9945 2639 9979
rect 3525 9945 3559 9979
rect 9873 9945 9907 9979
rect 8953 9877 8987 9911
rect 9965 9877 9999 9911
rect 12817 9877 12851 9911
rect 13553 9877 13587 9911
rect 14381 9877 14415 9911
rect 11529 9673 11563 9707
rect 8125 9605 8159 9639
rect 8953 9605 8987 9639
rect 13277 9605 13311 9639
rect 5917 9537 5951 9571
rect 8677 9537 8711 9571
rect 9505 9537 9539 9571
rect 9873 9537 9907 9571
rect 10701 9537 10735 9571
rect 12173 9537 12207 9571
rect 13001 9537 13035 9571
rect 13737 9537 13771 9571
rect 13829 9537 13863 9571
rect 2973 9469 3007 9503
rect 5825 9469 5859 9503
rect 9413 9469 9447 9503
rect 10425 9469 10459 9503
rect 11069 9469 11103 9503
rect 11897 9469 11931 9503
rect 13645 9469 13679 9503
rect 3240 9401 3274 9435
rect 8493 9401 8527 9435
rect 9321 9401 9355 9435
rect 10977 9401 11011 9435
rect 12817 9401 12851 9435
rect 4353 9333 4387 9367
rect 4997 9333 5031 9367
rect 6193 9333 6227 9367
rect 8585 9333 8619 9367
rect 10057 9333 10091 9367
rect 10517 9333 10551 9367
rect 11989 9333 12023 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 14473 9333 14507 9367
rect 7757 9129 7791 9163
rect 8401 9129 8435 9163
rect 8585 9129 8619 9163
rect 9045 9129 9079 9163
rect 9689 9129 9723 9163
rect 10149 9129 10183 9163
rect 10609 9129 10643 9163
rect 12173 9129 12207 9163
rect 12541 9129 12575 9163
rect 13369 9129 13403 9163
rect 4690 9061 4724 9095
rect 10057 9061 10091 9095
rect 10968 9061 11002 9095
rect 4445 8993 4479 9027
rect 5917 8993 5951 9027
rect 6184 8993 6218 9027
rect 7849 8993 7883 9027
rect 8953 8993 8987 9027
rect 9505 8993 9539 9027
rect 12909 8993 12943 9027
rect 13737 8993 13771 9027
rect 14197 8993 14231 9027
rect 7941 8925 7975 8959
rect 9137 8925 9171 8959
rect 10241 8925 10275 8959
rect 10701 8925 10735 8959
rect 12357 8925 12391 8959
rect 13001 8925 13035 8959
rect 13093 8925 13127 8959
rect 13829 8925 13863 8959
rect 13921 8925 13955 8959
rect 7297 8857 7331 8891
rect 12081 8857 12115 8891
rect 5825 8789 5859 8823
rect 7389 8789 7423 8823
rect 8309 8789 8343 8823
rect 11161 8585 11195 8619
rect 11529 8585 11563 8619
rect 14381 8585 14415 8619
rect 5733 8517 5767 8551
rect 2329 8449 2363 8483
rect 3801 8449 3835 8483
rect 4629 8449 4663 8483
rect 5457 8449 5491 8483
rect 6285 8449 6319 8483
rect 6837 8449 6871 8483
rect 8953 8449 8987 8483
rect 12081 8449 12115 8483
rect 13001 8449 13035 8483
rect 1501 8381 1535 8415
rect 2053 8381 2087 8415
rect 3617 8381 3651 8415
rect 5273 8381 5307 8415
rect 6101 8381 6135 8415
rect 6193 8381 6227 8415
rect 7104 8381 7138 8415
rect 8769 8381 8803 8415
rect 9781 8381 9815 8415
rect 11897 8381 11931 8415
rect 12633 8381 12667 8415
rect 13257 8381 13291 8415
rect 1777 8313 1811 8347
rect 4537 8313 4571 8347
rect 5365 8313 5399 8347
rect 10048 8313 10082 8347
rect 11989 8313 12023 8347
rect 12449 8313 12483 8347
rect 3249 8245 3283 8279
rect 3709 8245 3743 8279
rect 4077 8245 4111 8279
rect 4445 8245 4479 8279
rect 4905 8245 4939 8279
rect 6561 8245 6595 8279
rect 8217 8245 8251 8279
rect 8401 8245 8435 8279
rect 8861 8245 8895 8279
rect 9229 8245 9263 8279
rect 9597 8245 9631 8279
rect 11345 8245 11379 8279
rect 2697 8041 2731 8075
rect 3617 8041 3651 8075
rect 4813 8041 4847 8075
rect 5181 8041 5215 8075
rect 5641 8041 5675 8075
rect 6653 8041 6687 8075
rect 7297 8041 7331 8075
rect 8125 8041 8159 8075
rect 8585 8041 8619 8075
rect 8953 8041 8987 8075
rect 9781 8041 9815 8075
rect 10057 8041 10091 8075
rect 11345 8041 11379 8075
rect 12541 8041 12575 8075
rect 3525 7973 3559 8007
rect 5273 7973 5307 8007
rect 6009 7973 6043 8007
rect 12265 7973 12299 8007
rect 1501 7905 1535 7939
rect 4721 7905 4755 7939
rect 7205 7905 7239 7939
rect 9973 7905 10007 7939
rect 10425 7905 10459 7939
rect 11253 7905 11287 7939
rect 11713 7905 11747 7939
rect 12909 7905 12943 7939
rect 1685 7837 1719 7871
rect 2789 7837 2823 7871
rect 2973 7837 3007 7871
rect 3801 7837 3835 7871
rect 5365 7837 5399 7871
rect 6101 7837 6135 7871
rect 6193 7837 6227 7871
rect 7389 7837 7423 7871
rect 8217 7837 8251 7871
rect 8309 7837 8343 7871
rect 9045 7837 9079 7871
rect 9137 7837 9171 7871
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 11437 7837 11471 7871
rect 13001 7837 13035 7871
rect 13093 7837 13127 7871
rect 2329 7769 2363 7803
rect 3157 7769 3191 7803
rect 6837 7769 6871 7803
rect 10885 7769 10919 7803
rect 4537 7701 4571 7735
rect 6561 7701 6595 7735
rect 7757 7701 7791 7735
rect 9505 7701 9539 7735
rect 12357 7701 12391 7735
rect 4813 7497 4847 7531
rect 5089 7497 5123 7531
rect 5641 7497 5675 7531
rect 6561 7497 6595 7531
rect 8953 7497 8987 7531
rect 10609 7497 10643 7531
rect 11437 7497 11471 7531
rect 7021 7429 7055 7463
rect 8861 7429 8895 7463
rect 6193 7361 6227 7395
rect 9413 7361 9447 7395
rect 9505 7361 9539 7395
rect 10333 7361 10367 7395
rect 11161 7361 11195 7395
rect 12081 7361 12115 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 1961 7293 1995 7327
rect 3433 7293 3467 7327
rect 6101 7293 6135 7327
rect 7389 7293 7423 7327
rect 7481 7293 7515 7327
rect 7748 7293 7782 7327
rect 10241 7293 10275 7327
rect 13461 7293 13495 7327
rect 2206 7225 2240 7259
rect 3678 7225 3712 7259
rect 9321 7225 9355 7259
rect 11069 7225 11103 7259
rect 11805 7225 11839 7259
rect 3341 7157 3375 7191
rect 6009 7157 6043 7191
rect 6837 7157 6871 7191
rect 7205 7157 7239 7191
rect 9781 7157 9815 7191
rect 10149 7157 10183 7191
rect 10977 7157 11011 7191
rect 11897 7157 11931 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 13277 7157 13311 7191
rect 1869 6953 1903 6987
rect 2237 6953 2271 6987
rect 4353 6953 4387 6987
rect 4721 6953 4755 6987
rect 5181 6953 5215 6987
rect 8309 6953 8343 6987
rect 11069 6953 11103 6987
rect 12909 6953 12943 6987
rect 1777 6885 1811 6919
rect 6377 6885 6411 6919
rect 7196 6885 7230 6919
rect 9956 6885 9990 6919
rect 2605 6817 2639 6851
rect 2697 6817 2731 6851
rect 5549 6817 5583 6851
rect 5641 6817 5675 6851
rect 6469 6817 6503 6851
rect 6929 6817 6963 6851
rect 11704 6817 11738 6851
rect 13277 6817 13311 6851
rect 13369 6817 13403 6851
rect 13737 6817 13771 6851
rect 2053 6749 2087 6783
rect 2789 6749 2823 6783
rect 4813 6749 4847 6783
rect 4905 6749 4939 6783
rect 5733 6749 5767 6783
rect 6561 6749 6595 6783
rect 9413 6749 9447 6783
rect 9689 6749 9723 6783
rect 11437 6749 11471 6783
rect 13553 6749 13587 6783
rect 6009 6681 6043 6715
rect 9321 6681 9355 6715
rect 1409 6613 1443 6647
rect 11253 6613 11287 6647
rect 12817 6613 12851 6647
rect 2789 6409 2823 6443
rect 4629 6409 4663 6443
rect 5181 6409 5215 6443
rect 6009 6409 6043 6443
rect 6561 6409 6595 6443
rect 9689 6409 9723 6443
rect 9781 6409 9815 6443
rect 10241 6409 10275 6443
rect 10425 6409 10459 6443
rect 6837 6341 6871 6375
rect 1409 6273 1443 6307
rect 5733 6273 5767 6307
rect 6285 6273 6319 6307
rect 10977 6273 11011 6307
rect 12081 6273 12115 6307
rect 1665 6205 1699 6239
rect 3249 6205 3283 6239
rect 5549 6205 5583 6239
rect 6193 6205 6227 6239
rect 7941 6205 7975 6239
rect 8309 6205 8343 6239
rect 8576 6205 8610 6239
rect 9965 6205 9999 6239
rect 3494 6137 3528 6171
rect 10793 6137 10827 6171
rect 5641 6069 5675 6103
rect 7021 6069 7055 6103
rect 7205 6069 7239 6103
rect 10885 6069 10919 6103
rect 11345 6069 11379 6103
rect 2053 5865 2087 5899
rect 2881 5865 2915 5899
rect 3801 5865 3835 5899
rect 5641 5865 5675 5899
rect 6377 5865 6411 5899
rect 1777 5797 1811 5831
rect 2421 5797 2455 5831
rect 8769 5797 8803 5831
rect 9505 5797 9539 5831
rect 9689 5797 9723 5831
rect 9873 5797 9907 5831
rect 10701 5797 10735 5831
rect 14933 5797 14967 5831
rect 1501 5729 1535 5763
rect 3249 5729 3283 5763
rect 4344 5729 4378 5763
rect 6469 5729 6503 5763
rect 7104 5729 7138 5763
rect 8677 5729 8711 5763
rect 9229 5729 9263 5763
rect 2513 5661 2547 5695
rect 2697 5661 2731 5695
rect 3341 5661 3375 5695
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 8861 5661 8895 5695
rect 10333 5729 10367 5763
rect 14657 5729 14691 5763
rect 10149 5593 10183 5627
rect 5457 5525 5491 5559
rect 6009 5525 6043 5559
rect 8217 5525 8251 5559
rect 8309 5525 8343 5559
rect 9321 5525 9355 5559
rect 9505 5525 9539 5559
rect 10517 5525 10551 5559
rect 2605 5321 2639 5355
rect 3433 5321 3467 5355
rect 4261 5321 4295 5355
rect 6929 5321 6963 5355
rect 8217 5321 8251 5355
rect 9781 5321 9815 5355
rect 9965 5321 9999 5355
rect 15301 5321 15335 5355
rect 12173 5253 12207 5287
rect 13829 5253 13863 5287
rect 3249 5185 3283 5219
rect 4077 5185 4111 5219
rect 4813 5185 4847 5219
rect 7481 5185 7515 5219
rect 8401 5185 8435 5219
rect 10609 5185 10643 5219
rect 3801 5117 3835 5151
rect 5181 5117 5215 5151
rect 5448 5117 5482 5151
rect 7297 5117 7331 5151
rect 8033 5117 8067 5151
rect 10793 5117 10827 5151
rect 12449 5117 12483 5151
rect 13921 5117 13955 5151
rect 4629 5049 4663 5083
rect 7389 5049 7423 5083
rect 8668 5049 8702 5083
rect 10333 5049 10367 5083
rect 11060 5049 11094 5083
rect 12694 5049 12728 5083
rect 14188 5049 14222 5083
rect 2973 4981 3007 5015
rect 3065 4981 3099 5015
rect 3893 4981 3927 5015
rect 4721 4981 4755 5015
rect 6561 4981 6595 5015
rect 7757 4981 7791 5015
rect 10425 4981 10459 5015
rect 6009 4777 6043 4811
rect 6377 4777 6411 4811
rect 6837 4777 6871 4811
rect 7021 4777 7055 4811
rect 7389 4777 7423 4811
rect 8309 4777 8343 4811
rect 8677 4777 8711 4811
rect 10149 4777 10183 4811
rect 10977 4777 11011 4811
rect 13553 4777 13587 4811
rect 14381 4777 14415 4811
rect 2329 4709 2363 4743
rect 3617 4709 3651 4743
rect 5273 4709 5307 4743
rect 5825 4709 5859 4743
rect 7481 4709 7515 4743
rect 8217 4709 8251 4743
rect 9045 4709 9079 4743
rect 10517 4709 10551 4743
rect 12164 4709 12198 4743
rect 14749 4709 14783 4743
rect 1501 4641 1535 4675
rect 2053 4641 2087 4675
rect 3065 4641 3099 4675
rect 3157 4641 3191 4675
rect 4721 4641 4755 4675
rect 6469 4641 6503 4675
rect 11345 4641 11379 4675
rect 11897 4641 11931 4675
rect 13921 4641 13955 4675
rect 14841 4641 14875 4675
rect 1685 4573 1719 4607
rect 3249 4573 3283 4607
rect 4261 4573 4295 4607
rect 6561 4573 6595 4607
rect 7573 4573 7607 4607
rect 8401 4573 8435 4607
rect 9137 4573 9171 4607
rect 9321 4573 9355 4607
rect 10609 4573 10643 4607
rect 10793 4573 10827 4607
rect 11437 4573 11471 4607
rect 11621 4573 11655 4607
rect 14013 4573 14047 4607
rect 14105 4573 14139 4607
rect 14933 4573 14967 4607
rect 15301 4573 15335 4607
rect 2697 4505 2731 4539
rect 3801 4505 3835 4539
rect 4537 4505 4571 4539
rect 5549 4505 5583 4539
rect 9965 4505 9999 4539
rect 13277 4505 13311 4539
rect 4905 4437 4939 4471
rect 5181 4437 5215 4471
rect 7849 4437 7883 4471
rect 9781 4437 9815 4471
rect 2881 4233 2915 4267
rect 4353 4233 4387 4267
rect 4905 4233 4939 4267
rect 5825 4233 5859 4267
rect 7297 4233 7331 4267
rect 11529 4233 11563 4267
rect 13277 4233 13311 4267
rect 14013 4233 14047 4267
rect 4813 4165 4847 4199
rect 7573 4165 7607 4199
rect 11345 4165 11379 4199
rect 1501 4097 1535 4131
rect 5549 4097 5583 4131
rect 6009 4097 6043 4131
rect 7113 4097 7147 4131
rect 8125 4097 8159 4131
rect 8217 4097 8251 4131
rect 10057 4097 10091 4131
rect 10977 4097 11011 4131
rect 11253 4097 11287 4131
rect 12081 4097 12115 4131
rect 13001 4097 13035 4131
rect 14565 4097 14599 4131
rect 15393 4097 15427 4131
rect 2973 4029 3007 4063
rect 3240 4029 3274 4063
rect 6193 4029 6227 4063
rect 8033 4029 8067 4063
rect 8493 4029 8527 4063
rect 8861 4029 8895 4063
rect 9965 4029 9999 4063
rect 13829 4029 13863 4063
rect 14473 4029 14507 4063
rect 15209 4029 15243 4063
rect 1768 3961 1802 3995
rect 7021 3961 7055 3995
rect 10701 3961 10735 3995
rect 13461 3961 13495 3995
rect 4445 3893 4479 3927
rect 5273 3893 5307 3927
rect 5365 3893 5399 3927
rect 6285 3893 6319 3927
rect 6469 3893 6503 3927
rect 7665 3893 7699 3927
rect 8677 3893 8711 3927
rect 9045 3893 9079 3927
rect 9321 3893 9355 3927
rect 9505 3893 9539 3927
rect 9873 3893 9907 3927
rect 10333 3893 10367 3927
rect 10793 3893 10827 3927
rect 11897 3893 11931 3927
rect 11989 3893 12023 3927
rect 12449 3893 12483 3927
rect 12817 3893 12851 3927
rect 12909 3893 12943 3927
rect 14381 3893 14415 3927
rect 14841 3893 14875 3927
rect 15301 3893 15335 3927
rect 2053 3689 2087 3723
rect 3157 3689 3191 3723
rect 5549 3689 5583 3723
rect 7665 3689 7699 3723
rect 9413 3689 9447 3723
rect 10057 3689 10091 3723
rect 10517 3689 10551 3723
rect 11345 3689 11379 3723
rect 11713 3689 11747 3723
rect 12541 3689 12575 3723
rect 14841 3689 14875 3723
rect 15577 3689 15611 3723
rect 3525 3621 3559 3655
rect 6276 3621 6310 3655
rect 11253 3621 11287 3655
rect 12081 3621 12115 3655
rect 13001 3621 13035 3655
rect 1593 3553 1627 3587
rect 2789 3553 2823 3587
rect 3617 3553 3651 3587
rect 4436 3553 4470 3587
rect 5641 3553 5675 3587
rect 7481 3553 7515 3587
rect 8033 3553 8067 3587
rect 8300 3553 8334 3587
rect 10425 3553 10459 3587
rect 12909 3553 12943 3587
rect 13553 3553 13587 3587
rect 3709 3485 3743 3519
rect 4169 3485 4203 3519
rect 6009 3485 6043 3519
rect 9689 3485 9723 3519
rect 9965 3485 9999 3519
rect 10701 3485 10735 3519
rect 11437 3485 11471 3519
rect 12173 3485 12207 3519
rect 12357 3485 12391 3519
rect 13185 3485 13219 3519
rect 3065 3417 3099 3451
rect 5825 3417 5859 3451
rect 1777 3349 1811 3383
rect 2421 3349 2455 3383
rect 7389 3349 7423 3383
rect 7941 3349 7975 3383
rect 10885 3349 10919 3383
rect 13369 3349 13403 3383
rect 13829 3349 13863 3383
rect 3341 3145 3375 3179
rect 4077 3145 4111 3179
rect 5089 3145 5123 3179
rect 8309 3145 8343 3179
rect 9873 3145 9907 3179
rect 11529 3145 11563 3179
rect 14381 3145 14415 3179
rect 14841 3145 14875 3179
rect 2605 3077 2639 3111
rect 2973 3077 3007 3111
rect 3985 3077 4019 3111
rect 4997 3077 5031 3111
rect 12909 3077 12943 3111
rect 1685 3009 1719 3043
rect 4721 3009 4755 3043
rect 5641 3009 5675 3043
rect 6377 3009 6411 3043
rect 6561 3009 6595 3043
rect 8493 3009 8527 3043
rect 9965 3009 9999 3043
rect 11989 3009 12023 3043
rect 12173 3009 12207 3043
rect 12725 3009 12759 3043
rect 1501 2941 1535 2975
rect 2053 2941 2087 2975
rect 2421 2941 2455 2975
rect 2789 2941 2823 2975
rect 3157 2941 3191 2975
rect 3525 2941 3559 2975
rect 5457 2941 5491 2975
rect 6837 2941 6871 2975
rect 7104 2941 7138 2975
rect 8760 2941 8794 2975
rect 10232 2941 10266 2975
rect 11897 2941 11931 2975
rect 12449 2941 12483 2975
rect 4445 2873 4479 2907
rect 5549 2873 5583 2907
rect 13001 2941 13035 2975
rect 15025 2941 15059 2975
rect 13246 2873 13280 2907
rect 15301 2873 15335 2907
rect 2237 2805 2271 2839
rect 3709 2805 3743 2839
rect 4537 2805 4571 2839
rect 5917 2805 5951 2839
rect 6285 2805 6319 2839
rect 8217 2805 8251 2839
rect 11345 2805 11379 2839
rect 12909 2805 12943 2839
rect 1501 2601 1535 2635
rect 4169 2601 4203 2635
rect 5641 2601 5675 2635
rect 6009 2601 6043 2635
rect 6653 2601 6687 2635
rect 8217 2601 8251 2635
rect 8585 2601 8619 2635
rect 8861 2601 8895 2635
rect 9229 2601 9263 2635
rect 10241 2601 10275 2635
rect 11069 2601 11103 2635
rect 12081 2601 12115 2635
rect 12633 2601 12667 2635
rect 13001 2601 13035 2635
rect 14381 2601 14415 2635
rect 3893 2533 3927 2567
rect 4629 2533 4663 2567
rect 6101 2533 6135 2567
rect 9321 2533 9355 2567
rect 11437 2533 11471 2567
rect 13737 2533 13771 2567
rect 13921 2533 13955 2567
rect 1593 2465 1627 2499
rect 2493 2465 2527 2499
rect 4537 2465 4571 2499
rect 4997 2465 5031 2499
rect 6469 2465 6503 2499
rect 6929 2465 6963 2499
rect 7297 2465 7331 2499
rect 7665 2465 7699 2499
rect 8033 2465 8067 2499
rect 8401 2465 8435 2499
rect 9781 2465 9815 2499
rect 10609 2465 10643 2499
rect 10701 2465 10735 2499
rect 11529 2465 11563 2499
rect 11897 2465 11931 2499
rect 2237 2397 2271 2431
rect 4721 2397 4755 2431
rect 5365 2397 5399 2431
rect 6285 2397 6319 2431
rect 9505 2397 9539 2431
rect 10793 2397 10827 2431
rect 11621 2397 11655 2431
rect 12357 2397 12391 2431
rect 13093 2397 13127 2431
rect 13277 2397 13311 2431
rect 1777 2329 1811 2363
rect 5181 2329 5215 2363
rect 7481 2329 7515 2363
rect 9965 2329 9999 2363
rect 13461 2329 13495 2363
rect 2053 2261 2087 2295
rect 3617 2261 3651 2295
rect 7113 2261 7147 2295
rect 7849 2261 7883 2295
rect 14105 2261 14139 2295
rect 14197 2261 14231 2295
<< metal1 >>
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 12894 18136 12900 18148
rect 9732 18108 12900 18136
rect 9732 18096 9738 18108
rect 12894 18096 12900 18108
rect 12952 18136 12958 18148
rect 14274 18136 14280 18148
rect 12952 18108 14280 18136
rect 12952 18096 12958 18108
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 4062 17960 4068 18012
rect 4120 18000 4126 18012
rect 12894 18000 12900 18012
rect 4120 17972 12900 18000
rect 4120 17960 4126 17972
rect 12894 17960 12900 17972
rect 12952 17960 12958 18012
rect 2222 17620 2228 17672
rect 2280 17660 2286 17672
rect 2958 17660 2964 17672
rect 2280 17632 2964 17660
rect 2280 17620 2286 17632
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 13262 17660 13268 17672
rect 12584 17632 13268 17660
rect 12584 17620 12590 17632
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 12986 17552 12992 17604
rect 13044 17592 13050 17604
rect 13630 17592 13636 17604
rect 13044 17564 13636 17592
rect 13044 17552 13050 17564
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 198 17484 204 17536
rect 256 17524 262 17536
rect 14366 17524 14372 17536
rect 256 17496 14372 17524
rect 256 17484 262 17496
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 1104 17434 16008 17456
rect 1104 17382 3480 17434
rect 3532 17382 3544 17434
rect 3596 17382 3608 17434
rect 3660 17382 3672 17434
rect 3724 17382 8478 17434
rect 8530 17382 8542 17434
rect 8594 17382 8606 17434
rect 8658 17382 8670 17434
rect 8722 17382 13475 17434
rect 13527 17382 13539 17434
rect 13591 17382 13603 17434
rect 13655 17382 13667 17434
rect 13719 17382 16008 17434
rect 1104 17360 16008 17382
rect 1765 17323 1823 17329
rect 1765 17289 1777 17323
rect 1811 17320 1823 17323
rect 2774 17320 2780 17332
rect 1811 17292 2780 17320
rect 1811 17289 1823 17292
rect 1765 17283 1823 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 7285 17323 7343 17329
rect 7285 17320 7297 17323
rect 7156 17292 7297 17320
rect 7156 17280 7162 17292
rect 7285 17289 7297 17292
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 7558 17280 7564 17332
rect 7616 17320 7622 17332
rect 8113 17323 8171 17329
rect 8113 17320 8125 17323
rect 7616 17292 8125 17320
rect 7616 17280 7622 17292
rect 8113 17289 8125 17292
rect 8159 17289 8171 17323
rect 8113 17283 8171 17289
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 8389 17323 8447 17329
rect 8389 17320 8401 17323
rect 8260 17292 8401 17320
rect 8260 17280 8266 17292
rect 8389 17289 8401 17292
rect 8435 17320 8447 17323
rect 12802 17320 12808 17332
rect 8435 17292 12808 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 14366 17320 14372 17332
rect 14327 17292 14372 17320
rect 14366 17280 14372 17292
rect 14424 17320 14430 17332
rect 14424 17292 14596 17320
rect 14424 17280 14430 17292
rect 1486 17212 1492 17264
rect 1544 17252 1550 17264
rect 12618 17252 12624 17264
rect 1544 17224 12624 17252
rect 1544 17212 1550 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 14568 17261 14596 17292
rect 14553 17255 14611 17261
rect 14553 17221 14565 17255
rect 14599 17221 14611 17255
rect 14553 17215 14611 17221
rect 2498 17144 2504 17196
rect 2556 17184 2562 17196
rect 9493 17187 9551 17193
rect 9493 17184 9505 17187
rect 2556 17156 9505 17184
rect 2556 17144 2562 17156
rect 9493 17153 9505 17156
rect 9539 17184 9551 17187
rect 10134 17184 10140 17196
rect 9539 17156 10140 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 10594 17184 10600 17196
rect 10555 17156 10600 17184
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 11238 17144 11244 17196
rect 11296 17144 11302 17196
rect 11422 17184 11428 17196
rect 11383 17156 11428 17184
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17116 1639 17119
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1627 17088 2053 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 2041 17085 2053 17088
rect 2087 17116 2099 17119
rect 4062 17116 4068 17128
rect 2087 17088 4068 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 7929 17119 7987 17125
rect 7147 17088 7604 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 3234 17008 3240 17060
rect 3292 17048 3298 17060
rect 3605 17051 3663 17057
rect 3605 17048 3617 17051
rect 3292 17020 3617 17048
rect 3292 17008 3298 17020
rect 3605 17017 3617 17020
rect 3651 17048 3663 17051
rect 6546 17048 6552 17060
rect 3651 17020 6552 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 6546 17008 6552 17020
rect 6604 17008 6610 17060
rect 6638 17008 6644 17060
rect 6696 17048 6702 17060
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 6696 17020 7481 17048
rect 6696 17008 6702 17020
rect 7469 17017 7481 17020
rect 7515 17017 7527 17051
rect 7469 17011 7527 17017
rect 7576 16992 7604 17088
rect 7929 17085 7941 17119
rect 7975 17116 7987 17119
rect 8202 17116 8208 17128
rect 7975 17088 8208 17116
rect 7975 17085 7987 17088
rect 7929 17079 7987 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 11256 17116 11284 17144
rect 8312 17088 11284 17116
rect 12621 17119 12679 17125
rect 7834 17008 7840 17060
rect 7892 17048 7898 17060
rect 8312 17048 8340 17088
rect 12621 17085 12633 17119
rect 12667 17085 12679 17119
rect 14918 17116 14924 17128
rect 14879 17088 14924 17116
rect 12621 17079 12679 17085
rect 7892 17020 8340 17048
rect 10413 17051 10471 17057
rect 7892 17008 7898 17020
rect 10413 17017 10425 17051
rect 10459 17048 10471 17051
rect 11241 17051 11299 17057
rect 10459 17020 10916 17048
rect 10459 17017 10471 17020
rect 10413 17011 10471 17017
rect 2774 16940 2780 16992
rect 2832 16980 2838 16992
rect 3145 16983 3203 16989
rect 3145 16980 3157 16983
rect 2832 16952 3157 16980
rect 2832 16940 2838 16952
rect 3145 16949 3157 16952
rect 3191 16980 3203 16983
rect 4982 16980 4988 16992
rect 3191 16952 4988 16980
rect 3191 16949 3203 16952
rect 3145 16943 3203 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 5997 16983 6055 16989
rect 5997 16980 6009 16983
rect 5776 16952 6009 16980
rect 5776 16940 5782 16952
rect 5997 16949 6009 16952
rect 6043 16949 6055 16983
rect 5997 16943 6055 16949
rect 6362 16940 6368 16992
rect 6420 16980 6426 16992
rect 6917 16983 6975 16989
rect 6917 16980 6929 16983
rect 6420 16952 6929 16980
rect 6420 16940 6426 16952
rect 6917 16949 6929 16952
rect 6963 16949 6975 16983
rect 6917 16943 6975 16949
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 7653 16983 7711 16989
rect 7653 16980 7665 16983
rect 7616 16952 7665 16980
rect 7616 16940 7622 16952
rect 7653 16949 7665 16952
rect 7699 16949 7711 16983
rect 7653 16943 7711 16949
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 9217 16983 9275 16989
rect 9217 16980 9229 16983
rect 8904 16952 9229 16980
rect 8904 16940 8910 16952
rect 9217 16949 9229 16952
rect 9263 16949 9275 16983
rect 9858 16980 9864 16992
rect 9819 16952 9864 16980
rect 9217 16943 9275 16949
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 10042 16980 10048 16992
rect 10003 16952 10048 16980
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 10888 16989 10916 17020
rect 11241 17017 11253 17051
rect 11287 17048 11299 17051
rect 12434 17048 12440 17060
rect 11287 17020 12440 17048
rect 11287 17017 11299 17020
rect 11241 17011 11299 17017
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 10873 16983 10931 16989
rect 10560 16952 10605 16980
rect 10560 16940 10566 16952
rect 10873 16949 10885 16983
rect 10919 16949 10931 16983
rect 10873 16943 10931 16949
rect 11330 16940 11336 16992
rect 11388 16980 11394 16992
rect 12636 16980 12664 17079
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 12888 17051 12946 17057
rect 12888 17017 12900 17051
rect 12934 17048 12946 17051
rect 13354 17048 13360 17060
rect 12934 17020 13360 17048
rect 12934 17017 12946 17020
rect 12888 17011 12946 17017
rect 13354 17008 13360 17020
rect 13412 17008 13418 17060
rect 13078 16980 13084 16992
rect 11388 16952 11433 16980
rect 12636 16952 13084 16980
rect 11388 16940 11394 16952
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 13998 16980 14004 16992
rect 13959 16952 14004 16980
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 15013 16983 15071 16989
rect 15013 16980 15025 16983
rect 14792 16952 15025 16980
rect 14792 16940 14798 16952
rect 15013 16949 15025 16952
rect 15059 16949 15071 16983
rect 15013 16943 15071 16949
rect 1104 16890 16008 16912
rect 1104 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 10976 16890
rect 11028 16838 11040 16890
rect 11092 16838 11104 16890
rect 11156 16838 11168 16890
rect 11220 16838 16008 16890
rect 1104 16816 16008 16838
rect 1854 16736 1860 16788
rect 1912 16776 1918 16788
rect 2593 16779 2651 16785
rect 2593 16776 2605 16779
rect 1912 16748 2605 16776
rect 1912 16736 1918 16748
rect 2593 16745 2605 16748
rect 2639 16745 2651 16779
rect 2958 16776 2964 16788
rect 2919 16748 2964 16776
rect 2593 16739 2651 16745
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 3697 16779 3755 16785
rect 3697 16776 3709 16779
rect 3384 16748 3709 16776
rect 3384 16736 3390 16748
rect 3697 16745 3709 16748
rect 3743 16745 3755 16779
rect 3697 16739 3755 16745
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 4709 16779 4767 16785
rect 4709 16776 4721 16779
rect 4304 16748 4721 16776
rect 4304 16736 4310 16748
rect 4709 16745 4721 16748
rect 4755 16745 4767 16779
rect 4709 16739 4767 16745
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 5132 16748 5457 16776
rect 5132 16736 5138 16748
rect 5445 16745 5457 16748
rect 5491 16745 5503 16779
rect 5445 16739 5503 16745
rect 5810 16736 5816 16788
rect 5868 16776 5874 16788
rect 6181 16779 6239 16785
rect 6181 16776 6193 16779
rect 5868 16748 6193 16776
rect 5868 16736 5874 16748
rect 6181 16745 6193 16748
rect 6227 16745 6239 16779
rect 6181 16739 6239 16745
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 6328 16748 6561 16776
rect 6328 16736 6334 16748
rect 6549 16745 6561 16748
rect 6595 16745 6607 16779
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 6549 16739 6607 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 8352 16748 9413 16776
rect 8352 16736 8358 16748
rect 9401 16745 9413 16748
rect 9447 16745 9459 16779
rect 10134 16776 10140 16788
rect 10095 16748 10140 16776
rect 9401 16739 9459 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10318 16736 10324 16788
rect 10376 16776 10382 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 10376 16748 10885 16776
rect 10376 16736 10382 16748
rect 10873 16745 10885 16748
rect 10919 16745 10931 16779
rect 10873 16739 10931 16745
rect 1762 16708 1768 16720
rect 1723 16680 1768 16708
rect 1762 16668 1768 16680
rect 1820 16668 1826 16720
rect 2866 16708 2872 16720
rect 2424 16680 2872 16708
rect 1486 16640 1492 16652
rect 1447 16612 1492 16640
rect 1486 16600 1492 16612
rect 1544 16600 1550 16652
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2314 16640 2320 16652
rect 2087 16612 2320 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 2424 16649 2452 16680
rect 2866 16668 2872 16680
rect 2924 16668 2930 16720
rect 7193 16711 7251 16717
rect 7193 16708 7205 16711
rect 6012 16680 7205 16708
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16609 2467 16643
rect 2774 16640 2780 16652
rect 2735 16612 2780 16640
rect 2409 16603 2467 16609
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 3234 16640 3240 16652
rect 3191 16612 3240 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 3326 16600 3332 16652
rect 3384 16640 3390 16652
rect 3513 16643 3571 16649
rect 3513 16640 3525 16643
rect 3384 16612 3525 16640
rect 3384 16600 3390 16612
rect 3513 16609 3525 16612
rect 3559 16609 3571 16643
rect 3513 16603 3571 16609
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 4798 16640 4804 16652
rect 4571 16612 4804 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 4080 16572 4108 16603
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 4893 16643 4951 16649
rect 4893 16609 4905 16643
rect 4939 16640 4951 16643
rect 5166 16640 5172 16652
rect 4939 16612 5172 16640
rect 4939 16609 4951 16612
rect 4893 16603 4951 16609
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 5534 16640 5540 16652
rect 5307 16612 5540 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 5810 16640 5816 16652
rect 5675 16612 5816 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 6012 16649 6040 16680
rect 7193 16677 7205 16680
rect 7239 16708 7251 16711
rect 8754 16708 8760 16720
rect 7239 16680 8760 16708
rect 7239 16677 7251 16680
rect 7193 16671 7251 16677
rect 8754 16668 8760 16680
rect 8812 16668 8818 16720
rect 9122 16668 9128 16720
rect 9180 16708 9186 16720
rect 9490 16708 9496 16720
rect 9180 16680 9496 16708
rect 9180 16668 9186 16680
rect 9490 16668 9496 16680
rect 9548 16708 9554 16720
rect 10045 16711 10103 16717
rect 10045 16708 10057 16711
rect 9548 16680 10057 16708
rect 9548 16668 9554 16680
rect 10045 16677 10057 16680
rect 10091 16708 10103 16711
rect 10689 16711 10747 16717
rect 10689 16708 10701 16711
rect 10091 16680 10701 16708
rect 10091 16677 10103 16680
rect 10045 16671 10103 16677
rect 10689 16677 10701 16680
rect 10735 16677 10747 16711
rect 10888 16708 10916 16739
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 12437 16779 12495 16785
rect 12437 16776 12449 16779
rect 11480 16748 12449 16776
rect 11480 16736 11486 16748
rect 12437 16745 12449 16748
rect 12483 16745 12495 16779
rect 12437 16739 12495 16745
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 12805 16779 12863 16785
rect 12805 16776 12817 16779
rect 12676 16748 12817 16776
rect 12676 16736 12682 16748
rect 12805 16745 12817 16748
rect 12851 16745 12863 16779
rect 12805 16739 12863 16745
rect 11146 16708 11152 16720
rect 10888 16680 11152 16708
rect 10689 16671 10747 16677
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 11238 16668 11244 16720
rect 11296 16717 11302 16720
rect 11296 16711 11360 16717
rect 11296 16677 11314 16711
rect 11348 16677 11360 16711
rect 13170 16708 13176 16720
rect 13131 16680 13176 16708
rect 11296 16671 11360 16677
rect 11296 16668 11302 16671
rect 13170 16668 13176 16680
rect 13228 16668 13234 16720
rect 13900 16711 13958 16717
rect 13900 16708 13912 16711
rect 13832 16680 13912 16708
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16609 6055 16643
rect 6362 16640 6368 16652
rect 6323 16612 6368 16640
rect 5997 16603 6055 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 6730 16640 6736 16652
rect 6691 16612 6736 16640
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 7644 16643 7702 16649
rect 7644 16609 7656 16643
rect 7690 16640 7702 16643
rect 8202 16640 8208 16652
rect 7690 16612 8208 16640
rect 7690 16609 7702 16612
rect 7644 16603 7702 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8846 16640 8852 16652
rect 8807 16612 8852 16640
rect 8846 16600 8852 16612
rect 8904 16600 8910 16652
rect 9217 16643 9275 16649
rect 9217 16609 9229 16643
rect 9263 16640 9275 16643
rect 9858 16640 9864 16652
rect 9263 16612 9864 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 10152 16612 11069 16640
rect 4080 16544 4568 16572
rect 4540 16516 4568 16544
rect 5442 16532 5448 16584
rect 5500 16532 5506 16584
rect 6822 16532 6828 16584
rect 6880 16572 6886 16584
rect 7377 16575 7435 16581
rect 7377 16572 7389 16575
rect 6880 16544 7389 16572
rect 6880 16532 6886 16544
rect 7377 16541 7389 16544
rect 7423 16541 7435 16575
rect 7377 16535 7435 16541
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 10152 16572 10180 16612
rect 11057 16609 11069 16612
rect 11103 16640 11115 16643
rect 13262 16640 13268 16652
rect 11103 16612 12112 16640
rect 13223 16612 13268 16640
rect 11103 16609 11115 16612
rect 11057 16603 11115 16609
rect 9456 16544 10180 16572
rect 10229 16575 10287 16581
rect 9456 16532 9462 16544
rect 10229 16541 10241 16575
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 2225 16507 2283 16513
rect 2225 16504 2237 16507
rect 992 16476 2237 16504
rect 992 16464 998 16476
rect 2225 16473 2237 16476
rect 2271 16473 2283 16507
rect 3329 16507 3387 16513
rect 3329 16504 3341 16507
rect 2225 16467 2283 16473
rect 2884 16476 3341 16504
rect 2590 16396 2596 16448
rect 2648 16436 2654 16448
rect 2884 16436 2912 16476
rect 3329 16473 3341 16476
rect 3375 16473 3387 16507
rect 3329 16467 3387 16473
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 4249 16507 4307 16513
rect 4249 16504 4261 16507
rect 3936 16476 4261 16504
rect 3936 16464 3942 16476
rect 4249 16473 4261 16476
rect 4295 16473 4307 16507
rect 4249 16467 4307 16473
rect 4522 16464 4528 16516
rect 4580 16464 4586 16516
rect 4614 16464 4620 16516
rect 4672 16504 4678 16516
rect 5077 16507 5135 16513
rect 5077 16504 5089 16507
rect 4672 16476 5089 16504
rect 4672 16464 4678 16476
rect 5077 16473 5089 16476
rect 5123 16473 5135 16507
rect 5460 16504 5488 16532
rect 5813 16507 5871 16513
rect 5813 16504 5825 16507
rect 5460 16476 5825 16504
rect 5077 16467 5135 16473
rect 5813 16473 5825 16476
rect 5859 16473 5871 16507
rect 5813 16467 5871 16473
rect 8757 16507 8815 16513
rect 8757 16473 8769 16507
rect 8803 16504 8815 16507
rect 8938 16504 8944 16516
rect 8803 16476 8944 16504
rect 8803 16473 8815 16476
rect 8757 16467 8815 16473
rect 8938 16464 8944 16476
rect 8996 16504 9002 16516
rect 10244 16504 10272 16535
rect 8996 16476 10272 16504
rect 12084 16504 12112 16612
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13832 16640 13860 16680
rect 13900 16677 13912 16680
rect 13946 16708 13958 16711
rect 13998 16708 14004 16720
rect 13946 16680 14004 16708
rect 13946 16677 13958 16680
rect 13900 16671 13958 16677
rect 13998 16668 14004 16680
rect 14056 16668 14062 16720
rect 13556 16612 13860 16640
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13556 16572 13584 16612
rect 13495 16544 13584 16572
rect 13633 16575 13691 16581
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 13633 16541 13645 16575
rect 13679 16541 13691 16575
rect 13633 16535 13691 16541
rect 13078 16504 13084 16516
rect 12084 16476 13084 16504
rect 8996 16464 9002 16476
rect 13078 16464 13084 16476
rect 13136 16504 13142 16516
rect 13648 16504 13676 16535
rect 13136 16476 13676 16504
rect 13136 16464 13142 16476
rect 2648 16408 2912 16436
rect 2648 16396 2654 16408
rect 8018 16396 8024 16448
rect 8076 16436 8082 16448
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 8076 16408 9045 16436
rect 8076 16396 8082 16408
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 9033 16399 9091 16405
rect 9677 16439 9735 16445
rect 9677 16405 9689 16439
rect 9723 16436 9735 16439
rect 10134 16436 10140 16448
rect 9723 16408 10140 16436
rect 9723 16405 9735 16408
rect 9677 16399 9735 16405
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 10376 16408 10517 16436
rect 10376 16396 10382 16408
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 10505 16399 10563 16405
rect 14918 16396 14924 16448
rect 14976 16436 14982 16448
rect 15013 16439 15071 16445
rect 15013 16436 15025 16439
rect 14976 16408 15025 16436
rect 14976 16396 14982 16408
rect 15013 16405 15025 16408
rect 15059 16405 15071 16439
rect 15013 16399 15071 16405
rect 1104 16346 16008 16368
rect 1104 16294 3480 16346
rect 3532 16294 3544 16346
rect 3596 16294 3608 16346
rect 3660 16294 3672 16346
rect 3724 16294 8478 16346
rect 8530 16294 8542 16346
rect 8594 16294 8606 16346
rect 8658 16294 8670 16346
rect 8722 16294 13475 16346
rect 13527 16294 13539 16346
rect 13591 16294 13603 16346
rect 13655 16294 13667 16346
rect 13719 16294 16008 16346
rect 1104 16272 16008 16294
rect 3050 16192 3056 16244
rect 3108 16232 3114 16244
rect 3421 16235 3479 16241
rect 3421 16232 3433 16235
rect 3108 16204 3433 16232
rect 3108 16192 3114 16204
rect 3421 16201 3433 16204
rect 3467 16201 3479 16235
rect 8202 16232 8208 16244
rect 3421 16195 3479 16201
rect 6840 16204 8208 16232
rect 5534 16124 5540 16176
rect 5592 16164 5598 16176
rect 5721 16167 5779 16173
rect 5721 16164 5733 16167
rect 5592 16136 5733 16164
rect 5592 16124 5598 16136
rect 5721 16133 5733 16136
rect 5767 16164 5779 16167
rect 6638 16164 6644 16176
rect 5767 16136 6644 16164
rect 5767 16133 5779 16136
rect 5721 16127 5779 16133
rect 6638 16124 6644 16136
rect 6696 16124 6702 16176
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16096 6607 16099
rect 6840 16096 6868 16204
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 10042 16232 10048 16244
rect 8312 16204 10048 16232
rect 6595 16068 6868 16096
rect 6595 16065 6607 16068
rect 6549 16059 6607 16065
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 15997 1547 16031
rect 1489 15991 1547 15997
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 3605 16031 3663 16037
rect 3605 16028 3617 16031
rect 3283 16000 3617 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 3605 15997 3617 16000
rect 3651 16028 3663 16031
rect 3878 16028 3884 16040
rect 3651 16000 3884 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 1504 15960 1532 15991
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 6822 16028 6828 16040
rect 6783 16000 6828 16028
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 8312 16028 8340 16204
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16201 10195 16235
rect 10137 16195 10195 16201
rect 10152 16164 10180 16195
rect 10410 16192 10416 16244
rect 10468 16232 10474 16244
rect 11606 16232 11612 16244
rect 10468 16204 11612 16232
rect 10468 16192 10474 16204
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 11882 16192 11888 16244
rect 11940 16232 11946 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 11940 16204 12173 16232
rect 11940 16192 11946 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12492 16204 12537 16232
rect 12492 16192 12498 16204
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13228 16204 13737 16232
rect 13228 16192 13234 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 10152 16136 10824 16164
rect 8662 16096 8668 16108
rect 8623 16068 8668 16096
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10796 16105 10824 16136
rect 12894 16124 12900 16176
rect 12952 16164 12958 16176
rect 13541 16167 13599 16173
rect 13541 16164 13553 16167
rect 12952 16136 13553 16164
rect 12952 16124 12958 16136
rect 13541 16133 13553 16136
rect 13587 16164 13599 16167
rect 13587 16136 14688 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 10689 16099 10747 16105
rect 10689 16096 10701 16099
rect 10192 16068 10701 16096
rect 10192 16056 10198 16068
rect 10689 16065 10701 16068
rect 10735 16065 10747 16099
rect 10689 16059 10747 16065
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16096 10839 16099
rect 11238 16096 11244 16108
rect 10827 16068 11244 16096
rect 10827 16065 10839 16068
rect 10781 16059 10839 16065
rect 11238 16056 11244 16068
rect 11296 16096 11302 16108
rect 11514 16096 11520 16108
rect 11296 16068 11520 16096
rect 11296 16056 11302 16068
rect 11514 16056 11520 16068
rect 11572 16096 11578 16108
rect 11609 16099 11667 16105
rect 11609 16096 11621 16099
rect 11572 16068 11621 16096
rect 11572 16056 11578 16068
rect 11609 16065 11621 16068
rect 11655 16096 11667 16099
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 11655 16068 13001 16096
rect 11655 16065 11667 16068
rect 11609 16059 11667 16065
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13722 16096 13728 16108
rect 13412 16068 13728 16096
rect 13412 16056 13418 16068
rect 13722 16056 13728 16068
rect 13780 16096 13786 16108
rect 14660 16105 14688 16136
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13780 16068 14289 16096
rect 13780 16056 13786 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 15654 16096 15660 16108
rect 15615 16068 15660 16096
rect 14645 16059 14703 16065
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 8757 16031 8815 16037
rect 8757 16028 8769 16031
rect 6932 16000 8340 16028
rect 8404 16000 8769 16028
rect 6932 15960 6960 16000
rect 7098 15969 7104 15972
rect 7092 15960 7104 15969
rect 1504 15932 6960 15960
rect 7059 15932 7104 15960
rect 7092 15923 7104 15932
rect 7098 15920 7104 15923
rect 7156 15920 7162 15972
rect 8110 15920 8116 15972
rect 8168 15960 8174 15972
rect 8404 15960 8432 16000
rect 8757 15997 8769 16000
rect 8803 15997 8815 16031
rect 12158 16028 12164 16040
rect 8757 15991 8815 15997
rect 8864 16000 12164 16028
rect 8168 15932 8432 15960
rect 8168 15920 8174 15932
rect 2498 15892 2504 15904
rect 2459 15864 2504 15892
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 2866 15892 2872 15904
rect 2779 15864 2872 15892
rect 2866 15852 2872 15864
rect 2924 15892 2930 15904
rect 3142 15892 3148 15904
rect 2924 15864 3148 15892
rect 2924 15852 2930 15864
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 3881 15895 3939 15901
rect 3881 15892 3893 15895
rect 3292 15864 3893 15892
rect 3292 15852 3298 15864
rect 3881 15861 3893 15864
rect 3927 15861 3939 15895
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 3881 15855 3939 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 4798 15852 4804 15904
rect 4856 15892 4862 15904
rect 4893 15895 4951 15901
rect 4893 15892 4905 15895
rect 4856 15864 4905 15892
rect 4856 15852 4862 15864
rect 4893 15861 4905 15864
rect 4939 15861 4951 15895
rect 4893 15855 4951 15861
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5353 15895 5411 15901
rect 5353 15892 5365 15895
rect 5224 15864 5365 15892
rect 5224 15852 5230 15864
rect 5353 15861 5365 15864
rect 5399 15892 5411 15895
rect 5442 15892 5448 15904
rect 5399 15864 5448 15892
rect 5399 15861 5411 15864
rect 5353 15855 5411 15861
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 5905 15895 5963 15901
rect 5905 15892 5917 15895
rect 5776 15864 5917 15892
rect 5776 15852 5782 15864
rect 5905 15861 5917 15864
rect 5951 15861 5963 15895
rect 6270 15892 6276 15904
rect 6231 15864 6276 15892
rect 5905 15855 5963 15861
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 6365 15895 6423 15901
rect 6365 15861 6377 15895
rect 6411 15892 6423 15895
rect 7190 15892 7196 15904
rect 6411 15864 7196 15892
rect 6411 15861 6423 15864
rect 6365 15855 6423 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 8404 15892 8432 15932
rect 8481 15963 8539 15969
rect 8481 15929 8493 15963
rect 8527 15960 8539 15963
rect 8864 15960 8892 16000
rect 9140 15972 9168 16000
rect 12158 15988 12164 16000
rect 12216 15988 12222 16040
rect 8527 15932 8892 15960
rect 8527 15929 8539 15932
rect 8481 15923 8539 15929
rect 8938 15920 8944 15972
rect 8996 15969 9002 15972
rect 8996 15963 9060 15969
rect 8996 15929 9014 15963
rect 9048 15929 9060 15963
rect 8996 15923 9060 15929
rect 8996 15920 9002 15923
rect 9122 15920 9128 15972
rect 9180 15920 9186 15972
rect 9214 15920 9220 15972
rect 9272 15960 9278 15972
rect 9674 15960 9680 15972
rect 9272 15932 9680 15960
rect 9272 15920 9278 15932
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 10960 15932 11100 15960
rect 9398 15892 9404 15904
rect 8404 15864 9404 15892
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 10226 15852 10232 15904
rect 10284 15892 10290 15904
rect 10284 15864 10329 15892
rect 10284 15852 10290 15864
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10597 15895 10655 15901
rect 10597 15892 10609 15895
rect 10468 15864 10609 15892
rect 10468 15852 10474 15864
rect 10597 15861 10609 15864
rect 10643 15861 10655 15895
rect 10597 15855 10655 15861
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 10960 15892 10988 15932
rect 11072 15901 11100 15932
rect 11146 15920 11152 15972
rect 11204 15960 11210 15972
rect 11425 15963 11483 15969
rect 11204 15932 11284 15960
rect 11204 15920 11210 15932
rect 10744 15864 10988 15892
rect 11057 15895 11115 15901
rect 10744 15852 10750 15864
rect 11057 15861 11069 15895
rect 11103 15861 11115 15895
rect 11256 15892 11284 15932
rect 11425 15929 11437 15963
rect 11471 15960 11483 15963
rect 11790 15960 11796 15972
rect 11471 15932 11796 15960
rect 11471 15929 11483 15932
rect 11425 15923 11483 15929
rect 11790 15920 11796 15932
rect 11848 15920 11854 15972
rect 11885 15963 11943 15969
rect 11885 15929 11897 15963
rect 11931 15960 11943 15963
rect 12805 15963 12863 15969
rect 12805 15960 12817 15963
rect 11931 15932 12817 15960
rect 11931 15929 11943 15932
rect 11885 15923 11943 15929
rect 12805 15929 12817 15932
rect 12851 15929 12863 15963
rect 12805 15923 12863 15929
rect 12897 15963 12955 15969
rect 12897 15929 12909 15963
rect 12943 15960 12955 15963
rect 13357 15963 13415 15969
rect 13357 15960 13369 15963
rect 12943 15932 13369 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 13357 15929 13369 15932
rect 13403 15960 13415 15963
rect 13403 15932 14412 15960
rect 13403 15929 13415 15932
rect 13357 15923 13415 15929
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11256 15864 11529 15892
rect 11057 15855 11115 15861
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 12710 15852 12716 15904
rect 12768 15892 12774 15904
rect 12912 15892 12940 15923
rect 14090 15892 14096 15904
rect 12768 15864 12940 15892
rect 14051 15864 14096 15892
rect 12768 15852 12774 15864
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14384 15892 14412 15932
rect 14734 15920 14740 15972
rect 14792 15960 14798 15972
rect 14792 15932 14837 15960
rect 14792 15920 14798 15932
rect 16574 15892 16580 15904
rect 14240 15864 14285 15892
rect 14384 15864 16580 15892
rect 14240 15852 14246 15864
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 1104 15802 16008 15824
rect 1104 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 10976 15802
rect 11028 15750 11040 15802
rect 11092 15750 11104 15802
rect 11156 15750 11168 15802
rect 11220 15750 16008 15802
rect 1104 15728 16008 15750
rect 5718 15688 5724 15700
rect 1504 15660 5724 15688
rect 1504 15561 1532 15660
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 7190 15688 7196 15700
rect 7151 15660 7196 15688
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 8018 15688 8024 15700
rect 7979 15660 8024 15688
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 8312 15660 8493 15688
rect 1762 15620 1768 15632
rect 1723 15592 1768 15620
rect 1762 15580 1768 15592
rect 1820 15580 1826 15632
rect 3513 15623 3571 15629
rect 3513 15589 3525 15623
rect 3559 15620 3571 15623
rect 3970 15620 3976 15632
rect 3559 15592 3976 15620
rect 3559 15589 3571 15592
rect 3513 15583 3571 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 8312 15620 8340 15660
rect 8481 15657 8493 15660
rect 8527 15657 8539 15691
rect 8481 15651 8539 15657
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 8628 15660 10149 15688
rect 8628 15648 8634 15660
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 10502 15688 10508 15700
rect 10463 15660 10508 15688
rect 10137 15651 10195 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10873 15691 10931 15697
rect 10873 15688 10885 15691
rect 10744 15660 10885 15688
rect 10744 15648 10750 15660
rect 10873 15657 10885 15660
rect 10919 15657 10931 15691
rect 11330 15688 11336 15700
rect 11291 15660 11336 15688
rect 10873 15651 10931 15657
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 11793 15691 11851 15697
rect 11793 15657 11805 15691
rect 11839 15688 11851 15691
rect 12437 15691 12495 15697
rect 12437 15688 12449 15691
rect 11839 15660 12449 15688
rect 11839 15657 11851 15660
rect 11793 15651 11851 15657
rect 12437 15657 12449 15660
rect 12483 15688 12495 15691
rect 12526 15688 12532 15700
rect 12483 15660 12532 15688
rect 12483 15657 12495 15660
rect 12437 15651 12495 15657
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 12820 15660 13216 15688
rect 8260 15592 8340 15620
rect 8389 15623 8447 15629
rect 8260 15580 8266 15592
rect 8389 15589 8401 15623
rect 8435 15620 8447 15623
rect 8846 15620 8852 15632
rect 8435 15592 8852 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 8846 15580 8852 15592
rect 8904 15620 8910 15632
rect 9582 15620 9588 15632
rect 8904 15592 9588 15620
rect 8904 15580 8910 15592
rect 9582 15580 9588 15592
rect 9640 15580 9646 15632
rect 9858 15580 9864 15632
rect 9916 15620 9922 15632
rect 9916 15592 10180 15620
rect 9916 15580 9922 15592
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15521 1547 15555
rect 1489 15515 1547 15521
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15552 3663 15555
rect 4154 15552 4160 15564
rect 3651 15524 4160 15552
rect 3651 15521 3663 15524
rect 3605 15515 3663 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 5528 15555 5586 15561
rect 5528 15521 5540 15555
rect 5574 15552 5586 15555
rect 7374 15552 7380 15564
rect 5574 15524 7380 15552
rect 5574 15521 5586 15524
rect 5528 15515 5586 15521
rect 7374 15512 7380 15524
rect 7432 15512 7438 15564
rect 7558 15552 7564 15564
rect 7519 15524 7564 15552
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15552 7711 15555
rect 8294 15552 8300 15564
rect 7699 15524 8300 15552
rect 7699 15521 7711 15524
rect 7653 15515 7711 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 8662 15512 8668 15564
rect 8720 15552 8726 15564
rect 8720 15524 8984 15552
rect 8720 15512 8726 15524
rect 3050 15444 3056 15496
rect 3108 15484 3114 15496
rect 3786 15484 3792 15496
rect 3108 15456 3792 15484
rect 3108 15444 3114 15456
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 5258 15484 5264 15496
rect 5219 15456 5264 15484
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8846 15484 8852 15496
rect 8807 15456 8852 15484
rect 8573 15447 8631 15453
rect 6641 15419 6699 15425
rect 6641 15385 6653 15419
rect 6687 15416 6699 15419
rect 7098 15416 7104 15428
rect 6687 15388 7104 15416
rect 6687 15385 6699 15388
rect 6641 15379 6699 15385
rect 7098 15376 7104 15388
rect 7156 15416 7162 15428
rect 7852 15416 7880 15447
rect 8478 15416 8484 15428
rect 7156 15388 8484 15416
rect 7156 15376 7162 15388
rect 8478 15376 8484 15388
rect 8536 15376 8542 15428
rect 2958 15308 2964 15360
rect 3016 15348 3022 15360
rect 3145 15351 3203 15357
rect 3145 15348 3157 15351
rect 3016 15320 3157 15348
rect 3016 15308 3022 15320
rect 3145 15317 3157 15320
rect 3191 15317 3203 15351
rect 3145 15311 3203 15317
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 7650 15348 7656 15360
rect 5500 15320 7656 15348
rect 5500 15308 5506 15320
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 8202 15308 8208 15360
rect 8260 15348 8266 15360
rect 8588 15348 8616 15447
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 8956 15484 8984 15524
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9088 15524 10057 15552
rect 9088 15512 9094 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10152 15552 10180 15592
rect 10226 15580 10232 15632
rect 10284 15620 10290 15632
rect 10965 15623 11023 15629
rect 10965 15620 10977 15623
rect 10284 15592 10977 15620
rect 10284 15580 10290 15592
rect 10965 15589 10977 15592
rect 11011 15589 11023 15623
rect 10965 15583 11023 15589
rect 12158 15580 12164 15632
rect 12216 15620 12222 15632
rect 12820 15620 12848 15660
rect 13078 15620 13084 15632
rect 12216 15592 12848 15620
rect 12912 15592 13084 15620
rect 12216 15580 12222 15592
rect 12912 15561 12940 15592
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 13188 15620 13216 15660
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 14148 15660 14381 15688
rect 14148 15648 14154 15660
rect 14369 15657 14381 15660
rect 14415 15657 14427 15691
rect 14369 15651 14427 15657
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15286 15688 15292 15700
rect 14884 15660 15292 15688
rect 14884 15648 14890 15660
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 16114 15620 16120 15632
rect 13188 15592 16120 15620
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 13170 15561 13176 15564
rect 11701 15555 11759 15561
rect 11701 15552 11713 15555
rect 10152 15524 11713 15552
rect 10045 15515 10103 15521
rect 11701 15521 11713 15524
rect 11747 15552 11759 15555
rect 12897 15555 12955 15561
rect 11747 15524 12296 15552
rect 11747 15521 11759 15524
rect 11701 15515 11759 15521
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 8956 15456 10241 15484
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 11054 15484 11060 15496
rect 11015 15456 11060 15484
rect 10229 15447 10287 15453
rect 11054 15444 11060 15456
rect 11112 15484 11118 15496
rect 11422 15484 11428 15496
rect 11112 15456 11428 15484
rect 11112 15444 11118 15456
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 11514 15444 11520 15496
rect 11572 15484 11578 15496
rect 12268 15493 12296 15524
rect 12897 15521 12909 15555
rect 12943 15521 12955 15555
rect 13164 15552 13176 15561
rect 13131 15524 13176 15552
rect 12897 15515 12955 15521
rect 13164 15515 13176 15524
rect 13170 15512 13176 15515
rect 13228 15512 13234 15564
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 14737 15555 14795 15561
rect 13780 15524 13952 15552
rect 13780 15512 13786 15524
rect 11885 15487 11943 15493
rect 11885 15484 11897 15487
rect 11572 15456 11897 15484
rect 11572 15444 11578 15456
rect 11885 15453 11897 15456
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12618 15484 12624 15496
rect 12299 15456 12624 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 9677 15419 9735 15425
rect 9677 15416 9689 15419
rect 8812 15388 9689 15416
rect 8812 15376 8818 15388
rect 9677 15385 9689 15388
rect 9723 15385 9735 15419
rect 9677 15379 9735 15385
rect 10042 15376 10048 15428
rect 10100 15416 10106 15428
rect 10410 15416 10416 15428
rect 10100 15388 10416 15416
rect 10100 15376 10106 15388
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 10870 15376 10876 15428
rect 10928 15416 10934 15428
rect 10928 15388 11928 15416
rect 10928 15376 10934 15388
rect 8260 15320 8616 15348
rect 8260 15308 8266 15320
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8996 15320 9137 15348
rect 8996 15308 9002 15320
rect 9125 15317 9137 15320
rect 9171 15317 9183 15351
rect 9125 15311 9183 15317
rect 9401 15351 9459 15357
rect 9401 15317 9413 15351
rect 9447 15348 9459 15351
rect 9582 15348 9588 15360
rect 9447 15320 9588 15348
rect 9447 15317 9459 15320
rect 9401 15311 9459 15317
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 10778 15348 10784 15360
rect 10376 15320 10784 15348
rect 10376 15308 10382 15320
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 11900 15348 11928 15388
rect 12158 15376 12164 15428
rect 12216 15416 12222 15428
rect 13924 15416 13952 15524
rect 14737 15521 14749 15555
rect 14783 15552 14795 15555
rect 15010 15552 15016 15564
rect 14783 15524 15016 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 14090 15444 14096 15496
rect 14148 15484 14154 15496
rect 14826 15484 14832 15496
rect 14148 15456 14832 15484
rect 14148 15444 14154 15456
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15453 14979 15487
rect 14921 15447 14979 15453
rect 14277 15419 14335 15425
rect 14277 15416 14289 15419
rect 12216 15388 12940 15416
rect 13924 15388 14289 15416
rect 12216 15376 12222 15388
rect 12710 15348 12716 15360
rect 11900 15320 12716 15348
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 12912 15348 12940 15388
rect 14277 15385 14289 15388
rect 14323 15385 14335 15419
rect 14936 15416 14964 15447
rect 14277 15379 14335 15385
rect 14844 15388 14964 15416
rect 14844 15360 14872 15388
rect 14458 15348 14464 15360
rect 12912 15320 14464 15348
rect 14458 15308 14464 15320
rect 14516 15308 14522 15360
rect 14826 15308 14832 15360
rect 14884 15308 14890 15360
rect 1104 15258 16008 15280
rect 1104 15206 3480 15258
rect 3532 15206 3544 15258
rect 3596 15206 3608 15258
rect 3660 15206 3672 15258
rect 3724 15206 8478 15258
rect 8530 15206 8542 15258
rect 8594 15206 8606 15258
rect 8658 15206 8670 15258
rect 8722 15206 13475 15258
rect 13527 15206 13539 15258
rect 13591 15206 13603 15258
rect 13655 15206 13667 15258
rect 13719 15206 16008 15258
rect 1104 15184 16008 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 2133 15147 2191 15153
rect 2133 15144 2145 15147
rect 1452 15116 2145 15144
rect 1452 15104 1458 15116
rect 2133 15113 2145 15116
rect 2179 15113 2191 15147
rect 4154 15144 4160 15156
rect 4115 15116 4160 15144
rect 2133 15107 2191 15113
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 6822 15144 6828 15156
rect 5276 15116 6828 15144
rect 5276 15088 5304 15116
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 6917 15147 6975 15153
rect 6917 15113 6929 15147
rect 6963 15144 6975 15147
rect 9398 15144 9404 15156
rect 6963 15116 9404 15144
rect 6963 15113 6975 15116
rect 6917 15107 6975 15113
rect 566 15036 572 15088
rect 624 15076 630 15088
rect 1765 15079 1823 15085
rect 1765 15076 1777 15079
rect 624 15048 1777 15076
rect 624 15036 630 15048
rect 1765 15045 1777 15048
rect 1811 15045 1823 15079
rect 1765 15039 1823 15045
rect 3694 15036 3700 15088
rect 3752 15076 3758 15088
rect 4062 15076 4068 15088
rect 3752 15048 4068 15076
rect 3752 15036 3758 15048
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 5258 15076 5264 15088
rect 4448 15048 5264 15076
rect 2317 15011 2375 15017
rect 2317 15008 2329 15011
rect 1596 14980 2329 15008
rect 1596 14949 1624 14980
rect 2317 14977 2329 14980
rect 2363 15008 2375 15011
rect 2363 14980 2820 15008
rect 2363 14977 2375 14980
rect 2317 14971 2375 14977
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14909 2007 14943
rect 2682 14940 2688 14952
rect 2643 14912 2688 14940
rect 1949 14903 2007 14909
rect 1964 14872 1992 14903
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 2792 14940 2820 14980
rect 4246 14940 4252 14952
rect 2792 14912 4252 14940
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 2590 14872 2596 14884
rect 1964 14844 2596 14872
rect 2590 14832 2596 14844
rect 2648 14832 2654 14884
rect 2952 14875 3010 14881
rect 2952 14841 2964 14875
rect 2998 14872 3010 14875
rect 3050 14872 3056 14884
rect 2998 14844 3056 14872
rect 2998 14841 3010 14844
rect 2952 14835 3010 14841
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 4154 14832 4160 14884
rect 4212 14872 4218 14884
rect 4448 14872 4476 15048
rect 5258 15036 5264 15048
rect 5316 15036 5322 15088
rect 6270 15036 6276 15088
rect 6328 15076 6334 15088
rect 6932 15076 6960 15107
rect 9398 15104 9404 15116
rect 9456 15144 9462 15156
rect 9674 15144 9680 15156
rect 9456 15116 9680 15144
rect 9456 15104 9462 15116
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 10410 15144 10416 15156
rect 9824 15116 10416 15144
rect 9824 15104 9830 15116
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 10652 15116 11621 15144
rect 10652 15104 10658 15116
rect 11609 15113 11621 15116
rect 11655 15113 11667 15147
rect 13262 15144 13268 15156
rect 13223 15116 13268 15144
rect 11609 15107 11667 15113
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 14182 15144 14188 15156
rect 14143 15116 14188 15144
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 6328 15048 6960 15076
rect 7561 15079 7619 15085
rect 6328 15036 6334 15048
rect 7561 15045 7573 15079
rect 7607 15076 7619 15079
rect 9030 15076 9036 15088
rect 7607 15048 9036 15076
rect 7607 15045 7619 15048
rect 7561 15039 7619 15045
rect 9030 15036 9036 15048
rect 9088 15036 9094 15088
rect 14642 15076 14648 15088
rect 13004 15048 14648 15076
rect 4614 14968 4620 15020
rect 4672 15008 4678 15020
rect 4709 15011 4767 15017
rect 4709 15008 4721 15011
rect 4672 14980 4721 15008
rect 4672 14968 4678 14980
rect 4709 14977 4721 14980
rect 4755 14977 4767 15011
rect 5537 15011 5595 15017
rect 5537 15008 5549 15011
rect 4709 14971 4767 14977
rect 4908 14980 5549 15008
rect 4908 14952 4936 14980
rect 5537 14977 5549 14980
rect 5583 15008 5595 15011
rect 6730 15008 6736 15020
rect 5583 14980 6736 15008
rect 5583 14977 5595 14980
rect 5537 14971 5595 14977
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7432 14980 8125 15008
rect 7432 14968 7438 14980
rect 8113 14977 8125 14980
rect 8159 15008 8171 15011
rect 8202 15008 8208 15020
rect 8159 14980 8208 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8202 14968 8208 14980
rect 8260 15008 8266 15020
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8260 14980 8953 15008
rect 8260 14968 8266 14980
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 9766 15008 9772 15020
rect 9727 14980 9772 15008
rect 8941 14971 8999 14977
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 11330 14968 11336 15020
rect 11388 15008 11394 15020
rect 13004 15008 13032 15048
rect 14642 15036 14648 15048
rect 14700 15036 14706 15088
rect 11388 14980 13032 15008
rect 13081 15011 13139 15017
rect 11388 14968 11394 14980
rect 13081 14977 13093 15011
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4890 14940 4896 14952
rect 4571 14912 4896 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5442 14940 5448 14952
rect 5403 14912 5448 14940
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8846 14940 8852 14952
rect 7975 14912 8852 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 9030 14900 9036 14952
rect 9088 14940 9094 14952
rect 9088 14912 9260 14940
rect 9088 14900 9094 14912
rect 4212 14844 4476 14872
rect 4617 14875 4675 14881
rect 4212 14832 4218 14844
rect 4617 14841 4629 14875
rect 4663 14872 4675 14875
rect 5721 14875 5779 14881
rect 5721 14872 5733 14875
rect 4663 14844 5733 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 5721 14841 5733 14844
rect 5767 14872 5779 14875
rect 6730 14872 6736 14884
rect 5767 14844 6736 14872
rect 5767 14841 5779 14844
rect 5721 14835 5779 14841
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 8021 14875 8079 14881
rect 7239 14844 7972 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7944 14816 7972 14844
rect 8021 14841 8033 14875
rect 8067 14872 8079 14875
rect 9122 14872 9128 14884
rect 8067 14844 9128 14872
rect 8067 14841 8079 14844
rect 8021 14835 8079 14841
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 9232 14872 9260 14912
rect 9398 14900 9404 14952
rect 9456 14940 9462 14952
rect 9585 14943 9643 14949
rect 9585 14940 9597 14943
rect 9456 14912 9597 14940
rect 9456 14900 9462 14912
rect 9585 14909 9597 14912
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 10229 14943 10287 14949
rect 10229 14909 10241 14943
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 10496 14943 10554 14949
rect 10496 14909 10508 14943
rect 10542 14940 10554 14943
rect 11054 14940 11060 14952
rect 10542 14912 11060 14940
rect 10542 14909 10554 14912
rect 10496 14903 10554 14909
rect 9677 14875 9735 14881
rect 9677 14872 9689 14875
rect 9232 14844 9689 14872
rect 9677 14841 9689 14844
rect 9723 14841 9735 14875
rect 10244 14872 10272 14903
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 11885 14943 11943 14949
rect 11885 14940 11897 14943
rect 11756 14912 11897 14940
rect 11756 14900 11762 14912
rect 11885 14909 11897 14912
rect 11931 14909 11943 14943
rect 11885 14903 11943 14909
rect 12250 14900 12256 14952
rect 12308 14940 12314 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12308 14912 12909 14940
rect 12308 14900 12314 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 13096 14940 13124 14971
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13817 15011 13875 15017
rect 13817 15008 13829 15011
rect 13412 14980 13829 15008
rect 13412 14968 13418 14980
rect 13817 14977 13829 14980
rect 13863 14977 13875 15011
rect 14826 15008 14832 15020
rect 14787 14980 14832 15008
rect 13817 14971 13875 14977
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 15010 15008 15016 15020
rect 14971 14980 15016 15008
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 13170 14940 13176 14952
rect 13083 14912 13176 14940
rect 12897 14903 12955 14909
rect 13170 14900 13176 14912
rect 13228 14940 13234 14952
rect 14844 14940 14872 14968
rect 13228 14912 14872 14940
rect 13228 14900 13234 14912
rect 12158 14872 12164 14884
rect 9677 14835 9735 14841
rect 9968 14844 10272 14872
rect 12119 14844 12164 14872
rect 3326 14764 3332 14816
rect 3384 14804 3390 14816
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 3384 14776 4077 14804
rect 3384 14764 3390 14776
rect 4065 14773 4077 14776
rect 4111 14804 4123 14807
rect 4430 14804 4436 14816
rect 4111 14776 4436 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 4982 14804 4988 14816
rect 4943 14776 4988 14804
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 7374 14804 7380 14816
rect 7335 14776 7380 14804
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 7926 14764 7932 14816
rect 7984 14764 7990 14816
rect 8294 14764 8300 14816
rect 8352 14804 8358 14816
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 8352 14776 8401 14804
rect 8352 14764 8358 14776
rect 8389 14773 8401 14776
rect 8435 14773 8447 14807
rect 8754 14804 8760 14816
rect 8715 14776 8760 14804
rect 8389 14767 8447 14773
rect 8754 14764 8760 14776
rect 8812 14764 8818 14816
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14804 8907 14807
rect 9217 14807 9275 14813
rect 9217 14804 9229 14807
rect 8895 14776 9229 14804
rect 8895 14773 8907 14776
rect 8849 14767 8907 14773
rect 9217 14773 9229 14776
rect 9263 14773 9275 14807
rect 9217 14767 9275 14773
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9968 14804 9996 14844
rect 10134 14804 10140 14816
rect 9364 14776 9996 14804
rect 10095 14776 10140 14804
rect 9364 14764 9370 14776
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 10244 14804 10272 14844
rect 12158 14832 12164 14844
rect 12216 14832 12222 14884
rect 13633 14875 13691 14881
rect 13633 14872 13645 14875
rect 12452 14844 13645 14872
rect 12452 14813 12480 14844
rect 13633 14841 13645 14844
rect 13679 14841 13691 14875
rect 13633 14835 13691 14841
rect 14458 14832 14464 14884
rect 14516 14872 14522 14884
rect 14553 14875 14611 14881
rect 14553 14872 14565 14875
rect 14516 14844 14565 14872
rect 14516 14832 14522 14844
rect 14553 14841 14565 14844
rect 14599 14872 14611 14875
rect 15289 14875 15347 14881
rect 15289 14872 15301 14875
rect 14599 14844 15301 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 15289 14841 15301 14844
rect 15335 14841 15347 14875
rect 15289 14835 15347 14841
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 10244 14776 11713 14804
rect 11701 14773 11713 14776
rect 11747 14773 11759 14807
rect 11701 14767 11759 14773
rect 12437 14807 12495 14813
rect 12437 14773 12449 14807
rect 12483 14773 12495 14807
rect 12802 14804 12808 14816
rect 12763 14776 12808 14804
rect 12437 14767 12495 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 12894 14764 12900 14816
rect 12952 14804 12958 14816
rect 13725 14807 13783 14813
rect 13725 14804 13737 14807
rect 12952 14776 13737 14804
rect 12952 14764 12958 14776
rect 13725 14773 13737 14776
rect 13771 14773 13783 14807
rect 13725 14767 13783 14773
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 14645 14807 14703 14813
rect 14645 14804 14657 14807
rect 14332 14776 14657 14804
rect 14332 14764 14338 14776
rect 14645 14773 14657 14776
rect 14691 14804 14703 14807
rect 15473 14807 15531 14813
rect 15473 14804 15485 14807
rect 14691 14776 15485 14804
rect 14691 14773 14703 14776
rect 14645 14767 14703 14773
rect 15473 14773 15485 14776
rect 15519 14773 15531 14807
rect 15473 14767 15531 14773
rect 1104 14714 16008 14736
rect 1104 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 10976 14714
rect 11028 14662 11040 14714
rect 11092 14662 11104 14714
rect 11156 14662 11168 14714
rect 11220 14662 16008 14714
rect 1104 14640 16008 14662
rect 3053 14603 3111 14609
rect 3053 14569 3065 14603
rect 3099 14600 3111 14603
rect 3786 14600 3792 14612
rect 3099 14572 3792 14600
rect 3099 14569 3111 14572
rect 3053 14563 3111 14569
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 5258 14600 5264 14612
rect 3936 14572 5264 14600
rect 3936 14560 3942 14572
rect 5258 14560 5264 14572
rect 5316 14600 5322 14612
rect 5718 14600 5724 14612
rect 5316 14572 5724 14600
rect 5316 14560 5322 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 5997 14603 6055 14609
rect 5997 14569 6009 14603
rect 6043 14600 6055 14603
rect 6270 14600 6276 14612
rect 6043 14572 6276 14600
rect 6043 14569 6055 14572
rect 5997 14563 6055 14569
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 6917 14603 6975 14609
rect 6917 14569 6929 14603
rect 6963 14600 6975 14603
rect 7374 14600 7380 14612
rect 6963 14572 7380 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 7558 14600 7564 14612
rect 7515 14572 7564 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7837 14603 7895 14609
rect 7837 14600 7849 14603
rect 7708 14572 7849 14600
rect 7708 14560 7714 14572
rect 7837 14569 7849 14572
rect 7883 14600 7895 14603
rect 9398 14600 9404 14612
rect 7883 14572 9404 14600
rect 7883 14569 7895 14572
rect 7837 14563 7895 14569
rect 9398 14560 9404 14572
rect 9456 14600 9462 14612
rect 12802 14600 12808 14612
rect 9456 14572 12808 14600
rect 9456 14560 9462 14572
rect 12802 14560 12808 14572
rect 12860 14600 12866 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 12860 14572 13553 14600
rect 12860 14560 12866 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 13541 14563 13599 14569
rect 2682 14532 2688 14544
rect 1688 14504 2688 14532
rect 1688 14473 1716 14504
rect 2682 14492 2688 14504
rect 2740 14532 2746 14544
rect 4062 14532 4068 14544
rect 2740 14504 4068 14532
rect 2740 14492 2746 14504
rect 4062 14492 4068 14504
rect 4120 14492 4126 14544
rect 4246 14492 4252 14544
rect 4304 14532 4310 14544
rect 4304 14504 5120 14532
rect 4304 14492 4310 14504
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14433 1731 14467
rect 1673 14427 1731 14433
rect 1940 14467 1998 14473
rect 1940 14433 1952 14467
rect 1986 14464 1998 14467
rect 3510 14464 3516 14476
rect 1986 14436 2728 14464
rect 3471 14436 3516 14464
rect 1986 14433 1998 14436
rect 1940 14427 1998 14433
rect 2700 14260 2728 14436
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 3605 14399 3663 14405
rect 3605 14396 3617 14399
rect 2924 14368 3617 14396
rect 2924 14356 2930 14368
rect 3605 14365 3617 14368
rect 3651 14365 3663 14399
rect 3786 14396 3792 14408
rect 3747 14368 3792 14396
rect 3605 14359 3663 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 4080 14396 4108 14492
rect 4430 14473 4436 14476
rect 4424 14464 4436 14473
rect 4391 14436 4436 14464
rect 4424 14427 4436 14436
rect 4430 14424 4436 14427
rect 4488 14424 4494 14476
rect 5092 14464 5120 14504
rect 5166 14492 5172 14544
rect 5224 14532 5230 14544
rect 8297 14535 8355 14541
rect 8297 14532 8309 14535
rect 5224 14504 8309 14532
rect 5224 14492 5230 14504
rect 8297 14501 8309 14504
rect 8343 14501 8355 14535
rect 10502 14532 10508 14544
rect 8297 14495 8355 14501
rect 8956 14504 9076 14532
rect 8956 14476 8984 14504
rect 6089 14467 6147 14473
rect 6089 14464 6101 14467
rect 5092 14436 6101 14464
rect 6089 14433 6101 14436
rect 6135 14464 6147 14467
rect 6638 14464 6644 14476
rect 6135 14436 6644 14464
rect 6135 14433 6147 14436
rect 6089 14427 6147 14433
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14464 6883 14467
rect 7926 14464 7932 14476
rect 6871 14436 7932 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 8754 14424 8760 14476
rect 8812 14464 8818 14476
rect 8812 14436 8857 14464
rect 8812 14424 8818 14436
rect 8938 14424 8944 14476
rect 8996 14424 9002 14476
rect 4157 14399 4215 14405
rect 4157 14396 4169 14399
rect 4080 14368 4169 14396
rect 4157 14365 4169 14368
rect 4203 14365 4215 14399
rect 6178 14396 6184 14408
rect 4157 14359 4215 14365
rect 5552 14368 6184 14396
rect 2774 14288 2780 14340
rect 2832 14328 2838 14340
rect 5552 14337 5580 14368
rect 6178 14356 6184 14368
rect 6236 14396 6242 14408
rect 7009 14399 7067 14405
rect 6236 14368 6684 14396
rect 6236 14356 6242 14368
rect 3145 14331 3203 14337
rect 3145 14328 3157 14331
rect 2832 14300 3157 14328
rect 2832 14288 2838 14300
rect 3145 14297 3157 14300
rect 3191 14297 3203 14331
rect 3145 14291 3203 14297
rect 5537 14331 5595 14337
rect 5537 14297 5549 14331
rect 5583 14297 5595 14331
rect 6656 14328 6684 14368
rect 7009 14365 7021 14399
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8202 14396 8208 14408
rect 8159 14368 8208 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 7024 14328 7052 14359
rect 8202 14356 8208 14368
rect 8260 14396 8266 14408
rect 8846 14396 8852 14408
rect 8260 14368 8708 14396
rect 8807 14368 8852 14396
rect 8260 14356 8266 14368
rect 6656 14300 7052 14328
rect 8297 14331 8355 14337
rect 5537 14291 5595 14297
rect 8297 14297 8309 14331
rect 8343 14328 8355 14331
rect 8389 14331 8447 14337
rect 8389 14328 8401 14331
rect 8343 14300 8401 14328
rect 8343 14297 8355 14300
rect 8297 14291 8355 14297
rect 8389 14297 8401 14300
rect 8435 14297 8447 14331
rect 8680 14328 8708 14368
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9048 14405 9076 14504
rect 9784 14504 10508 14532
rect 9122 14424 9128 14476
rect 9180 14424 9186 14476
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9364 14436 9689 14464
rect 9364 14424 9370 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9033 14399 9091 14405
rect 9033 14365 9045 14399
rect 9079 14365 9091 14399
rect 9140 14396 9168 14424
rect 9784 14396 9812 14504
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 10594 14492 10600 14544
rect 10652 14532 10658 14544
rect 11394 14535 11452 14541
rect 11394 14532 11406 14535
rect 10652 14504 11406 14532
rect 10652 14492 10658 14504
rect 11394 14501 11406 14504
rect 11440 14501 11452 14535
rect 11394 14495 11452 14501
rect 12158 14492 12164 14544
rect 12216 14532 12222 14544
rect 13081 14535 13139 14541
rect 13081 14532 13093 14535
rect 12216 14504 13093 14532
rect 12216 14492 12222 14504
rect 13081 14501 13093 14504
rect 13127 14501 13139 14535
rect 13081 14495 13139 14501
rect 14185 14535 14243 14541
rect 14185 14501 14197 14535
rect 14231 14532 14243 14535
rect 15010 14532 15016 14544
rect 14231 14504 15016 14532
rect 14231 14501 14243 14504
rect 14185 14495 14243 14501
rect 15010 14492 15016 14504
rect 15068 14492 15074 14544
rect 9944 14467 10002 14473
rect 9944 14433 9956 14467
rect 9990 14464 10002 14467
rect 10410 14464 10416 14476
rect 9990 14436 10416 14464
rect 9990 14433 10002 14436
rect 9944 14427 10002 14433
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 11149 14467 11207 14473
rect 11149 14433 11161 14467
rect 11195 14464 11207 14467
rect 11238 14464 11244 14476
rect 11195 14436 11244 14464
rect 11195 14433 11207 14436
rect 11149 14427 11207 14433
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13725 14467 13783 14473
rect 13725 14464 13737 14467
rect 13228 14436 13737 14464
rect 13228 14424 13234 14436
rect 13725 14433 13737 14436
rect 13771 14433 13783 14467
rect 13725 14427 13783 14433
rect 9140 14368 9812 14396
rect 13265 14399 13323 14405
rect 9033 14359 9091 14365
rect 13265 14365 13277 14399
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14365 14151 14399
rect 14366 14396 14372 14408
rect 14327 14368 14372 14396
rect 14093 14359 14151 14365
rect 9309 14331 9367 14337
rect 8680 14300 9168 14328
rect 8389 14291 8447 14297
rect 4154 14260 4160 14272
rect 2700 14232 4160 14260
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 5684 14232 5729 14260
rect 5684 14220 5690 14232
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6457 14263 6515 14269
rect 6457 14260 6469 14263
rect 5868 14232 6469 14260
rect 5868 14220 5874 14232
rect 6457 14229 6469 14232
rect 6503 14229 6515 14263
rect 6457 14223 6515 14229
rect 6638 14220 6644 14272
rect 6696 14260 6702 14272
rect 7285 14263 7343 14269
rect 7285 14260 7297 14263
rect 6696 14232 7297 14260
rect 6696 14220 6702 14232
rect 7285 14229 7297 14232
rect 7331 14260 7343 14263
rect 9030 14260 9036 14272
rect 7331 14232 9036 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 9140 14260 9168 14300
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 9398 14328 9404 14340
rect 9355 14300 9404 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14328 9551 14331
rect 9674 14328 9680 14340
rect 9539 14300 9680 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 12529 14331 12587 14337
rect 12529 14297 12541 14331
rect 12575 14328 12587 14331
rect 13078 14328 13084 14340
rect 12575 14300 13084 14328
rect 12575 14297 12587 14300
rect 12529 14291 12587 14297
rect 13078 14288 13084 14300
rect 13136 14328 13142 14340
rect 13280 14328 13308 14359
rect 13136 14300 13308 14328
rect 14108 14328 14136 14359
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 14108 14300 15424 14328
rect 13136 14288 13142 14300
rect 15396 14272 15424 14300
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 9140 14232 11069 14260
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 12710 14260 12716 14272
rect 12671 14232 12716 14260
rect 11057 14223 11115 14229
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 15378 14260 15384 14272
rect 15339 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 1104 14170 16008 14192
rect 1104 14118 3480 14170
rect 3532 14118 3544 14170
rect 3596 14118 3608 14170
rect 3660 14118 3672 14170
rect 3724 14118 8478 14170
rect 8530 14118 8542 14170
rect 8594 14118 8606 14170
rect 8658 14118 8670 14170
rect 8722 14118 13475 14170
rect 13527 14118 13539 14170
rect 13591 14118 13603 14170
rect 13655 14118 13667 14170
rect 13719 14118 16008 14170
rect 1104 14096 16008 14118
rect 3142 14056 3148 14068
rect 3103 14028 3148 14056
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 5534 14056 5540 14068
rect 4847 14028 5540 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 9766 14056 9772 14068
rect 6420 14028 9352 14056
rect 9727 14028 9772 14056
rect 6420 14016 6426 14028
rect 5166 13988 5172 14000
rect 1514 13960 5172 13988
rect 1514 13861 1542 13960
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 5626 13988 5632 14000
rect 5276 13960 5632 13988
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 2961 13923 3019 13929
rect 2832 13892 2877 13920
rect 2832 13880 2838 13892
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3326 13920 3332 13932
rect 3007 13892 3332 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 4154 13920 4160 13932
rect 3835 13892 4160 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 4154 13880 4160 13892
rect 4212 13920 4218 13932
rect 4614 13920 4620 13932
rect 4212 13892 4620 13920
rect 4212 13880 4218 13892
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 5276 13929 5304 13960
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 6454 13988 6460 14000
rect 6012 13960 6460 13988
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13920 5503 13923
rect 6012 13920 6040 13960
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 9324 13988 9352 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 11330 14056 11336 14068
rect 9876 14028 11336 14056
rect 9876 13988 9904 14028
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 14366 14056 14372 14068
rect 11572 14028 14372 14056
rect 11572 14016 11578 14028
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 15010 14016 15016 14068
rect 15068 14065 15074 14068
rect 15068 14059 15117 14065
rect 15068 14025 15071 14059
rect 15105 14025 15117 14059
rect 15068 14019 15117 14025
rect 15068 14016 15074 14019
rect 9324 13960 9904 13988
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 13170 13988 13176 14000
rect 10192 13960 13176 13988
rect 10192 13948 10198 13960
rect 13170 13948 13176 13960
rect 13228 13948 13234 14000
rect 14737 13991 14795 13997
rect 14737 13988 14749 13991
rect 14384 13960 14749 13988
rect 6178 13920 6184 13932
rect 5491 13892 6040 13920
rect 6139 13892 6184 13920
rect 5491 13889 5503 13892
rect 5445 13883 5503 13889
rect 6178 13880 6184 13892
rect 6236 13920 6242 13932
rect 6236 13892 6960 13920
rect 6236 13880 6242 13892
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13821 1547 13855
rect 1489 13815 1547 13821
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 4246 13852 4252 13864
rect 3651 13824 4252 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13852 4399 13855
rect 4982 13852 4988 13864
rect 4387 13824 4988 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5718 13812 5724 13864
rect 5776 13852 5782 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5776 13824 6101 13852
rect 5776 13812 5782 13824
rect 6089 13821 6101 13824
rect 6135 13852 6147 13855
rect 6457 13855 6515 13861
rect 6457 13852 6469 13855
rect 6135 13824 6469 13852
rect 6135 13821 6147 13824
rect 6089 13815 6147 13821
rect 6457 13821 6469 13824
rect 6503 13821 6515 13855
rect 6822 13852 6828 13864
rect 6783 13824 6828 13852
rect 6457 13815 6515 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 6932 13852 6960 13892
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 9732 13892 11989 13920
rect 9732 13880 9738 13892
rect 11977 13889 11989 13892
rect 12023 13920 12035 13923
rect 12158 13920 12164 13932
rect 12023 13892 12164 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 13078 13920 13084 13932
rect 13039 13892 13084 13920
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 13136 13892 13492 13920
rect 13136 13880 13142 13892
rect 7081 13855 7139 13861
rect 7081 13852 7093 13855
rect 6932 13824 7093 13852
rect 7081 13821 7093 13824
rect 7127 13821 7139 13855
rect 7081 13815 7139 13821
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 8110 13852 8116 13864
rect 7616 13824 8116 13852
rect 7616 13812 7622 13824
rect 8110 13812 8116 13824
rect 8168 13852 8174 13864
rect 8386 13852 8392 13864
rect 8168 13824 8392 13852
rect 8168 13812 8174 13824
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 8656 13855 8714 13861
rect 8656 13821 8668 13855
rect 8702 13852 8714 13855
rect 8938 13852 8944 13864
rect 8702 13824 8944 13852
rect 8702 13821 8714 13824
rect 8656 13815 8714 13821
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 9030 13812 9036 13864
rect 9088 13852 9094 13864
rect 12253 13855 12311 13861
rect 12253 13852 12265 13855
rect 9088 13824 12265 13852
rect 9088 13812 9094 13824
rect 12253 13821 12265 13824
rect 12299 13852 12311 13855
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12299 13824 13001 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12989 13821 13001 13824
rect 13035 13821 13047 13855
rect 12989 13815 13047 13821
rect 13262 13812 13268 13864
rect 13320 13852 13326 13864
rect 13357 13855 13415 13861
rect 13357 13852 13369 13855
rect 13320 13824 13369 13852
rect 13320 13812 13326 13824
rect 13357 13821 13369 13824
rect 13403 13821 13415 13855
rect 13464 13852 13492 13892
rect 13613 13855 13671 13861
rect 13613 13852 13625 13855
rect 13464 13824 13625 13852
rect 13357 13815 13415 13821
rect 13613 13821 13625 13824
rect 13659 13821 13671 13855
rect 14384 13852 14412 13960
rect 14737 13957 14749 13960
rect 14783 13988 14795 13991
rect 14826 13988 14832 14000
rect 14783 13960 14832 13988
rect 14783 13957 14795 13960
rect 14737 13951 14795 13957
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 13613 13815 13671 13821
rect 13740 13824 14412 13852
rect 13740 13796 13768 13824
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15010 13861 15016 13864
rect 14988 13855 15016 13861
rect 14988 13852 15000 13855
rect 14792 13824 15000 13852
rect 14792 13812 14798 13824
rect 14988 13821 15000 13824
rect 14988 13815 15016 13821
rect 15010 13812 15016 13815
rect 15068 13812 15074 13864
rect 2685 13787 2743 13793
rect 2685 13753 2697 13787
rect 2731 13784 2743 13787
rect 2958 13784 2964 13796
rect 2731 13756 2964 13784
rect 2731 13753 2743 13756
rect 2685 13747 2743 13753
rect 2958 13744 2964 13756
rect 3016 13744 3022 13796
rect 5169 13787 5227 13793
rect 5169 13753 5181 13787
rect 5215 13784 5227 13787
rect 5810 13784 5816 13796
rect 5215 13756 5816 13784
rect 5215 13753 5227 13756
rect 5169 13747 5227 13753
rect 5810 13744 5816 13756
rect 5868 13744 5874 13796
rect 5902 13744 5908 13796
rect 5960 13784 5966 13796
rect 6638 13784 6644 13796
rect 5960 13756 6644 13784
rect 5960 13744 5966 13756
rect 6638 13744 6644 13756
rect 6696 13784 6702 13796
rect 6696 13756 10916 13784
rect 6696 13744 6702 13756
rect 1486 13676 1492 13728
rect 1544 13716 1550 13728
rect 2317 13719 2375 13725
rect 2317 13716 2329 13719
rect 1544 13688 2329 13716
rect 1544 13676 1550 13688
rect 2317 13685 2329 13688
rect 2363 13685 2375 13719
rect 2317 13679 2375 13685
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3513 13719 3571 13725
rect 3513 13716 3525 13719
rect 3292 13688 3525 13716
rect 3292 13676 3298 13688
rect 3513 13685 3525 13688
rect 3559 13716 3571 13719
rect 3602 13716 3608 13728
rect 3559 13688 3608 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 3602 13676 3608 13688
rect 3660 13676 3666 13728
rect 4433 13719 4491 13725
rect 4433 13685 4445 13719
rect 4479 13716 4491 13719
rect 4522 13716 4528 13728
rect 4479 13688 4528 13716
rect 4479 13685 4491 13688
rect 4433 13679 4491 13685
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 5626 13716 5632 13728
rect 5587 13688 5632 13716
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 5718 13676 5724 13728
rect 5776 13716 5782 13728
rect 5997 13719 6055 13725
rect 5997 13716 6009 13719
rect 5776 13688 6009 13716
rect 5776 13676 5782 13688
rect 5997 13685 6009 13688
rect 6043 13716 6055 13719
rect 6822 13716 6828 13728
rect 6043 13688 6828 13716
rect 6043 13685 6055 13688
rect 5997 13679 6055 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 8202 13716 8208 13728
rect 8163 13688 8208 13716
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 10778 13716 10784 13728
rect 9088 13688 10784 13716
rect 9088 13676 9094 13688
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 10888 13716 10916 13756
rect 12158 13744 12164 13796
rect 12216 13784 12222 13796
rect 12897 13787 12955 13793
rect 12897 13784 12909 13787
rect 12216 13756 12909 13784
rect 12216 13744 12222 13756
rect 12897 13753 12909 13756
rect 12943 13753 12955 13787
rect 12897 13747 12955 13753
rect 13722 13744 13728 13796
rect 13780 13744 13786 13796
rect 12342 13716 12348 13728
rect 10888 13688 12348 13716
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12529 13719 12587 13725
rect 12529 13685 12541 13719
rect 12575 13716 12587 13719
rect 13354 13716 13360 13728
rect 12575 13688 13360 13716
rect 12575 13685 12587 13688
rect 12529 13679 12587 13685
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 1104 13626 16008 13648
rect 1104 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 10976 13626
rect 11028 13574 11040 13626
rect 11092 13574 11104 13626
rect 11156 13574 11168 13626
rect 11220 13574 16008 13626
rect 1104 13552 16008 13574
rect 2866 13512 2872 13524
rect 2827 13484 2872 13512
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5629 13515 5687 13521
rect 5629 13512 5641 13515
rect 5592 13484 5641 13512
rect 5592 13472 5598 13484
rect 5629 13481 5641 13484
rect 5675 13481 5687 13515
rect 5629 13475 5687 13481
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 8938 13512 8944 13524
rect 6595 13484 8524 13512
rect 8899 13484 8944 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 3050 13404 3056 13456
rect 3108 13444 3114 13456
rect 3237 13447 3295 13453
rect 3237 13444 3249 13447
rect 3108 13416 3249 13444
rect 3108 13404 3114 13416
rect 3237 13413 3249 13416
rect 3283 13444 3295 13447
rect 3789 13447 3847 13453
rect 3789 13444 3801 13447
rect 3283 13416 3801 13444
rect 3283 13413 3295 13416
rect 3237 13407 3295 13413
rect 3789 13413 3801 13416
rect 3835 13444 3847 13447
rect 3970 13444 3976 13456
rect 3835 13416 3976 13444
rect 3835 13413 3847 13416
rect 3789 13407 3847 13413
rect 3970 13404 3976 13416
rect 4028 13404 4034 13456
rect 4522 13404 4528 13456
rect 4580 13444 4586 13456
rect 4893 13447 4951 13453
rect 4893 13444 4905 13447
rect 4580 13416 4905 13444
rect 4580 13404 4586 13416
rect 4893 13413 4905 13416
rect 4939 13444 4951 13447
rect 6362 13444 6368 13456
rect 4939 13416 6368 13444
rect 4939 13413 4951 13416
rect 4893 13407 4951 13413
rect 6362 13404 6368 13416
rect 6420 13404 6426 13456
rect 6733 13447 6791 13453
rect 6733 13413 6745 13447
rect 6779 13444 6791 13447
rect 6822 13444 6828 13456
rect 6779 13416 6828 13444
rect 6779 13413 6791 13416
rect 6733 13407 6791 13413
rect 6822 13404 6828 13416
rect 6880 13444 6886 13456
rect 7926 13444 7932 13456
rect 6880 13416 7932 13444
rect 6880 13404 6886 13416
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 8496 13444 8524 13484
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 9539 13484 11437 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 11425 13481 11437 13484
rect 11471 13512 11483 13515
rect 11606 13512 11612 13524
rect 11471 13484 11612 13512
rect 11471 13481 11483 13484
rect 11425 13475 11483 13481
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 13265 13515 13323 13521
rect 13265 13512 13277 13515
rect 12768 13484 13277 13512
rect 12768 13472 12774 13484
rect 13265 13481 13277 13484
rect 13311 13481 13323 13515
rect 13265 13475 13323 13481
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13412 13484 13457 13512
rect 13412 13472 13418 13484
rect 9674 13444 9680 13456
rect 8496 13416 9680 13444
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 11330 13444 11336 13456
rect 10060 13416 11336 13444
rect 1486 13376 1492 13388
rect 1447 13348 1492 13376
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 5350 13336 5356 13388
rect 5408 13376 5414 13388
rect 5537 13379 5595 13385
rect 5537 13376 5549 13379
rect 5408 13348 5549 13376
rect 5408 13336 5414 13348
rect 5537 13345 5549 13348
rect 5583 13345 5595 13379
rect 5537 13339 5595 13345
rect 7828 13379 7886 13385
rect 7828 13345 7840 13379
rect 7874 13376 7886 13379
rect 9122 13376 9128 13388
rect 7874 13348 9128 13376
rect 7874 13345 7886 13348
rect 7828 13339 7886 13345
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 10060 13385 10088 13416
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 11701 13447 11759 13453
rect 11701 13444 11713 13447
rect 11572 13416 11713 13444
rect 11572 13404 11578 13416
rect 11701 13413 11713 13416
rect 11747 13444 11759 13447
rect 12437 13447 12495 13453
rect 12437 13444 12449 13447
rect 11747 13416 12449 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 12437 13413 12449 13416
rect 12483 13413 12495 13447
rect 12437 13407 12495 13413
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13413 12587 13447
rect 12529 13407 12587 13413
rect 9861 13379 9919 13385
rect 9861 13345 9873 13379
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 10045 13379 10103 13385
rect 10045 13345 10057 13379
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 10312 13379 10370 13385
rect 10312 13345 10324 13379
rect 10358 13376 10370 13379
rect 10594 13376 10600 13388
rect 10358 13348 10600 13376
rect 10358 13345 10370 13348
rect 10312 13339 10370 13345
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2406 13268 2412 13320
rect 2464 13308 2470 13320
rect 3329 13311 3387 13317
rect 3329 13308 3341 13311
rect 2464 13280 3341 13308
rect 2464 13268 2470 13280
rect 3329 13277 3341 13280
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 4154 13308 4160 13320
rect 3559 13280 4160 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4246 13268 4252 13320
rect 4304 13308 4310 13320
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 4304 13280 4353 13308
rect 4304 13268 4310 13280
rect 4341 13277 4353 13280
rect 4387 13308 4399 13311
rect 4522 13308 4528 13320
rect 4387 13280 4528 13308
rect 4387 13277 4399 13280
rect 4341 13271 4399 13277
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 5810 13308 5816 13320
rect 5771 13280 5816 13308
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 7558 13308 7564 13320
rect 7519 13280 7564 13308
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 9214 13308 9220 13320
rect 9175 13280 9220 13308
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 3602 13200 3608 13252
rect 3660 13240 3666 13252
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 3660 13212 4077 13240
rect 3660 13200 3666 13212
rect 4065 13209 4077 13212
rect 4111 13240 4123 13243
rect 6549 13243 6607 13249
rect 6549 13240 6561 13243
rect 4111 13212 6561 13240
rect 4111 13209 4123 13212
rect 4065 13203 4123 13209
rect 6549 13209 6561 13212
rect 6595 13209 6607 13243
rect 9876 13240 9904 13339
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 12544 13320 12572 13407
rect 11514 13268 11520 13320
rect 11572 13308 11578 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11572 13280 11897 13308
rect 11572 13268 11578 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 13078 13308 13084 13320
rect 12759 13280 13084 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 13722 13308 13728 13320
rect 13587 13280 13728 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 6549 13203 6607 13209
rect 8496 13212 9904 13240
rect 12069 13243 12127 13249
rect 5166 13172 5172 13184
rect 5127 13144 5172 13172
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 7282 13172 7288 13184
rect 7243 13144 7288 13172
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7926 13132 7932 13184
rect 7984 13172 7990 13184
rect 8496 13172 8524 13212
rect 12069 13209 12081 13243
rect 12115 13240 12127 13243
rect 12250 13240 12256 13252
rect 12115 13212 12256 13240
rect 12115 13209 12127 13212
rect 12069 13203 12127 13209
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12894 13240 12900 13252
rect 12855 13212 12900 13240
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 7984 13144 8524 13172
rect 7984 13132 7990 13144
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8996 13144 9045 13172
rect 8996 13132 9002 13144
rect 9033 13141 9045 13144
rect 9079 13141 9091 13175
rect 9033 13135 9091 13141
rect 9122 13132 9128 13184
rect 9180 13172 9186 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9180 13144 9505 13172
rect 9180 13132 9186 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 11698 13172 11704 13184
rect 9723 13144 11704 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 1104 13082 16008 13104
rect 1104 13030 3480 13082
rect 3532 13030 3544 13082
rect 3596 13030 3608 13082
rect 3660 13030 3672 13082
rect 3724 13030 8478 13082
rect 8530 13030 8542 13082
rect 8594 13030 8606 13082
rect 8658 13030 8670 13082
rect 8722 13030 13475 13082
rect 13527 13030 13539 13082
rect 13591 13030 13603 13082
rect 13655 13030 13667 13082
rect 13719 13030 16008 13082
rect 1104 13008 16008 13030
rect 2406 12968 2412 12980
rect 2367 12940 2412 12968
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3878 12968 3884 12980
rect 2832 12940 3884 12968
rect 2832 12928 2838 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 5350 12968 5356 12980
rect 5311 12940 5356 12968
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 6638 12968 6644 12980
rect 6595 12940 6644 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 8573 12971 8631 12977
rect 8573 12937 8585 12971
rect 8619 12968 8631 12971
rect 8846 12968 8852 12980
rect 8619 12940 8852 12968
rect 8619 12937 8631 12940
rect 8573 12931 8631 12937
rect 8846 12928 8852 12940
rect 8904 12928 8910 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10410 12968 10416 12980
rect 10008 12940 10416 12968
rect 10008 12928 10014 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 10560 12940 11069 12968
rect 10560 12928 10566 12940
rect 11057 12937 11069 12940
rect 11103 12937 11115 12971
rect 13541 12971 13599 12977
rect 11057 12931 11115 12937
rect 11164 12940 13492 12968
rect 6178 12900 6184 12912
rect 1504 12872 3280 12900
rect 6139 12872 6184 12900
rect 1504 12773 1532 12872
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1636 12804 1685 12832
rect 1636 12792 1642 12804
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12801 3111 12835
rect 3252 12832 3280 12872
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 7190 12860 7196 12912
rect 7248 12900 7254 12912
rect 7466 12900 7472 12912
rect 7248 12872 7472 12900
rect 7248 12860 7254 12872
rect 7466 12860 7472 12872
rect 7524 12900 7530 12912
rect 11164 12900 11192 12940
rect 7524 12872 11192 12900
rect 11256 12872 12388 12900
rect 7524 12860 7530 12872
rect 3252 12804 3372 12832
rect 3053 12795 3111 12801
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12733 1547 12767
rect 1489 12727 1547 12733
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 2832 12736 2877 12764
rect 2832 12724 2838 12736
rect 3068 12696 3096 12795
rect 3234 12764 3240 12776
rect 3195 12736 3240 12764
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3344 12764 3372 12804
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5684 12804 5825 12832
rect 5684 12792 5690 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12832 6055 12835
rect 6454 12832 6460 12844
rect 6043 12804 6460 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 4982 12764 4988 12776
rect 3344 12736 4988 12764
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 6012 12764 6040 12795
rect 6454 12792 6460 12804
rect 6512 12832 6518 12844
rect 6512 12804 6592 12832
rect 6512 12792 6518 12804
rect 5408 12736 6040 12764
rect 6365 12767 6423 12773
rect 5408 12724 5414 12736
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6564 12764 6592 12804
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 7282 12832 7288 12844
rect 7064 12804 7288 12832
rect 7064 12792 7070 12804
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 8202 12832 8208 12844
rect 7423 12804 8208 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7392 12764 7420 12795
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 9122 12832 9128 12844
rect 9083 12804 9128 12832
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12832 10103 12835
rect 10502 12832 10508 12844
rect 10091 12804 10508 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 10873 12835 10931 12841
rect 10873 12832 10885 12835
rect 10836 12804 10885 12832
rect 10836 12792 10842 12804
rect 10873 12801 10885 12804
rect 10919 12832 10931 12835
rect 11256 12832 11284 12872
rect 12360 12844 12388 12872
rect 12434 12860 12440 12912
rect 12492 12900 12498 12912
rect 13170 12900 13176 12912
rect 12492 12872 13176 12900
rect 12492 12860 12498 12872
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 13464 12900 13492 12940
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13998 12968 14004 12980
rect 13587 12940 14004 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14458 12900 14464 12912
rect 13464 12872 14464 12900
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 11606 12832 11612 12844
rect 10919 12804 11284 12832
rect 11567 12804 11612 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12400 12804 13001 12832
rect 12400 12792 12406 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 16942 12832 16948 12844
rect 15335 12804 16948 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 6564 12736 7420 12764
rect 9769 12767 9827 12773
rect 6365 12727 6423 12733
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 10594 12764 10600 12776
rect 9815 12736 10600 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 3510 12705 3516 12708
rect 3504 12696 3516 12705
rect 3068 12668 3516 12696
rect 3504 12659 3516 12668
rect 3510 12656 3516 12659
rect 3568 12656 3574 12708
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 5442 12696 5448 12708
rect 4764 12668 5448 12696
rect 4764 12656 4770 12668
rect 5442 12656 5448 12668
rect 5500 12696 5506 12708
rect 6178 12696 6184 12708
rect 5500 12668 6184 12696
rect 5500 12656 5506 12668
rect 6178 12656 6184 12668
rect 6236 12656 6242 12708
rect 6380 12696 6408 12727
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 11425 12767 11483 12773
rect 11425 12733 11437 12767
rect 11471 12764 11483 12767
rect 12434 12764 12440 12776
rect 11471 12736 12440 12764
rect 11471 12733 11483 12736
rect 11425 12727 11483 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12894 12764 12900 12776
rect 12807 12736 12900 12764
rect 12894 12724 12900 12736
rect 12952 12764 12958 12776
rect 13998 12764 14004 12776
rect 12952 12736 14004 12764
rect 12952 12724 12958 12736
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14844 12736 15025 12764
rect 7926 12696 7932 12708
rect 6380 12668 7932 12696
rect 7926 12656 7932 12668
rect 7984 12656 7990 12708
rect 8941 12699 8999 12705
rect 8941 12665 8953 12699
rect 8987 12696 8999 12699
rect 11517 12699 11575 12705
rect 8987 12668 10272 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2556 12600 2881 12628
rect 2556 12588 2562 12600
rect 2869 12597 2881 12600
rect 2915 12628 2927 12631
rect 3602 12628 3608 12640
rect 2915 12600 3608 12628
rect 2915 12597 2927 12600
rect 2869 12591 2927 12597
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4617 12631 4675 12637
rect 4617 12628 4629 12631
rect 4212 12600 4629 12628
rect 4212 12588 4218 12600
rect 4617 12597 4629 12600
rect 4663 12597 4675 12631
rect 4617 12591 4675 12597
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 6638 12628 6644 12640
rect 5767 12600 6644 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 6825 12631 6883 12637
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 6914 12628 6920 12640
rect 6871 12600 6920 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7190 12628 7196 12640
rect 7151 12600 7196 12628
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 7524 12600 7665 12628
rect 7524 12588 7530 12600
rect 7653 12597 7665 12600
rect 7699 12597 7711 12631
rect 8018 12628 8024 12640
rect 7979 12600 8024 12628
rect 7653 12591 7711 12597
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8846 12628 8852 12640
rect 8159 12600 8852 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9033 12631 9091 12637
rect 9033 12597 9045 12631
rect 9079 12628 9091 12631
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 9079 12600 9413 12628
rect 9079 12597 9091 12600
rect 9033 12591 9091 12597
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9858 12628 9864 12640
rect 9819 12600 9864 12628
rect 9401 12591 9459 12597
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10244 12637 10272 12668
rect 10612 12668 10916 12696
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12597 10287 12631
rect 10229 12591 10287 12597
rect 10410 12588 10416 12640
rect 10468 12628 10474 12640
rect 10612 12637 10640 12668
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10468 12600 10609 12628
rect 10468 12588 10474 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 10597 12591 10655 12597
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 10888 12628 10916 12668
rect 11517 12665 11529 12699
rect 11563 12696 11575 12699
rect 11563 12668 12480 12696
rect 11563 12665 11575 12668
rect 11517 12659 11575 12665
rect 12452 12637 12480 12668
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12802 12696 12808 12708
rect 12584 12668 12808 12696
rect 12584 12656 12590 12668
rect 12802 12656 12808 12668
rect 12860 12696 12866 12708
rect 13265 12699 13323 12705
rect 13265 12696 13277 12699
rect 12860 12668 13277 12696
rect 12860 12656 12866 12668
rect 13265 12665 13277 12668
rect 13311 12665 13323 12699
rect 13265 12659 13323 12665
rect 14844 12640 14872 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 10744 12600 10789 12628
rect 10888 12600 11897 12628
rect 10744 12588 10750 12600
rect 11885 12597 11897 12600
rect 11931 12597 11943 12631
rect 11885 12591 11943 12597
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12597 12495 12631
rect 12437 12591 12495 12597
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 12894 12628 12900 12640
rect 12676 12600 12900 12628
rect 12676 12588 12682 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 14826 12628 14832 12640
rect 14787 12600 14832 12628
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 1104 12538 16008 12560
rect 1104 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 10976 12538
rect 11028 12486 11040 12538
rect 11092 12486 11104 12538
rect 11156 12486 11168 12538
rect 11220 12486 16008 12538
rect 1104 12464 16008 12486
rect 3602 12424 3608 12436
rect 3563 12396 3608 12424
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 9861 12427 9919 12433
rect 6788 12396 8136 12424
rect 6788 12384 6794 12396
rect 2866 12356 2872 12368
rect 2148 12328 2872 12356
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12288 1547 12291
rect 2038 12288 2044 12300
rect 1535 12260 2044 12288
rect 1535 12257 1547 12260
rect 1489 12251 1547 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2148 12297 2176 12328
rect 2866 12316 2872 12328
rect 2924 12356 2930 12368
rect 3234 12356 3240 12368
rect 2924 12328 3240 12356
rect 2924 12316 2930 12328
rect 3234 12316 3240 12328
rect 3292 12316 3298 12368
rect 5068 12359 5126 12365
rect 5068 12325 5080 12359
rect 5114 12356 5126 12359
rect 5350 12356 5356 12368
rect 5114 12328 5356 12356
rect 5114 12325 5126 12328
rect 5068 12319 5126 12325
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 6270 12316 6276 12368
rect 6328 12356 6334 12368
rect 6454 12356 6460 12368
rect 6328 12328 6460 12356
rect 6328 12316 6334 12328
rect 6454 12316 6460 12328
rect 6512 12356 6518 12368
rect 6512 12328 7788 12356
rect 6512 12316 6518 12328
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12257 2191 12291
rect 2133 12251 2191 12257
rect 2400 12291 2458 12297
rect 2400 12257 2412 12291
rect 2446 12288 2458 12291
rect 2774 12288 2780 12300
rect 2446 12260 2780 12288
rect 2446 12257 2458 12260
rect 2400 12251 2458 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 4617 12291 4675 12297
rect 4617 12257 4629 12291
rect 4663 12288 4675 12291
rect 4706 12288 4712 12300
rect 4663 12260 4712 12288
rect 4663 12257 4675 12260
rect 4617 12251 4675 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5810 12248 5816 12300
rect 5868 12288 5874 12300
rect 6540 12291 6598 12297
rect 6540 12288 6552 12291
rect 5868 12260 6552 12288
rect 5868 12248 5874 12260
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 4801 12223 4859 12229
rect 3292 12192 4108 12220
rect 3292 12180 3298 12192
rect 3510 12152 3516 12164
rect 3471 12124 3516 12152
rect 3510 12112 3516 12124
rect 3568 12112 3574 12164
rect 4080 12096 4108 12192
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 4120 12056 4445 12084
rect 4120 12044 4126 12056
rect 4433 12053 4445 12056
rect 4479 12084 4491 12087
rect 4816 12084 4844 12183
rect 6196 12161 6224 12260
rect 6540 12257 6552 12260
rect 6586 12288 6598 12291
rect 7098 12288 7104 12300
rect 6586 12260 7104 12288
rect 6586 12257 6598 12260
rect 6540 12251 6598 12257
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7760 12297 7788 12328
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12257 7803 12291
rect 8001 12291 8059 12297
rect 8001 12288 8013 12291
rect 7745 12251 7803 12257
rect 7852 12260 8013 12288
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 7852 12220 7880 12260
rect 8001 12257 8013 12260
rect 8047 12257 8059 12291
rect 8108 12288 8136 12396
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 10686 12424 10692 12436
rect 9907 12396 10692 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 12069 12427 12127 12433
rect 12069 12393 12081 12427
rect 12115 12424 12127 12427
rect 12342 12424 12348 12436
rect 12115 12396 12348 12424
rect 12115 12393 12127 12396
rect 12069 12387 12127 12393
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 9030 12316 9036 12368
rect 9088 12356 9094 12368
rect 9950 12356 9956 12368
rect 9088 12328 9956 12356
rect 9088 12316 9094 12328
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 10229 12359 10287 12365
rect 10229 12325 10241 12359
rect 10275 12356 10287 12359
rect 11974 12356 11980 12368
rect 10275 12328 11980 12356
rect 10275 12325 10287 12328
rect 10229 12319 10287 12325
rect 10244 12288 10272 12319
rect 11974 12316 11980 12328
rect 12032 12356 12038 12368
rect 12621 12359 12679 12365
rect 12621 12356 12633 12359
rect 12032 12328 12633 12356
rect 12032 12316 12038 12328
rect 12621 12325 12633 12328
rect 12667 12325 12679 12359
rect 12621 12319 12679 12325
rect 10962 12297 10968 12300
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 8108 12260 10272 12288
rect 10612 12260 10701 12288
rect 8001 12251 8059 12257
rect 6328 12192 6373 12220
rect 7668 12192 7880 12220
rect 6328 12180 6334 12192
rect 6181 12155 6239 12161
rect 6181 12121 6193 12155
rect 6227 12121 6239 12155
rect 6181 12115 6239 12121
rect 6086 12084 6092 12096
rect 4479 12056 6092 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 6270 12044 6276 12096
rect 6328 12084 6334 12096
rect 7668 12093 7696 12192
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 9950 12220 9956 12232
rect 9732 12192 9956 12220
rect 9732 12180 9738 12192
rect 9950 12180 9956 12192
rect 10008 12220 10014 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10008 12192 10333 12220
rect 10008 12180 10014 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12189 10563 12223
rect 10505 12183 10563 12189
rect 9125 12155 9183 12161
rect 9125 12121 9137 12155
rect 9171 12152 9183 12155
rect 9171 12124 10364 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 7653 12087 7711 12093
rect 7653 12084 7665 12087
rect 6328 12056 7665 12084
rect 6328 12044 6334 12056
rect 7653 12053 7665 12056
rect 7699 12053 7711 12087
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 7653 12047 7711 12053
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10134 12084 10140 12096
rect 9732 12056 10140 12084
rect 9732 12044 9738 12056
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 10336 12084 10364 12124
rect 10410 12084 10416 12096
rect 10323 12056 10416 12084
rect 10410 12044 10416 12056
rect 10468 12084 10474 12096
rect 10520 12084 10548 12183
rect 10468 12056 10548 12084
rect 10612 12084 10640 12260
rect 10689 12257 10701 12260
rect 10735 12257 10747 12291
rect 10956 12288 10968 12297
rect 10923 12260 10968 12288
rect 10689 12251 10747 12257
rect 10956 12251 10968 12260
rect 10962 12248 10968 12251
rect 11020 12248 11026 12300
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13814 12288 13820 12300
rect 13127 12260 13820 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13814 12248 13820 12260
rect 13872 12288 13878 12300
rect 14826 12288 14832 12300
rect 13872 12260 14832 12288
rect 13872 12248 13878 12260
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12220 12219 12223
rect 12618 12220 12624 12232
rect 12207 12192 12624 12220
rect 12207 12189 12219 12192
rect 12161 12183 12219 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 11330 12084 11336 12096
rect 10612 12056 11336 12084
rect 10468 12044 10474 12056
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 12437 12087 12495 12093
rect 12437 12084 12449 12087
rect 12308 12056 12449 12084
rect 12308 12044 12314 12056
rect 12437 12053 12449 12056
rect 12483 12053 12495 12087
rect 12437 12047 12495 12053
rect 1104 11994 16008 12016
rect 1104 11942 3480 11994
rect 3532 11942 3544 11994
rect 3596 11942 3608 11994
rect 3660 11942 3672 11994
rect 3724 11942 8478 11994
rect 8530 11942 8542 11994
rect 8594 11942 8606 11994
rect 8658 11942 8670 11994
rect 8722 11942 13475 11994
rect 13527 11942 13539 11994
rect 13591 11942 13603 11994
rect 13655 11942 13667 11994
rect 13719 11942 16008 11994
rect 1104 11920 16008 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2832 11852 2877 11880
rect 2832 11840 2838 11852
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 3844 11852 4077 11880
rect 3844 11840 3850 11852
rect 4065 11849 4077 11852
rect 4111 11880 4123 11883
rect 4338 11880 4344 11892
rect 4111 11852 4344 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4982 11880 4988 11892
rect 4943 11852 4988 11880
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 7926 11880 7932 11892
rect 5092 11852 7512 11880
rect 7887 11852 7932 11880
rect 3878 11772 3884 11824
rect 3936 11812 3942 11824
rect 5092 11812 5120 11852
rect 3936 11784 5120 11812
rect 3936 11772 3942 11784
rect 5718 11772 5724 11824
rect 5776 11812 5782 11824
rect 5776 11784 6408 11812
rect 5776 11772 5782 11784
rect 4706 11744 4712 11756
rect 2976 11716 4712 11744
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2866 11676 2872 11688
rect 1443 11648 2872 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 2976 11620 3004 11716
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5224 11716 5457 11744
rect 5224 11704 5230 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11744 5687 11747
rect 6270 11744 6276 11756
rect 5675 11716 6276 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 6380 11753 6408 11784
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 7484 11812 7512 11852
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 10594 11880 10600 11892
rect 9732 11852 9777 11880
rect 10555 11852 10600 11880
rect 9732 11840 9738 11852
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 11701 11883 11759 11889
rect 11701 11880 11713 11883
rect 11480 11852 11713 11880
rect 11480 11840 11486 11852
rect 11701 11849 11713 11852
rect 11747 11849 11759 11883
rect 11701 11843 11759 11849
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 13541 11883 13599 11889
rect 12492 11852 12537 11880
rect 12492 11840 12498 11852
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 13814 11880 13820 11892
rect 13587 11852 13820 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 9490 11812 9496 11824
rect 7156 11784 7420 11812
rect 7484 11784 9496 11812
rect 7156 11772 7162 11784
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7392 11753 7420 11784
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 6972 11716 7297 11744
rect 6972 11704 6978 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 8018 11744 8024 11756
rect 7699 11716 8024 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 9214 11744 9220 11756
rect 9175 11716 9220 11744
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 9692 11744 9720 11840
rect 9769 11815 9827 11821
rect 9769 11781 9781 11815
rect 9815 11812 9827 11815
rect 9858 11812 9864 11824
rect 9815 11784 9864 11812
rect 9815 11781 9827 11784
rect 9769 11775 9827 11781
rect 9858 11772 9864 11784
rect 9916 11772 9922 11824
rect 10226 11744 10232 11756
rect 9692 11716 10232 11744
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 10410 11744 10416 11756
rect 10371 11716 10416 11744
rect 10410 11704 10416 11716
rect 10468 11744 10474 11756
rect 10962 11744 10968 11756
rect 10468 11716 10968 11744
rect 10468 11704 10474 11716
rect 10962 11704 10968 11716
rect 11020 11744 11026 11756
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 11020 11716 11161 11744
rect 11020 11704 11026 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12400 11716 13001 11744
rect 12400 11704 12406 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 7193 11679 7251 11685
rect 5399 11648 6868 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 1664 11611 1722 11617
rect 1664 11577 1676 11611
rect 1710 11608 1722 11611
rect 2958 11608 2964 11620
rect 1710 11580 2964 11608
rect 1710 11577 1722 11580
rect 1664 11571 1722 11577
rect 2958 11568 2964 11580
rect 3016 11568 3022 11620
rect 4525 11611 4583 11617
rect 4525 11577 4537 11611
rect 4571 11608 4583 11611
rect 4571 11580 5212 11608
rect 4571 11577 4583 11580
rect 4525 11571 4583 11577
rect 4154 11540 4160 11552
rect 4115 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 5184 11540 5212 11580
rect 5626 11568 5632 11620
rect 5684 11608 5690 11620
rect 6181 11611 6239 11617
rect 6181 11608 6193 11611
rect 5684 11580 6193 11608
rect 5684 11568 5690 11580
rect 6181 11577 6193 11580
rect 6227 11577 6239 11611
rect 6181 11571 6239 11577
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 4672 11512 4717 11540
rect 5184 11512 5825 11540
rect 4672 11500 4678 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 6270 11540 6276 11552
rect 6231 11512 6276 11540
rect 5813 11503 5871 11509
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6840 11549 6868 11648
rect 7193 11645 7205 11679
rect 7239 11676 7251 11679
rect 7466 11676 7472 11688
rect 7239 11648 7472 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 8110 11676 8116 11688
rect 8071 11648 8116 11676
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10778 11676 10784 11688
rect 10100 11648 10784 11676
rect 10100 11636 10106 11648
rect 10778 11636 10784 11648
rect 10836 11676 10842 11688
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10836 11648 11069 11676
rect 10836 11636 10842 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11422 11636 11428 11688
rect 11480 11636 11486 11688
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 11698 11676 11704 11688
rect 11655 11648 11704 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12676 11648 12817 11676
rect 12676 11636 12682 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 9033 11611 9091 11617
rect 9033 11577 9045 11611
rect 9079 11608 9091 11611
rect 9674 11608 9680 11620
rect 9079 11580 9680 11608
rect 9079 11577 9091 11580
rect 9033 11571 9091 11577
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 10965 11611 11023 11617
rect 10965 11577 10977 11611
rect 11011 11608 11023 11611
rect 11440 11608 11468 11636
rect 11011 11580 11468 11608
rect 11011 11577 11023 11580
rect 10965 11571 11023 11577
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 6972 11512 8677 11540
rect 6972 11500 6978 11512
rect 8665 11509 8677 11512
rect 8711 11509 8723 11543
rect 8665 11503 8723 11509
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 9180 11512 9225 11540
rect 9180 11500 9186 11512
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9858 11540 9864 11552
rect 9548 11512 9864 11540
rect 9548 11500 9554 11512
rect 9858 11500 9864 11512
rect 9916 11540 9922 11552
rect 10137 11543 10195 11549
rect 10137 11540 10149 11543
rect 9916 11512 10149 11540
rect 9916 11500 9922 11512
rect 10137 11509 10149 11512
rect 10183 11509 10195 11543
rect 10137 11503 10195 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11425 11543 11483 11549
rect 11425 11540 11437 11543
rect 11388 11512 11437 11540
rect 11388 11500 11394 11512
rect 11425 11509 11437 11512
rect 11471 11509 11483 11543
rect 11425 11503 11483 11509
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 12342 11540 12348 11552
rect 12124 11512 12348 11540
rect 12124 11500 12130 11512
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 12943 11512 13369 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13357 11509 13369 11512
rect 13403 11540 13415 11543
rect 14182 11540 14188 11552
rect 13403 11512 14188 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 14182 11500 14188 11512
rect 14240 11540 14246 11552
rect 15746 11540 15752 11552
rect 14240 11512 15752 11540
rect 14240 11500 14246 11512
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 1104 11450 16008 11472
rect 1104 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 10976 11450
rect 11028 11398 11040 11450
rect 11092 11398 11104 11450
rect 11156 11398 11168 11450
rect 11220 11398 16008 11450
rect 1104 11376 16008 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 4154 11336 4160 11348
rect 2455 11308 4160 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 4764 11308 5457 11336
rect 4764 11296 4770 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5626 11336 5632 11348
rect 5587 11308 5632 11336
rect 5445 11299 5503 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 7006 11336 7012 11348
rect 6328 11308 7012 11336
rect 6328 11296 6334 11308
rect 7006 11296 7012 11308
rect 7064 11336 7070 11348
rect 7561 11339 7619 11345
rect 7561 11336 7573 11339
rect 7064 11308 7573 11336
rect 7064 11296 7070 11308
rect 7561 11305 7573 11308
rect 7607 11336 7619 11339
rect 7742 11336 7748 11348
rect 7607 11308 7748 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8297 11339 8355 11345
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 9766 11336 9772 11348
rect 8343 11308 9772 11336
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10468 11308 10517 11336
rect 10468 11296 10474 11308
rect 10505 11305 10517 11308
rect 10551 11336 10563 11339
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 10551 11308 11437 11336
rect 10551 11305 10563 11308
rect 10505 11299 10563 11305
rect 11425 11305 11437 11308
rect 11471 11336 11483 11339
rect 11514 11336 11520 11348
rect 11471 11308 11520 11336
rect 11471 11305 11483 11308
rect 11425 11299 11483 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 3513 11271 3571 11277
rect 3513 11237 3525 11271
rect 3559 11268 3571 11271
rect 3786 11268 3792 11280
rect 3559 11240 3792 11268
rect 3559 11237 3571 11240
rect 3513 11231 3571 11237
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 6454 11268 6460 11280
rect 6012 11240 6460 11268
rect 4332 11203 4390 11209
rect 4332 11200 4344 11203
rect 3804 11172 4344 11200
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 2774 11132 2780 11144
rect 2731 11104 2780 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 3804 11141 3832 11172
rect 4332 11169 4344 11172
rect 4378 11200 4390 11203
rect 5718 11200 5724 11212
rect 4378 11172 5724 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6012 11209 6040 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 6822 11268 6828 11280
rect 6604 11240 6828 11268
rect 6604 11228 6610 11240
rect 6822 11228 6828 11240
rect 6880 11228 6886 11280
rect 8389 11271 8447 11277
rect 8389 11237 8401 11271
rect 8435 11268 8447 11271
rect 9030 11268 9036 11280
rect 8435 11240 9036 11268
rect 8435 11237 8447 11240
rect 8389 11231 8447 11237
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 10870 11268 10876 11280
rect 9968 11240 10876 11268
rect 5997 11203 6055 11209
rect 5997 11169 6009 11203
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 6264 11203 6322 11209
rect 6264 11169 6276 11203
rect 6310 11200 6322 11203
rect 7558 11200 7564 11212
rect 6310 11172 7564 11200
rect 6310 11169 6322 11172
rect 6264 11163 6322 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 8846 11160 8852 11212
rect 8904 11200 8910 11212
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 8904 11172 9137 11200
rect 8904 11160 8910 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 9968 11200 9996 11240
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 11241 11271 11299 11277
rect 11241 11237 11253 11271
rect 11287 11268 11299 11271
rect 12066 11268 12072 11280
rect 11287 11240 12072 11268
rect 11287 11237 11299 11240
rect 11241 11231 11299 11237
rect 9263 11172 9996 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 3384 11104 3617 11132
rect 3384 11092 3390 11104
rect 3605 11101 3617 11104
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 4062 11132 4068 11144
rect 4023 11104 4068 11132
rect 3789 11095 3847 11101
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 3804 11064 3832 11095
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 7377 11067 7435 11073
rect 7377 11064 7389 11067
rect 3292 11036 3832 11064
rect 6932 11036 7389 11064
rect 3292 11024 3298 11036
rect 3050 10956 3056 11008
rect 3108 10996 3114 11008
rect 3145 10999 3203 11005
rect 3145 10996 3157 10999
rect 3108 10968 3157 10996
rect 3108 10956 3114 10968
rect 3145 10965 3157 10968
rect 3191 10965 3203 10999
rect 3145 10959 3203 10965
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 6932 10996 6960 11036
rect 7377 11033 7389 11036
rect 7423 11033 7435 11067
rect 8496 11064 8524 11095
rect 9416 11064 9444 11095
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 9968 11141 9996 11172
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 11256 11200 11284 11231
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 10643 11172 11284 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 11388 11172 11713 11200
rect 11388 11160 11394 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 11968 11203 12026 11209
rect 11968 11169 11980 11203
rect 12014 11200 12026 11203
rect 12250 11200 12256 11212
rect 12014 11172 12256 11200
rect 12014 11169 12026 11172
rect 11968 11163 12026 11169
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 10042 11132 10048 11144
rect 9999 11104 10048 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 11422 11132 11428 11144
rect 10928 11104 11428 11132
rect 10928 11092 10934 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 8496 11036 9444 11064
rect 7377 11027 7435 11033
rect 6696 10968 6960 10996
rect 6696 10956 6702 10968
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 7929 10999 7987 11005
rect 7929 10996 7941 10999
rect 7708 10968 7941 10996
rect 7708 10956 7714 10968
rect 7929 10965 7941 10968
rect 7975 10965 7987 10999
rect 7929 10959 7987 10965
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8757 10999 8815 11005
rect 8757 10996 8769 10999
rect 8076 10968 8769 10996
rect 8076 10956 8082 10968
rect 8757 10965 8769 10968
rect 8803 10965 8815 10999
rect 9416 10996 9444 11036
rect 9677 11067 9735 11073
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 9784 11064 9812 11092
rect 10134 11064 10140 11076
rect 9723 11036 9996 11064
rect 10095 11036 10140 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 9766 10996 9772 11008
rect 9416 10968 9772 10996
rect 8757 10959 8815 10965
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 9968 10996 9996 11036
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10778 11024 10784 11076
rect 10836 11064 10842 11076
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 10836 11036 10977 11064
rect 10836 11024 10842 11036
rect 10965 11033 10977 11036
rect 11011 11033 11023 11067
rect 10965 11027 11023 11033
rect 12434 10996 12440 11008
rect 9968 10968 12440 10996
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 13081 10999 13139 11005
rect 13081 10996 13093 10999
rect 12676 10968 13093 10996
rect 12676 10956 12682 10968
rect 13081 10965 13093 10968
rect 13127 10965 13139 10999
rect 16114 10996 16120 11008
rect 16075 10968 16120 10996
rect 13081 10959 13139 10965
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 1104 10906 16008 10928
rect 1104 10854 3480 10906
rect 3532 10854 3544 10906
rect 3596 10854 3608 10906
rect 3660 10854 3672 10906
rect 3724 10854 8478 10906
rect 8530 10854 8542 10906
rect 8594 10854 8606 10906
rect 8658 10854 8670 10906
rect 8722 10854 13475 10906
rect 13527 10854 13539 10906
rect 13591 10854 13603 10906
rect 13655 10854 13667 10906
rect 13719 10854 16008 10906
rect 1104 10832 16008 10854
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3421 10795 3479 10801
rect 3421 10792 3433 10795
rect 3384 10764 3433 10792
rect 3384 10752 3390 10764
rect 3421 10761 3433 10764
rect 3467 10761 3479 10795
rect 5905 10795 5963 10801
rect 5905 10792 5917 10795
rect 3421 10755 3479 10761
rect 3988 10764 5917 10792
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 3234 10656 3240 10668
rect 3195 10628 3240 10656
rect 3234 10616 3240 10628
rect 3292 10616 3298 10668
rect 3878 10656 3884 10668
rect 3839 10628 3884 10656
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10588 1547 10591
rect 3988 10588 4016 10764
rect 5905 10761 5917 10764
rect 5951 10761 5963 10795
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 5905 10755 5963 10761
rect 6012 10764 11529 10792
rect 5629 10727 5687 10733
rect 5629 10693 5641 10727
rect 5675 10724 5687 10727
rect 5718 10724 5724 10736
rect 5675 10696 5724 10724
rect 5675 10693 5687 10696
rect 5629 10687 5687 10693
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 6012 10724 6040 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 12308 10764 14105 10792
rect 12308 10752 12314 10764
rect 14093 10761 14105 10764
rect 14139 10761 14151 10795
rect 14093 10755 14151 10761
rect 9214 10724 9220 10736
rect 5868 10696 6040 10724
rect 8864 10696 9220 10724
rect 5868 10684 5874 10696
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 1535 10560 4016 10588
rect 1535 10557 1547 10560
rect 1489 10551 1547 10557
rect 2961 10523 3019 10529
rect 2961 10489 2973 10523
rect 3007 10520 3019 10523
rect 3510 10520 3516 10532
rect 3007 10492 3516 10520
rect 3007 10489 3019 10492
rect 2961 10483 3019 10489
rect 3510 10480 3516 10492
rect 3568 10480 3574 10532
rect 4080 10520 4108 10619
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4212 10628 4261 10656
rect 4212 10616 4218 10628
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4249 10619 4307 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6638 10656 6644 10668
rect 6595 10628 6644 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6638 10616 6644 10628
rect 6696 10616 6702 10668
rect 7558 10656 7564 10668
rect 7519 10628 7564 10656
rect 7558 10616 7564 10628
rect 7616 10656 7622 10668
rect 7616 10628 7972 10656
rect 7616 10616 7622 10628
rect 6365 10591 6423 10597
rect 6365 10557 6377 10591
rect 6411 10588 6423 10591
rect 6914 10588 6920 10600
rect 6411 10560 6920 10588
rect 6411 10557 6423 10560
rect 6365 10551 6423 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7650 10588 7656 10600
rect 7515 10560 7656 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 7834 10588 7840 10600
rect 7795 10560 7840 10588
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 7944 10588 7972 10628
rect 8864 10588 8892 10696
rect 9214 10684 9220 10696
rect 9272 10684 9278 10736
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 9088 10628 9321 10656
rect 9088 10616 9094 10628
rect 9309 10625 9321 10628
rect 9355 10656 9367 10659
rect 9490 10656 9496 10668
rect 9355 10628 9496 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12618 10656 12624 10668
rect 12207 10628 12624 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 7944 10560 8892 10588
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9858 10588 9864 10600
rect 9723 10560 9864 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10588 10103 10591
rect 11330 10588 11336 10600
rect 10091 10560 11336 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 4516 10523 4574 10529
rect 4516 10520 4528 10523
rect 4080 10492 4528 10520
rect 4516 10489 4528 10492
rect 4562 10520 4574 10523
rect 5166 10520 5172 10532
rect 4562 10492 5172 10520
rect 4562 10489 4574 10492
rect 4516 10483 4574 10489
rect 5166 10480 5172 10492
rect 5224 10480 5230 10532
rect 6273 10523 6331 10529
rect 6273 10489 6285 10523
rect 6319 10520 6331 10523
rect 8104 10523 8162 10529
rect 6319 10492 7052 10520
rect 6319 10489 6331 10492
rect 6273 10483 6331 10489
rect 2590 10452 2596 10464
rect 2551 10424 2596 10452
rect 2590 10412 2596 10424
rect 2648 10412 2654 10464
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 3602 10452 3608 10464
rect 3099 10424 3608 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 3789 10455 3847 10461
rect 3789 10421 3801 10455
rect 3835 10452 3847 10455
rect 4338 10452 4344 10464
rect 3835 10424 4344 10452
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 7024 10461 7052 10492
rect 8104 10489 8116 10523
rect 8150 10520 8162 10523
rect 8150 10492 8708 10520
rect 8150 10489 8162 10492
rect 8104 10483 8162 10489
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10421 7067 10455
rect 7009 10415 7067 10421
rect 7377 10455 7435 10461
rect 7377 10421 7389 10455
rect 7423 10452 7435 10455
rect 7926 10452 7932 10464
rect 7423 10424 7932 10452
rect 7423 10421 7435 10424
rect 7377 10415 7435 10421
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 8680 10452 8708 10492
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 10060 10520 10088 10551
rect 11330 10548 11336 10560
rect 11388 10588 11394 10600
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 11388 10560 12725 10588
rect 11388 10548 11394 10560
rect 12713 10557 12725 10560
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 8812 10492 10088 10520
rect 10312 10523 10370 10529
rect 8812 10480 8818 10492
rect 10312 10489 10324 10523
rect 10358 10520 10370 10523
rect 10686 10520 10692 10532
rect 10358 10492 10692 10520
rect 10358 10489 10370 10492
rect 10312 10483 10370 10489
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 11885 10523 11943 10529
rect 11885 10489 11897 10523
rect 11931 10520 11943 10523
rect 12802 10520 12808 10532
rect 11931 10492 12808 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 12986 10529 12992 10532
rect 12980 10483 12992 10529
rect 13044 10520 13050 10532
rect 13044 10492 13080 10520
rect 12986 10480 12992 10483
rect 13044 10480 13050 10492
rect 9766 10452 9772 10464
rect 8680 10424 9772 10452
rect 9766 10412 9772 10424
rect 9824 10452 9830 10464
rect 11425 10455 11483 10461
rect 11425 10452 11437 10455
rect 9824 10424 11437 10452
rect 9824 10412 9830 10424
rect 11425 10421 11437 10424
rect 11471 10421 11483 10455
rect 11974 10452 11980 10464
rect 11935 10424 11980 10452
rect 11425 10415 11483 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12894 10452 12900 10464
rect 12492 10424 12900 10452
rect 12492 10412 12498 10424
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 14734 10452 14740 10464
rect 14231 10424 14740 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 1104 10362 16008 10384
rect 1104 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 10976 10362
rect 11028 10310 11040 10362
rect 11092 10310 11104 10362
rect 11156 10310 11168 10362
rect 11220 10310 16008 10362
rect 1104 10288 16008 10310
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 2961 10251 3019 10257
rect 2961 10248 2973 10251
rect 2648 10220 2973 10248
rect 2648 10208 2654 10220
rect 2961 10217 2973 10220
rect 3007 10217 3019 10251
rect 2961 10211 3019 10217
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3602 10248 3608 10260
rect 3108 10220 3153 10248
rect 3563 10220 3608 10248
rect 3108 10208 3114 10220
rect 3602 10208 3608 10220
rect 3660 10248 3666 10260
rect 3970 10248 3976 10260
rect 3660 10220 3976 10248
rect 3660 10208 3666 10220
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 4672 10220 5089 10248
rect 4672 10208 4678 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 5077 10211 5135 10217
rect 5166 10208 5172 10260
rect 5224 10248 5230 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 5224 10220 7297 10248
rect 5224 10208 5230 10220
rect 7285 10217 7297 10220
rect 7331 10217 7343 10251
rect 7285 10211 7343 10217
rect 7377 10251 7435 10257
rect 7377 10217 7389 10251
rect 7423 10248 7435 10251
rect 8846 10248 8852 10260
rect 7423 10220 8852 10248
rect 7423 10217 7435 10220
rect 7377 10211 7435 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 13078 10248 13084 10260
rect 9539 10220 13084 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 13078 10208 13084 10220
rect 13136 10248 13142 10260
rect 14001 10251 14059 10257
rect 14001 10248 14013 10251
rect 13136 10220 14013 10248
rect 13136 10208 13142 10220
rect 14001 10217 14013 10220
rect 14047 10217 14059 10251
rect 14734 10248 14740 10260
rect 14695 10220 14740 10248
rect 14001 10211 14059 10217
rect 5810 10180 5816 10192
rect 1504 10152 5816 10180
rect 1504 10121 1532 10152
rect 5810 10140 5816 10152
rect 5868 10140 5874 10192
rect 6172 10183 6230 10189
rect 6172 10149 6184 10183
rect 6218 10180 6230 10183
rect 6638 10180 6644 10192
rect 6218 10152 6644 10180
rect 6218 10149 6230 10152
rect 6172 10143 6230 10149
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 7653 10183 7711 10189
rect 7653 10149 7665 10183
rect 7699 10180 7711 10183
rect 11692 10183 11750 10189
rect 7699 10152 10456 10180
rect 7699 10149 7711 10152
rect 7653 10143 7711 10149
rect 1499 10115 1557 10121
rect 1499 10081 1511 10115
rect 1545 10081 1557 10115
rect 1499 10075 1557 10081
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3936 10084 4261 10112
rect 3936 10072 3942 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4396 10084 4537 10112
rect 4396 10072 4402 10084
rect 4525 10081 4537 10084
rect 4571 10112 4583 10115
rect 5166 10112 5172 10124
rect 4571 10084 5172 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5442 10072 5448 10084
rect 5500 10112 5506 10124
rect 5626 10112 5632 10124
rect 5500 10084 5632 10112
rect 5500 10072 5506 10084
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6454 10112 6460 10124
rect 5951 10084 6460 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6454 10072 6460 10084
rect 6512 10072 6518 10124
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7926 10112 7932 10124
rect 7156 10084 7932 10112
rect 7156 10072 7162 10084
rect 7926 10072 7932 10084
rect 7984 10112 7990 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 7984 10084 9505 10112
rect 7984 10072 7990 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9858 10072 9864 10124
rect 9916 10112 9922 10124
rect 10318 10112 10324 10124
rect 9916 10084 10324 10112
rect 9916 10072 9922 10084
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10428 10112 10456 10152
rect 11692 10149 11704 10183
rect 11738 10180 11750 10183
rect 12618 10180 12624 10192
rect 11738 10152 12624 10180
rect 11738 10149 11750 10152
rect 11692 10143 11750 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 14016 10180 14044 10211
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 15289 10183 15347 10189
rect 15289 10180 15301 10183
rect 14016 10152 15301 10180
rect 15289 10149 15301 10152
rect 15335 10149 15347 10183
rect 15289 10143 15347 10149
rect 13262 10112 13268 10124
rect 10428 10084 13268 10112
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 13909 10115 13967 10121
rect 13909 10112 13921 10115
rect 13872 10084 13921 10112
rect 13872 10072 13878 10084
rect 13909 10081 13921 10084
rect 13955 10081 13967 10115
rect 14829 10115 14887 10121
rect 14829 10112 14841 10115
rect 13909 10075 13967 10081
rect 14016 10084 14841 10112
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3145 10047 3203 10053
rect 3145 10044 3157 10047
rect 3016 10016 3157 10044
rect 3016 10004 3022 10016
rect 3145 10013 3157 10016
rect 3191 10013 3203 10047
rect 5534 10044 5540 10056
rect 5495 10016 5540 10044
rect 3145 10007 3203 10013
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5718 10044 5724 10056
rect 5679 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 2498 9936 2504 9988
rect 2556 9976 2562 9988
rect 2593 9979 2651 9985
rect 2593 9976 2605 9979
rect 2556 9948 2605 9976
rect 2556 9936 2562 9948
rect 2593 9945 2605 9948
rect 2639 9945 2651 9979
rect 3510 9976 3516 9988
rect 3423 9948 3516 9976
rect 2593 9939 2651 9945
rect 3510 9936 3516 9948
rect 3568 9976 3574 9988
rect 5258 9976 5264 9988
rect 3568 9948 5264 9976
rect 3568 9936 3574 9948
rect 5258 9936 5264 9948
rect 5316 9976 5322 9988
rect 8202 9976 8208 9988
rect 5316 9948 5948 9976
rect 5316 9936 5322 9948
rect 5920 9908 5948 9948
rect 6840 9948 8208 9976
rect 6840 9908 6868 9948
rect 8202 9936 8208 9948
rect 8260 9936 8266 9988
rect 9861 9979 9919 9985
rect 9861 9945 9873 9979
rect 9907 9976 9919 9979
rect 10226 9976 10232 9988
rect 9907 9948 10232 9976
rect 9907 9945 9919 9948
rect 9861 9939 9919 9945
rect 10226 9936 10232 9948
rect 10284 9976 10290 9988
rect 10428 9976 10456 10007
rect 10284 9948 10456 9976
rect 10284 9936 10290 9948
rect 5920 9880 6868 9908
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 8110 9908 8116 9920
rect 7616 9880 8116 9908
rect 7616 9868 7622 9880
rect 8110 9868 8116 9880
rect 8168 9908 8174 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8168 9880 8953 9908
rect 8168 9868 8174 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 9950 9908 9956 9920
rect 9911 9880 9956 9908
rect 8941 9871 8999 9877
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 10612 9908 10640 10007
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11388 10016 11437 10044
rect 11388 10004 11394 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 14016 10044 14044 10084
rect 14829 10081 14841 10084
rect 14875 10112 14887 10115
rect 15473 10115 15531 10121
rect 15473 10112 15485 10115
rect 14875 10084 15485 10112
rect 14875 10081 14887 10084
rect 14829 10075 14887 10081
rect 15473 10081 15485 10084
rect 15519 10112 15531 10115
rect 16117 10115 16175 10121
rect 16117 10112 16129 10115
rect 15519 10084 16129 10112
rect 15519 10081 15531 10084
rect 15473 10075 15531 10081
rect 16117 10081 16129 10084
rect 16163 10081 16175 10115
rect 16117 10075 16175 10081
rect 12676 10016 14044 10044
rect 14093 10047 14151 10053
rect 12676 10004 12682 10016
rect 14093 10013 14105 10047
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 12986 9936 12992 9988
rect 13044 9976 13050 9988
rect 13906 9976 13912 9988
rect 13044 9948 13912 9976
rect 13044 9936 13050 9948
rect 13906 9936 13912 9948
rect 13964 9976 13970 9988
rect 14108 9976 14136 10007
rect 14936 9976 14964 10007
rect 13964 9948 14964 9976
rect 13964 9936 13970 9948
rect 10686 9908 10692 9920
rect 10599 9880 10692 9908
rect 10686 9868 10692 9880
rect 10744 9908 10750 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 10744 9880 12817 9908
rect 10744 9868 10750 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 13354 9868 13360 9920
rect 13412 9908 13418 9920
rect 13541 9911 13599 9917
rect 13541 9908 13553 9911
rect 13412 9880 13553 9908
rect 13412 9868 13418 9880
rect 13541 9877 13553 9880
rect 13587 9877 13599 9911
rect 14366 9908 14372 9920
rect 14327 9880 14372 9908
rect 13541 9871 13599 9877
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 1104 9818 16008 9840
rect 1104 9766 3480 9818
rect 3532 9766 3544 9818
rect 3596 9766 3608 9818
rect 3660 9766 3672 9818
rect 3724 9766 8478 9818
rect 8530 9766 8542 9818
rect 8594 9766 8606 9818
rect 8658 9766 8670 9818
rect 8722 9766 13475 9818
rect 13527 9766 13539 9818
rect 13591 9766 13603 9818
rect 13655 9766 13667 9818
rect 13719 9766 16008 9818
rect 1104 9744 16008 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 7650 9704 7656 9716
rect 3936 9676 7656 9704
rect 3936 9664 3942 9676
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 11517 9707 11575 9713
rect 9232 9676 11008 9704
rect 9232 9648 9260 9676
rect 4154 9596 4160 9648
rect 4212 9636 4218 9648
rect 4522 9636 4528 9648
rect 4212 9608 4528 9636
rect 4212 9596 4218 9608
rect 4522 9596 4528 9608
rect 4580 9636 4586 9648
rect 8113 9639 8171 9645
rect 4580 9608 6040 9636
rect 4580 9596 4586 9608
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 5626 9568 5632 9580
rect 5408 9540 5632 9568
rect 5408 9528 5414 9540
rect 5626 9528 5632 9540
rect 5684 9568 5690 9580
rect 5905 9571 5963 9577
rect 5905 9568 5917 9571
rect 5684 9540 5917 9568
rect 5684 9528 5690 9540
rect 5905 9537 5917 9540
rect 5951 9537 5963 9571
rect 5905 9531 5963 9537
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 4430 9500 4436 9512
rect 3007 9472 4436 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 4798 9460 4804 9512
rect 4856 9500 4862 9512
rect 5258 9500 5264 9512
rect 4856 9472 5264 9500
rect 4856 9460 4862 9472
rect 5258 9460 5264 9472
rect 5316 9500 5322 9512
rect 5810 9500 5816 9512
rect 5316 9472 5816 9500
rect 5316 9460 5322 9472
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 6012 9500 6040 9608
rect 8113 9605 8125 9639
rect 8159 9636 8171 9639
rect 8941 9639 8999 9645
rect 8159 9608 8892 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 8665 9571 8723 9577
rect 8665 9568 8677 9571
rect 8352 9540 8677 9568
rect 8352 9528 8358 9540
rect 8665 9537 8677 9540
rect 8711 9537 8723 9571
rect 8864 9568 8892 9608
rect 8941 9605 8953 9639
rect 8987 9636 8999 9639
rect 9122 9636 9128 9648
rect 8987 9608 9128 9636
rect 8987 9605 8999 9608
rect 8941 9599 8999 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 9214 9596 9220 9648
rect 9272 9596 9278 9648
rect 9306 9596 9312 9648
rect 9364 9636 9370 9648
rect 9364 9608 10272 9636
rect 9364 9596 9370 9608
rect 9030 9568 9036 9580
rect 8864 9540 9036 9568
rect 8665 9531 8723 9537
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 9324 9568 9352 9596
rect 9140 9540 9352 9568
rect 9493 9571 9551 9577
rect 9140 9512 9168 9540
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 9766 9568 9772 9580
rect 9539 9540 9772 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 9907 9540 10180 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 6012 9472 8984 9500
rect 3228 9435 3286 9441
rect 3228 9401 3240 9435
rect 3274 9432 3286 9435
rect 4614 9432 4620 9444
rect 3274 9404 4620 9432
rect 3274 9401 3286 9404
rect 3228 9395 3286 9401
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 5534 9392 5540 9444
rect 5592 9432 5598 9444
rect 8481 9435 8539 9441
rect 5592 9404 6224 9432
rect 5592 9392 5598 9404
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 3844 9336 4353 9364
rect 3844 9324 3850 9336
rect 4341 9333 4353 9336
rect 4387 9333 4399 9367
rect 4341 9327 4399 9333
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5810 9364 5816 9376
rect 5031 9336 5816 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6196 9373 6224 9404
rect 8481 9401 8493 9435
rect 8527 9432 8539 9435
rect 8846 9432 8852 9444
rect 8527 9404 8852 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6822 9364 6828 9376
rect 6227 9336 6828 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 8570 9364 8576 9376
rect 8531 9336 8576 9364
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 8956 9364 8984 9472
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9950 9500 9956 9512
rect 9447 9472 9956 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 9309 9435 9367 9441
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 9355 9404 10088 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9950 9364 9956 9376
rect 8956 9336 9956 9364
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10060 9373 10088 9404
rect 10045 9367 10103 9373
rect 10045 9333 10057 9367
rect 10091 9333 10103 9367
rect 10152 9364 10180 9540
rect 10244 9432 10272 9608
rect 10778 9596 10784 9648
rect 10836 9596 10842 9648
rect 10980 9636 11008 9676
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11974 9704 11980 9716
rect 11563 9676 11980 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11974 9664 11980 9676
rect 12032 9664 12038 9716
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 12308 9676 13860 9704
rect 12308 9664 12314 9676
rect 12066 9636 12072 9648
rect 10980 9608 12072 9636
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 10686 9568 10692 9580
rect 10647 9540 10692 9568
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 10796 9568 10824 9596
rect 12161 9571 12219 9577
rect 10796 9540 11192 9568
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 10870 9500 10876 9512
rect 10459 9472 10876 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 10870 9460 10876 9472
rect 10928 9500 10934 9512
rect 11057 9503 11115 9509
rect 11057 9500 11069 9503
rect 10928 9472 11069 9500
rect 10928 9460 10934 9472
rect 11057 9469 11069 9472
rect 11103 9469 11115 9503
rect 11057 9463 11115 9469
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10244 9404 10977 9432
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 10502 9364 10508 9376
rect 10152 9336 10508 9364
rect 10045 9327 10103 9333
rect 10502 9324 10508 9336
rect 10560 9364 10566 9376
rect 11164 9364 11192 9540
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 12268 9568 12296 9664
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 13265 9639 13323 9645
rect 13265 9636 13277 9639
rect 12860 9608 13277 9636
rect 12860 9596 12866 9608
rect 13265 9605 13277 9608
rect 13311 9605 13323 9639
rect 13265 9599 13323 9605
rect 12986 9568 12992 9580
rect 12207 9540 12296 9568
rect 12947 9540 12992 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 13832 9577 13860 9676
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13412 9540 13737 9568
rect 13412 9528 13418 9540
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 13078 9500 13084 9512
rect 11931 9472 13084 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9500 13691 9503
rect 14366 9500 14372 9512
rect 13679 9472 14372 9500
rect 13679 9469 13691 9472
rect 13633 9463 13691 9469
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 12802 9432 12808 9444
rect 12763 9404 12808 9432
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 10560 9336 11192 9364
rect 11977 9367 12035 9373
rect 10560 9324 10566 9336
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12023 9336 12449 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12437 9327 12495 9333
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 13872 9336 14473 9364
rect 13872 9324 13878 9336
rect 14461 9333 14473 9336
rect 14507 9364 14519 9367
rect 16114 9364 16120 9376
rect 14507 9336 16120 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 1104 9274 16008 9296
rect 1104 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 10976 9274
rect 11028 9222 11040 9274
rect 11092 9222 11104 9274
rect 11156 9222 11168 9274
rect 11220 9222 16008 9274
rect 1104 9200 16008 9222
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2096 9132 5120 9160
rect 2096 9120 2102 9132
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 4678 9095 4736 9101
rect 4678 9092 4690 9095
rect 3844 9064 4690 9092
rect 3844 9052 3850 9064
rect 4678 9061 4690 9064
rect 4724 9061 4736 9095
rect 5092 9092 5120 9132
rect 5166 9120 5172 9172
rect 5224 9160 5230 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 5224 9132 7757 9160
rect 5224 9120 5230 9132
rect 7745 9129 7757 9132
rect 7791 9160 7803 9163
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 7791 9132 8401 9160
rect 7791 9129 7803 9132
rect 7745 9123 7803 9129
rect 8389 9129 8401 9132
rect 8435 9129 8447 9163
rect 8570 9160 8576 9172
rect 8531 9132 8576 9160
rect 8389 9123 8447 9129
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 9033 9163 9091 9169
rect 9033 9129 9045 9163
rect 9079 9160 9091 9163
rect 9122 9160 9128 9172
rect 9079 9132 9128 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 10686 9160 10692 9172
rect 10643 9132 10692 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 9858 9092 9864 9104
rect 5092 9064 9864 9092
rect 4678 9055 4736 9061
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 10045 9095 10103 9101
rect 10045 9061 10057 9095
rect 10091 9092 10103 9095
rect 10612 9092 10640 9123
rect 10686 9120 10692 9132
rect 10744 9160 10750 9172
rect 12158 9160 12164 9172
rect 10744 9132 12020 9160
rect 12119 9132 12164 9160
rect 10744 9120 10750 9132
rect 10091 9064 10640 9092
rect 10956 9095 11014 9101
rect 10091 9061 10103 9064
rect 10045 9055 10103 9061
rect 10956 9061 10968 9095
rect 11002 9092 11014 9095
rect 11146 9092 11152 9104
rect 11002 9064 11152 9092
rect 11002 9061 11014 9064
rect 10956 9055 11014 9061
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 11992 9092 12020 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 12894 9160 12900 9172
rect 12575 9132 12900 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 13136 9132 13369 9160
rect 13136 9120 13142 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 14090 9092 14096 9104
rect 11992 9064 14096 9092
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 4430 9024 4436 9036
rect 4391 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 9024 4494 9036
rect 6178 9033 6184 9036
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 4488 8996 5917 9024
rect 4488 8984 4494 8996
rect 5828 8968 5856 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 6172 9024 6184 9033
rect 6139 8996 6184 9024
rect 5905 8987 5963 8993
rect 6172 8987 6184 8996
rect 6178 8984 6184 8987
rect 6236 8984 6242 9036
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 7837 9027 7895 9033
rect 7837 9024 7849 9027
rect 7708 8996 7849 9024
rect 7708 8984 7714 8996
rect 7837 8993 7849 8996
rect 7883 9024 7895 9027
rect 8941 9027 8999 9033
rect 7883 8996 8340 9024
rect 7883 8993 7895 8996
rect 7837 8987 7895 8993
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 7098 8848 7104 8900
rect 7156 8888 7162 8900
rect 7285 8891 7343 8897
rect 7285 8888 7297 8891
rect 7156 8860 7297 8888
rect 7156 8848 7162 8860
rect 7285 8857 7297 8860
rect 7331 8888 7343 8891
rect 7944 8888 7972 8919
rect 7331 8860 7972 8888
rect 7331 8857 7343 8860
rect 7285 8851 7343 8857
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5776 8792 5825 8820
rect 5776 8780 5782 8792
rect 5813 8789 5825 8792
rect 5859 8820 5871 8823
rect 6178 8820 6184 8832
rect 5859 8792 6184 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 8312 8829 8340 8996
rect 8941 8993 8953 9027
rect 8987 9024 8999 9027
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8987 8996 9505 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 9493 8993 9505 8996
rect 9539 9024 9551 9027
rect 9582 9024 9588 9036
rect 9539 8996 9588 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 9582 8984 9588 8996
rect 9640 9024 9646 9036
rect 9640 8996 11744 9024
rect 9640 8984 9646 8996
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9180 8928 9225 8956
rect 9180 8916 9186 8928
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 9824 8928 10241 8956
rect 9824 8916 9830 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10686 8956 10692 8968
rect 10647 8928 10692 8956
rect 10229 8919 10287 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 9950 8888 9956 8900
rect 9732 8860 9956 8888
rect 9732 8848 9738 8860
rect 9950 8848 9956 8860
rect 10008 8848 10014 8900
rect 8297 8823 8355 8829
rect 8297 8789 8309 8823
rect 8343 8820 8355 8823
rect 9214 8820 9220 8832
rect 8343 8792 9220 8820
rect 8343 8789 8355 8792
rect 8297 8783 8355 8789
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10686 8820 10692 8832
rect 9824 8792 10692 8820
rect 9824 8780 9830 8792
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11716 8820 11744 8996
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12897 9027 12955 9033
rect 12897 9024 12909 9027
rect 12216 8996 12909 9024
rect 12216 8984 12222 8996
rect 12897 8993 12909 8996
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13725 9027 13783 9033
rect 13725 9024 13737 9027
rect 13412 8996 13737 9024
rect 13412 8984 13418 8996
rect 13725 8993 13737 8996
rect 13771 9024 13783 9027
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13771 8996 14197 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 11848 8928 12357 8956
rect 11848 8916 11854 8928
rect 12345 8925 12357 8928
rect 12391 8956 12403 8959
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12391 8928 13001 8956
rect 12391 8925 12403 8928
rect 12345 8919 12403 8925
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 12066 8888 12072 8900
rect 11979 8860 12072 8888
rect 12066 8848 12072 8860
rect 12124 8888 12130 8900
rect 13096 8888 13124 8919
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13228 8928 13829 8956
rect 13228 8916 13234 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 13964 8928 14009 8956
rect 13964 8916 13970 8928
rect 12124 8860 13124 8888
rect 12124 8848 12130 8860
rect 13814 8820 13820 8832
rect 11716 8792 13820 8820
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 1104 8730 16008 8752
rect 1104 8678 3480 8730
rect 3532 8678 3544 8730
rect 3596 8678 3608 8730
rect 3660 8678 3672 8730
rect 3724 8678 8478 8730
rect 8530 8678 8542 8730
rect 8594 8678 8606 8730
rect 8658 8678 8670 8730
rect 8722 8678 13475 8730
rect 13527 8678 13539 8730
rect 13591 8678 13603 8730
rect 13655 8678 13667 8730
rect 13719 8678 16008 8730
rect 1104 8656 16008 8678
rect 8938 8616 8944 8628
rect 1504 8588 8944 8616
rect 1504 8421 1532 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 10410 8616 10416 8628
rect 9640 8588 10416 8616
rect 9640 8576 9646 8588
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8616 11210 8628
rect 11422 8616 11428 8628
rect 11204 8588 11428 8616
rect 11204 8576 11210 8588
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 13170 8616 13176 8628
rect 11563 8588 13176 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 13964 8588 14381 8616
rect 13964 8576 13970 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 14369 8579 14427 8585
rect 5721 8551 5779 8557
rect 5721 8548 5733 8551
rect 3620 8520 5733 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2774 8480 2780 8492
rect 2363 8452 2780 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 1489 8415 1547 8421
rect 1489 8381 1501 8415
rect 1535 8381 1547 8415
rect 2038 8412 2044 8424
rect 1999 8384 2044 8412
rect 1489 8375 1547 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 3620 8421 3648 8520
rect 5721 8517 5733 8520
rect 5767 8517 5779 8551
rect 5721 8511 5779 8517
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 10704 8548 10732 8576
rect 11330 8548 11336 8560
rect 5868 8520 6868 8548
rect 10704 8520 11336 8548
rect 5868 8508 5874 8520
rect 3786 8480 3792 8492
rect 3747 8452 3792 8480
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 4614 8480 4620 8492
rect 4575 8452 4620 8480
rect 4614 8440 4620 8452
rect 4672 8480 4678 8492
rect 6840 8489 6868 8520
rect 11330 8508 11336 8520
rect 11388 8548 11394 8560
rect 11388 8520 13032 8548
rect 11388 8508 11394 8520
rect 5445 8483 5503 8489
rect 5445 8480 5457 8483
rect 4672 8452 5457 8480
rect 4672 8440 4678 8452
rect 5445 8449 5457 8452
rect 5491 8480 5503 8483
rect 6273 8483 6331 8489
rect 6273 8480 6285 8483
rect 5491 8452 6285 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 6273 8449 6285 8452
rect 6319 8449 6331 8483
rect 6273 8443 6331 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 6825 8443 6883 8449
rect 8220 8452 8953 8480
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 4706 8412 4712 8424
rect 3605 8375 3663 8381
rect 4448 8384 4712 8412
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 4448 8288 4476 8384
rect 4706 8372 4712 8384
rect 4764 8412 4770 8424
rect 4764 8384 5212 8412
rect 4764 8372 4770 8384
rect 4525 8347 4583 8353
rect 4525 8313 4537 8347
rect 4571 8344 4583 8347
rect 5074 8344 5080 8356
rect 4571 8316 5080 8344
rect 4571 8313 4583 8316
rect 4525 8307 4583 8313
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 3234 8276 3240 8288
rect 3195 8248 3240 8276
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 3697 8279 3755 8285
rect 3697 8245 3709 8279
rect 3743 8276 3755 8279
rect 4065 8279 4123 8285
rect 4065 8276 4077 8279
rect 3743 8248 4077 8276
rect 3743 8245 3755 8248
rect 3697 8239 3755 8245
rect 4065 8245 4077 8248
rect 4111 8245 4123 8279
rect 4430 8276 4436 8288
rect 4391 8248 4436 8276
rect 4065 8239 4123 8245
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 4890 8276 4896 8288
rect 4851 8248 4896 8276
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5184 8276 5212 8384
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 5316 8384 5361 8412
rect 5316 8372 5322 8384
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 6089 8415 6147 8421
rect 6089 8412 6101 8415
rect 6052 8384 6101 8412
rect 6052 8372 6058 8384
rect 6089 8381 6101 8384
rect 6135 8381 6147 8415
rect 6089 8375 6147 8381
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8412 6239 8415
rect 6362 8412 6368 8424
rect 6227 8384 6368 8412
rect 6227 8381 6239 8384
rect 6181 8375 6239 8381
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 7098 8421 7104 8424
rect 7092 8412 7104 8421
rect 7059 8384 7104 8412
rect 7092 8375 7104 8384
rect 7098 8372 7104 8375
rect 7156 8372 7162 8424
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5810 8344 5816 8356
rect 5399 8316 5816 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 5184 8248 6561 8276
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6549 8239 6607 8245
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 8220 8285 8248 8452
rect 8941 8449 8953 8452
rect 8987 8480 8999 8483
rect 9122 8480 9128 8492
rect 8987 8452 9128 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 11790 8480 11796 8492
rect 9272 8452 9904 8480
rect 9272 8440 9278 8452
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8412 8815 8415
rect 9398 8412 9404 8424
rect 8803 8384 9404 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 9398 8372 9404 8384
rect 9456 8412 9462 8424
rect 9766 8412 9772 8424
rect 9456 8384 9628 8412
rect 9727 8384 9772 8412
rect 9456 8372 9462 8384
rect 9600 8288 9628 8384
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9876 8412 9904 8452
rect 11440 8452 11796 8480
rect 11440 8412 11468 8452
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 12066 8480 12072 8492
rect 12027 8452 12072 8480
rect 12066 8440 12072 8452
rect 12124 8480 12130 8492
rect 13004 8489 13032 8520
rect 12989 8483 13047 8489
rect 12124 8452 12940 8480
rect 12124 8440 12130 8452
rect 9876 8384 11468 8412
rect 11514 8372 11520 8424
rect 11572 8412 11578 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 11572 8384 11897 8412
rect 11572 8372 11578 8384
rect 11885 8381 11897 8384
rect 11931 8412 11943 8415
rect 12342 8412 12348 8424
rect 11931 8384 12348 8412
rect 11931 8381 11943 8384
rect 11885 8375 11943 8381
rect 12342 8372 12348 8384
rect 12400 8412 12406 8424
rect 12621 8415 12679 8421
rect 12621 8412 12633 8415
rect 12400 8384 12633 8412
rect 12400 8372 12406 8384
rect 12621 8381 12633 8384
rect 12667 8381 12679 8415
rect 12912 8412 12940 8452
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13078 8412 13084 8424
rect 12912 8384 13084 8412
rect 12621 8375 12679 8381
rect 13078 8372 13084 8384
rect 13136 8412 13142 8424
rect 13245 8415 13303 8421
rect 13245 8412 13257 8415
rect 13136 8384 13257 8412
rect 13136 8372 13142 8384
rect 13245 8381 13257 8384
rect 13291 8381 13303 8415
rect 13245 8375 13303 8381
rect 10036 8347 10094 8353
rect 10036 8313 10048 8347
rect 10082 8344 10094 8347
rect 10686 8344 10692 8356
rect 10082 8316 10692 8344
rect 10082 8313 10094 8316
rect 10036 8307 10094 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 11790 8304 11796 8356
rect 11848 8344 11854 8356
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 11848 8316 11989 8344
rect 11848 8304 11854 8316
rect 11977 8313 11989 8316
rect 12023 8344 12035 8347
rect 12437 8347 12495 8353
rect 12437 8344 12449 8347
rect 12023 8316 12449 8344
rect 12023 8313 12035 8316
rect 11977 8307 12035 8313
rect 12437 8313 12449 8316
rect 12483 8313 12495 8347
rect 12437 8307 12495 8313
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7524 8248 8217 8276
rect 7524 8236 7530 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8386 8276 8392 8288
rect 8347 8248 8392 8276
rect 8205 8239 8263 8245
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 8754 8276 8760 8288
rect 8536 8248 8760 8276
rect 8536 8236 8542 8248
rect 8754 8236 8760 8248
rect 8812 8276 8818 8288
rect 8849 8279 8907 8285
rect 8849 8276 8861 8279
rect 8812 8248 8861 8276
rect 8812 8236 8818 8248
rect 8849 8245 8861 8248
rect 8895 8245 8907 8279
rect 9214 8276 9220 8288
rect 9175 8248 9220 8276
rect 8849 8239 8907 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 9582 8276 9588 8288
rect 9543 8248 9588 8276
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10870 8276 10876 8288
rect 9916 8248 10876 8276
rect 9916 8236 9922 8248
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 11333 8279 11391 8285
rect 11333 8245 11345 8279
rect 11379 8276 11391 8279
rect 12250 8276 12256 8288
rect 11379 8248 12256 8276
rect 11379 8245 11391 8248
rect 11333 8239 11391 8245
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 1104 8186 16008 8208
rect 1104 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 10976 8186
rect 11028 8134 11040 8186
rect 11092 8134 11104 8186
rect 11156 8134 11168 8186
rect 11220 8134 16008 8186
rect 1104 8112 16008 8134
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 3234 8072 3240 8084
rect 2731 8044 3240 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 3651 8044 4813 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 5169 8075 5227 8081
rect 5169 8041 5181 8075
rect 5215 8072 5227 8075
rect 5629 8075 5687 8081
rect 5629 8072 5641 8075
rect 5215 8044 5641 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 5629 8041 5641 8044
rect 5675 8041 5687 8075
rect 5629 8035 5687 8041
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6420 8044 6653 8072
rect 6420 8032 6426 8044
rect 6641 8041 6653 8044
rect 6687 8072 6699 8075
rect 7098 8072 7104 8084
rect 6687 8044 7104 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7374 8072 7380 8084
rect 7331 8044 7380 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8386 8072 8392 8084
rect 8159 8044 8392 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8846 8072 8852 8084
rect 8619 8044 8852 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9214 8072 9220 8084
rect 8987 8044 9220 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 9490 8032 9496 8084
rect 9548 8032 9554 8084
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 9824 8044 9869 8072
rect 9824 8032 9830 8044
rect 9950 8032 9956 8084
rect 10008 8032 10014 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 10091 8044 11345 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 11333 8041 11345 8044
rect 11379 8041 11391 8075
rect 11333 8035 11391 8041
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12802 8072 12808 8084
rect 12575 8044 12808 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 3513 8007 3571 8013
rect 3513 7973 3525 8007
rect 3559 8004 3571 8007
rect 4890 8004 4896 8016
rect 3559 7976 4896 8004
rect 3559 7973 3571 7976
rect 3513 7967 3571 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 5258 8004 5264 8016
rect 5219 7976 5264 8004
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 5997 8007 6055 8013
rect 5997 7973 6009 8007
rect 6043 8004 6055 8007
rect 6914 8004 6920 8016
rect 6043 7976 6920 8004
rect 6043 7973 6055 7976
rect 5997 7967 6055 7973
rect 1489 7939 1547 7945
rect 1489 7905 1501 7939
rect 1535 7905 1547 7939
rect 1489 7899 1547 7905
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7936 4767 7939
rect 5442 7936 5448 7948
rect 4755 7908 5448 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 1504 7800 1532 7899
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 6012 7936 6040 7967
rect 6914 7964 6920 7976
rect 6972 8004 6978 8016
rect 6972 7976 9444 8004
rect 6972 7964 6978 7976
rect 7190 7936 7196 7948
rect 5684 7908 6040 7936
rect 7151 7908 7196 7936
rect 5684 7896 5690 7908
rect 7190 7896 7196 7908
rect 7248 7896 7254 7948
rect 7392 7908 8616 7936
rect 7392 7880 7420 7908
rect 1670 7868 1676 7880
rect 1631 7840 1676 7868
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3786 7868 3792 7880
rect 3007 7840 3648 7868
rect 3747 7840 3792 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 2317 7803 2375 7809
rect 2317 7800 2329 7803
rect 1504 7772 2329 7800
rect 2317 7769 2329 7772
rect 2363 7769 2375 7803
rect 2792 7800 2820 7831
rect 3145 7803 3203 7809
rect 3145 7800 3157 7803
rect 2792 7772 3157 7800
rect 2317 7763 2375 7769
rect 3145 7769 3157 7772
rect 3191 7769 3203 7803
rect 3620 7800 3648 7840
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 4614 7828 4620 7880
rect 4672 7868 4678 7880
rect 5353 7871 5411 7877
rect 5353 7868 5365 7871
rect 4672 7840 5365 7868
rect 4672 7828 4678 7840
rect 5353 7837 5365 7840
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 5718 7800 5724 7812
rect 3620 7772 5724 7800
rect 3145 7763 3203 7769
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 4522 7732 4528 7744
rect 4483 7704 4528 7732
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 6104 7732 6132 7831
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 7374 7868 7380 7880
rect 6236 7840 6281 7868
rect 7335 7840 7380 7868
rect 6236 7828 6242 7840
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 6825 7803 6883 7809
rect 6825 7769 6837 7803
rect 6871 7800 6883 7803
rect 8220 7800 8248 7831
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8352 7840 8397 7868
rect 8352 7828 8358 7840
rect 6871 7772 8248 7800
rect 8588 7800 8616 7908
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8720 7840 9045 7868
rect 8720 7828 8726 7840
rect 9033 7837 9045 7840
rect 9079 7837 9091 7871
rect 9033 7831 9091 7837
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9416 7868 9444 7976
rect 9508 7948 9536 8032
rect 9490 7896 9496 7948
rect 9548 7896 9554 7948
rect 9968 7945 9996 8032
rect 12250 8004 12256 8016
rect 12163 7976 12256 8004
rect 12250 7964 12256 7976
rect 12308 8004 12314 8016
rect 12308 7976 12848 8004
rect 12308 7964 12314 7976
rect 12820 7948 12848 7976
rect 9961 7939 10019 7945
rect 9961 7905 9973 7939
rect 10007 7905 10019 7939
rect 10410 7936 10416 7948
rect 10371 7908 10416 7936
rect 9961 7899 10019 7905
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 11238 7936 11244 7948
rect 11199 7908 11244 7936
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11698 7936 11704 7948
rect 11659 7908 11704 7936
rect 11698 7896 11704 7908
rect 11756 7936 11762 7948
rect 12618 7936 12624 7948
rect 11756 7908 12624 7936
rect 11756 7896 11762 7908
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12802 7896 12808 7948
rect 12860 7936 12866 7948
rect 12897 7939 12955 7945
rect 12897 7936 12909 7939
rect 12860 7908 12909 7936
rect 12860 7896 12866 7908
rect 12897 7905 12909 7908
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 10134 7868 10140 7880
rect 9416 7840 10140 7868
rect 9125 7831 9183 7837
rect 9140 7800 9168 7831
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10502 7868 10508 7880
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10686 7868 10692 7880
rect 10647 7840 10692 7868
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 11422 7868 11428 7880
rect 11383 7840 11428 7868
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12360 7840 13001 7868
rect 9306 7800 9312 7812
rect 8588 7772 9168 7800
rect 9232 7772 9312 7800
rect 6871 7769 6883 7772
rect 6825 7763 6883 7769
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 6104 7704 6561 7732
rect 6549 7701 6561 7704
rect 6595 7732 6607 7735
rect 7558 7732 7564 7744
rect 6595 7704 7564 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7745 7735 7803 7741
rect 7745 7701 7757 7735
rect 7791 7732 7803 7735
rect 9232 7732 9260 7772
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 10870 7800 10876 7812
rect 10831 7772 10876 7800
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 7791 7704 9260 7732
rect 9493 7735 9551 7741
rect 7791 7701 7803 7704
rect 7745 7695 7803 7701
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9582 7732 9588 7744
rect 9539 7704 9588 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9582 7692 9588 7704
rect 9640 7732 9646 7744
rect 12360 7741 12388 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 13136 7840 13181 7868
rect 13136 7828 13142 7840
rect 12345 7735 12403 7741
rect 12345 7732 12357 7735
rect 9640 7704 12357 7732
rect 9640 7692 9646 7704
rect 12345 7701 12357 7704
rect 12391 7701 12403 7735
rect 12345 7695 12403 7701
rect 1104 7642 16008 7664
rect 1104 7590 3480 7642
rect 3532 7590 3544 7642
rect 3596 7590 3608 7642
rect 3660 7590 3672 7642
rect 3724 7590 8478 7642
rect 8530 7590 8542 7642
rect 8594 7590 8606 7642
rect 8658 7590 8670 7642
rect 8722 7590 13475 7642
rect 13527 7590 13539 7642
rect 13591 7590 13603 7642
rect 13655 7590 13667 7642
rect 13719 7590 16008 7642
rect 1104 7568 16008 7590
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4672 7500 4813 7528
rect 4672 7488 4678 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 4801 7491 4859 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 5316 7500 5641 7528
rect 5316 7488 5322 7500
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 5629 7491 5687 7497
rect 6012 7500 6561 7528
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 1995 7296 3433 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 3421 7293 3433 7296
rect 3467 7324 3479 7327
rect 4522 7324 4528 7336
rect 3467 7296 4528 7324
rect 3467 7293 3479 7296
rect 3421 7287 3479 7293
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 6012 7324 6040 7500
rect 6549 7497 6561 7500
rect 6595 7528 6607 7531
rect 8938 7528 8944 7540
rect 6595 7500 8616 7528
rect 8899 7500 8944 7528
rect 6595 7497 6607 7500
rect 6549 7491 6607 7497
rect 8588 7472 8616 7500
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9858 7488 9864 7540
rect 9916 7528 9922 7540
rect 10318 7528 10324 7540
rect 9916 7500 10324 7528
rect 9916 7488 9922 7500
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 10502 7488 10508 7540
rect 10560 7528 10566 7540
rect 10597 7531 10655 7537
rect 10597 7528 10609 7531
rect 10560 7500 10609 7528
rect 10560 7488 10566 7500
rect 10597 7497 10609 7500
rect 10643 7497 10655 7531
rect 10597 7491 10655 7497
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11425 7531 11483 7537
rect 11425 7528 11437 7531
rect 11296 7500 11437 7528
rect 11296 7488 11302 7500
rect 11425 7497 11437 7500
rect 11471 7497 11483 7531
rect 11425 7491 11483 7497
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 7009 7463 7067 7469
rect 7009 7460 7021 7463
rect 6972 7432 7021 7460
rect 6972 7420 6978 7432
rect 7009 7429 7021 7432
rect 7055 7429 7067 7463
rect 7466 7460 7472 7472
rect 7009 7423 7067 7429
rect 7392 7432 7472 7460
rect 6178 7392 6184 7404
rect 6091 7364 6184 7392
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 6012 7296 6101 7324
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 2194 7259 2252 7265
rect 2194 7256 2206 7259
rect 2096 7228 2206 7256
rect 2096 7216 2102 7228
rect 2194 7225 2206 7228
rect 2240 7225 2252 7259
rect 3666 7259 3724 7265
rect 3666 7256 3678 7259
rect 2194 7219 2252 7225
rect 3344 7228 3678 7256
rect 3344 7197 3372 7228
rect 3666 7225 3678 7228
rect 3712 7256 3724 7259
rect 6196 7256 6224 7352
rect 7392 7333 7420 7432
rect 7466 7420 7472 7432
rect 7524 7420 7530 7472
rect 8570 7420 8576 7472
rect 8628 7420 8634 7472
rect 8849 7463 8907 7469
rect 8849 7429 8861 7463
rect 8895 7429 8907 7463
rect 8849 7423 8907 7429
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 7736 7327 7794 7333
rect 7524 7296 7569 7324
rect 7524 7284 7530 7296
rect 7736 7293 7748 7327
rect 7782 7324 7794 7327
rect 8294 7324 8300 7336
rect 7782 7296 8300 7324
rect 7782 7293 7794 7296
rect 7736 7287 7794 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 8864 7324 8892 7423
rect 9122 7420 9128 7472
rect 9180 7460 9186 7472
rect 9180 7432 9628 7460
rect 9180 7420 9186 7432
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9364 7364 9413 7392
rect 9364 7352 9370 7364
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 9508 7324 9536 7355
rect 8720 7296 9536 7324
rect 9600 7324 9628 7432
rect 10686 7420 10692 7472
rect 10744 7460 10750 7472
rect 10744 7432 12112 7460
rect 10744 7420 10750 7432
rect 12084 7404 12112 7432
rect 10318 7392 10324 7404
rect 10279 7364 10324 7392
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 10870 7352 10876 7404
rect 10928 7392 10934 7404
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10928 7364 11161 7392
rect 10928 7352 10934 7364
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 12066 7392 12072 7404
rect 12027 7364 12072 7392
rect 11149 7355 11207 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12768 7364 12909 7392
rect 12768 7352 12774 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 10226 7324 10232 7336
rect 9600 7296 10232 7324
rect 8720 7284 8726 7296
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 12912 7324 12940 7355
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13044 7364 13089 7392
rect 13044 7352 13050 7364
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 12912 7296 13461 7324
rect 13449 7293 13461 7296
rect 13495 7324 13507 7327
rect 13906 7324 13912 7336
rect 13495 7296 13912 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 6546 7256 6552 7268
rect 3712 7228 6552 7256
rect 3712 7225 3724 7228
rect 3666 7219 3724 7225
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 8754 7256 8760 7268
rect 6840 7228 8760 7256
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7157 3387 7191
rect 3329 7151 3387 7157
rect 5997 7191 6055 7197
rect 5997 7157 6009 7191
rect 6043 7188 6055 7191
rect 6270 7188 6276 7200
rect 6043 7160 6276 7188
rect 6043 7157 6055 7160
rect 5997 7151 6055 7157
rect 6270 7148 6276 7160
rect 6328 7188 6334 7200
rect 6840 7197 6868 7228
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 9030 7216 9036 7268
rect 9088 7256 9094 7268
rect 9309 7259 9367 7265
rect 9309 7256 9321 7259
rect 9088 7228 9321 7256
rect 9088 7216 9094 7228
rect 9309 7225 9321 7228
rect 9355 7225 9367 7259
rect 11057 7259 11115 7265
rect 11057 7256 11069 7259
rect 9309 7219 9367 7225
rect 9784 7228 11069 7256
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6328 7160 6837 7188
rect 6328 7148 6334 7160
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 6825 7151 6883 7157
rect 7193 7191 7251 7197
rect 7193 7157 7205 7191
rect 7239 7188 7251 7191
rect 7282 7188 7288 7200
rect 7239 7160 7288 7188
rect 7239 7157 7251 7160
rect 7193 7151 7251 7157
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 9674 7188 9680 7200
rect 7708 7160 9680 7188
rect 7708 7148 7714 7160
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9784 7197 9812 7228
rect 11057 7225 11069 7228
rect 11103 7225 11115 7259
rect 11057 7219 11115 7225
rect 11793 7259 11851 7265
rect 11793 7225 11805 7259
rect 11839 7256 11851 7259
rect 12618 7256 12624 7268
rect 11839 7228 12624 7256
rect 11839 7225 11851 7228
rect 11793 7219 11851 7225
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7157 9827 7191
rect 9769 7151 9827 7157
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10137 7191 10195 7197
rect 10137 7188 10149 7191
rect 9916 7160 10149 7188
rect 9916 7148 9922 7160
rect 10137 7157 10149 7160
rect 10183 7157 10195 7191
rect 10137 7151 10195 7157
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 10744 7160 10977 7188
rect 10744 7148 10750 7160
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 10965 7151 11023 7157
rect 11885 7191 11943 7197
rect 11885 7157 11897 7191
rect 11931 7188 11943 7191
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 11931 7160 12449 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12437 7151 12495 7157
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 13078 7188 13084 7200
rect 12851 7160 13084 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13078 7148 13084 7160
rect 13136 7188 13142 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 13136 7160 13277 7188
rect 13136 7148 13142 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 1104 7098 16008 7120
rect 1104 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 10976 7098
rect 11028 7046 11040 7098
rect 11092 7046 11104 7098
rect 11156 7046 11168 7098
rect 11220 7046 16008 7098
rect 1104 7024 16008 7046
rect 1857 6987 1915 6993
rect 1857 6953 1869 6987
rect 1903 6984 1915 6987
rect 2225 6987 2283 6993
rect 2225 6984 2237 6987
rect 1903 6956 2237 6984
rect 1903 6953 1915 6956
rect 1857 6947 1915 6953
rect 2225 6953 2237 6956
rect 2271 6953 2283 6987
rect 2225 6947 2283 6953
rect 4341 6987 4399 6993
rect 4341 6953 4353 6987
rect 4387 6953 4399 6987
rect 4341 6947 4399 6953
rect 4709 6987 4767 6993
rect 4709 6953 4721 6987
rect 4755 6984 4767 6987
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4755 6956 5181 6984
rect 4755 6953 4767 6956
rect 4709 6947 4767 6953
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 7650 6984 7656 6996
rect 5169 6947 5227 6953
rect 6656 6956 7656 6984
rect 1765 6919 1823 6925
rect 1765 6885 1777 6919
rect 1811 6916 1823 6919
rect 4356 6916 4384 6947
rect 6656 6928 6684 6956
rect 7650 6944 7656 6956
rect 7708 6944 7714 6996
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 10686 6984 10692 6996
rect 8404 6956 10692 6984
rect 1811 6888 4384 6916
rect 6365 6919 6423 6925
rect 1811 6885 1823 6888
rect 1765 6879 1823 6885
rect 6365 6885 6377 6919
rect 6411 6916 6423 6919
rect 6638 6916 6644 6928
rect 6411 6888 6644 6916
rect 6411 6885 6423 6888
rect 6365 6879 6423 6885
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 7184 6919 7242 6925
rect 7184 6885 7196 6919
rect 7230 6916 7242 6919
rect 7374 6916 7380 6928
rect 7230 6888 7380 6916
rect 7230 6885 7242 6888
rect 7184 6879 7242 6885
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 8404 6916 8432 6956
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 10870 6944 10876 6996
rect 10928 6984 10934 6996
rect 11057 6987 11115 6993
rect 11057 6984 11069 6987
rect 10928 6956 11069 6984
rect 10928 6944 10934 6956
rect 11057 6953 11069 6956
rect 11103 6953 11115 6987
rect 11057 6947 11115 6953
rect 7616 6888 8432 6916
rect 7616 6876 7622 6888
rect 8662 6876 8668 6928
rect 8720 6916 8726 6928
rect 8846 6916 8852 6928
rect 8720 6888 8852 6916
rect 8720 6876 8726 6888
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 9122 6876 9128 6928
rect 9180 6916 9186 6928
rect 9582 6916 9588 6928
rect 9180 6888 9588 6916
rect 9180 6876 9186 6888
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 9944 6919 10002 6925
rect 9944 6916 9956 6919
rect 9732 6888 9956 6916
rect 9732 6876 9738 6888
rect 9944 6885 9956 6888
rect 9990 6916 10002 6919
rect 10318 6916 10324 6928
rect 9990 6888 10324 6916
rect 9990 6885 10002 6888
rect 9944 6879 10002 6885
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 2590 6848 2596 6860
rect 2551 6820 2596 6848
rect 2590 6808 2596 6820
rect 2648 6808 2654 6860
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 2866 6848 2872 6860
rect 2731 6820 2872 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 5534 6848 5540 6860
rect 5495 6820 5540 6848
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6086 6848 6092 6860
rect 5675 6820 6092 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6848 6515 6851
rect 6730 6848 6736 6860
rect 6503 6820 6736 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7466 6848 7472 6860
rect 6963 6820 7472 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 7466 6808 7472 6820
rect 7524 6848 7530 6860
rect 9766 6848 9772 6860
rect 7524 6820 9772 6848
rect 7524 6808 7530 6820
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2608 6752 2789 6780
rect 1670 6672 1676 6724
rect 1728 6712 1734 6724
rect 2498 6712 2504 6724
rect 1728 6684 2504 6712
rect 1728 6672 1734 6684
rect 2498 6672 2504 6684
rect 2556 6712 2562 6724
rect 2608 6712 2636 6752
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 4798 6780 4804 6792
rect 4759 6752 4804 6780
rect 2777 6743 2835 6749
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 4893 6783 4951 6789
rect 4893 6749 4905 6783
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 2556 6684 2636 6712
rect 2556 6672 2562 6684
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 4908 6712 4936 6743
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 5776 6752 5821 6780
rect 5776 6740 5782 6752
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 6604 6752 6649 6780
rect 6604 6740 6610 6752
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9692 6789 9720 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9272 6752 9413 6780
rect 9272 6740 9278 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9401 6743 9459 6749
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 10704 6780 10732 6944
rect 11072 6848 11100 6947
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12676 6956 12909 6984
rect 12676 6944 12682 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 11692 6851 11750 6857
rect 11692 6848 11704 6851
rect 11072 6820 11704 6848
rect 11692 6817 11704 6820
rect 11738 6848 11750 6851
rect 13262 6848 13268 6860
rect 11738 6820 13032 6848
rect 13223 6820 13268 6848
rect 11738 6817 11750 6820
rect 11692 6811 11750 6817
rect 13004 6792 13032 6820
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13412 6820 13737 6848
rect 13412 6808 13418 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 9723 6752 9757 6780
rect 10704 6752 11284 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 4672 6684 4936 6712
rect 4672 6672 4678 6684
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 5868 6684 6009 6712
rect 5868 6672 5874 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 8570 6672 8576 6724
rect 8628 6672 8634 6724
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9309 6715 9367 6721
rect 9309 6712 9321 6715
rect 8812 6684 9321 6712
rect 8812 6672 8818 6684
rect 9309 6681 9321 6684
rect 9355 6712 9367 6715
rect 9355 6684 9720 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 1397 6647 1455 6653
rect 1397 6613 1409 6647
rect 1443 6644 1455 6647
rect 1486 6644 1492 6656
rect 1443 6616 1492 6644
rect 1443 6613 1455 6616
rect 1397 6607 1455 6613
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 8588 6644 8616 6672
rect 9214 6644 9220 6656
rect 8588 6616 9220 6644
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9692 6644 9720 6684
rect 9858 6644 9864 6656
rect 9692 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 11256 6653 11284 6752
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 11388 6752 11437 6780
rect 11388 6740 11394 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13044 6752 13553 6780
rect 13044 6740 13050 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 11241 6647 11299 6653
rect 11241 6613 11253 6647
rect 11287 6644 11299 6647
rect 11330 6644 11336 6656
rect 11287 6616 11336 6644
rect 11287 6613 11299 6616
rect 11241 6607 11299 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 12805 6647 12863 6653
rect 12805 6644 12817 6647
rect 12124 6616 12817 6644
rect 12124 6604 12130 6616
rect 12805 6613 12817 6616
rect 12851 6613 12863 6647
rect 12805 6607 12863 6613
rect 1104 6554 16008 6576
rect 1104 6502 3480 6554
rect 3532 6502 3544 6554
rect 3596 6502 3608 6554
rect 3660 6502 3672 6554
rect 3724 6502 8478 6554
rect 8530 6502 8542 6554
rect 8594 6502 8606 6554
rect 8658 6502 8670 6554
rect 8722 6502 13475 6554
rect 13527 6502 13539 6554
rect 13591 6502 13603 6554
rect 13655 6502 13667 6554
rect 13719 6502 16008 6554
rect 1104 6480 16008 6502
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2096 6412 2789 6440
rect 2096 6400 2102 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 4614 6440 4620 6452
rect 2777 6403 2835 6409
rect 3252 6412 4620 6440
rect 2498 6332 2504 6384
rect 2556 6372 2562 6384
rect 3252 6372 3280 6412
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 5169 6443 5227 6449
rect 5169 6440 5181 6443
rect 4856 6412 5181 6440
rect 4856 6400 4862 6412
rect 5169 6409 5181 6412
rect 5215 6409 5227 6443
rect 5169 6403 5227 6409
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5500 6412 6009 6440
rect 5500 6400 5506 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 5997 6403 6055 6409
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6144 6412 6561 6440
rect 6144 6400 6150 6412
rect 6549 6409 6561 6412
rect 6595 6440 6607 6443
rect 7006 6440 7012 6452
rect 6595 6412 7012 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 7006 6400 7012 6412
rect 7064 6440 7070 6452
rect 8018 6440 8024 6452
rect 7064 6412 8024 6440
rect 7064 6400 7070 6412
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 9674 6440 9680 6452
rect 8312 6412 9536 6440
rect 9635 6412 9680 6440
rect 2556 6344 3280 6372
rect 2556 6332 2562 6344
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 6825 6375 6883 6381
rect 6825 6372 6837 6375
rect 6788 6344 6837 6372
rect 6788 6332 6794 6344
rect 6825 6341 6837 6344
rect 6871 6372 6883 6375
rect 8312 6372 8340 6412
rect 6871 6344 8340 6372
rect 9508 6372 9536 6412
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 9950 6440 9956 6452
rect 9815 6412 9956 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10229 6443 10287 6449
rect 10229 6440 10241 6443
rect 10192 6412 10241 6440
rect 10192 6400 10198 6412
rect 10229 6409 10241 6412
rect 10275 6409 10287 6443
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 10229 6403 10287 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 10594 6372 10600 6384
rect 9508 6344 10600 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 5718 6304 5724 6316
rect 1443 6276 1532 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1394 6128 1400 6180
rect 1452 6168 1458 6180
rect 1504 6168 1532 6276
rect 4448 6276 5724 6304
rect 1670 6245 1676 6248
rect 1653 6239 1676 6245
rect 1653 6205 1665 6239
rect 1653 6199 1676 6205
rect 1670 6196 1676 6199
rect 1728 6196 1734 6248
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 4246 6236 4252 6248
rect 3283 6208 4252 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 3252 6168 3280 6199
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 1452 6140 3280 6168
rect 1452 6128 1458 6140
rect 3418 6128 3424 6180
rect 3476 6177 3482 6180
rect 3476 6171 3540 6177
rect 3476 6137 3494 6171
rect 3528 6168 3540 6171
rect 4448 6168 4476 6276
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6273 6307 6331 6313
rect 6273 6304 6285 6307
rect 6104 6276 6285 6304
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 5408 6208 5549 6236
rect 5408 6196 5414 6208
rect 5537 6205 5549 6208
rect 5583 6236 5595 6239
rect 6104 6236 6132 6276
rect 6273 6273 6285 6276
rect 6319 6304 6331 6307
rect 7190 6304 7196 6316
rect 6319 6276 7196 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 10870 6264 10876 6316
rect 10928 6304 10934 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10928 6276 10977 6304
rect 10928 6264 10934 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 13262 6304 13268 6316
rect 12115 6276 13268 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 5583 6208 6132 6236
rect 6181 6239 6239 6245
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 6181 6205 6193 6239
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 3528 6140 4476 6168
rect 6196 6168 6224 6199
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 6880 6208 7941 6236
rect 6880 6196 6886 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 7929 6199 7987 6205
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 8168 6208 8309 6236
rect 8168 6196 8174 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8564 6239 8622 6245
rect 8564 6205 8576 6239
rect 8610 6236 8622 6239
rect 8846 6236 8852 6248
rect 8610 6208 8852 6236
rect 8610 6205 8622 6208
rect 8564 6199 8622 6205
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 7282 6168 7288 6180
rect 6196 6140 7288 6168
rect 3528 6137 3540 6140
rect 3476 6131 3540 6137
rect 3476 6128 3482 6131
rect 7282 6128 7288 6140
rect 7340 6168 7346 6180
rect 9968 6168 9996 6199
rect 7340 6140 9996 6168
rect 10781 6171 10839 6177
rect 7340 6128 7346 6140
rect 10781 6137 10793 6171
rect 10827 6168 10839 6171
rect 10827 6140 11376 6168
rect 10827 6137 10839 6140
rect 10781 6131 10839 6137
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 6638 6100 6644 6112
rect 5675 6072 6644 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7009 6103 7067 6109
rect 7009 6100 7021 6103
rect 6788 6072 7021 6100
rect 6788 6060 6794 6072
rect 7009 6069 7021 6072
rect 7055 6069 7067 6103
rect 7009 6063 7067 6069
rect 7193 6103 7251 6109
rect 7193 6069 7205 6103
rect 7239 6100 7251 6103
rect 7374 6100 7380 6112
rect 7239 6072 7380 6100
rect 7239 6069 7251 6072
rect 7193 6063 7251 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10042 6100 10048 6112
rect 9732 6072 10048 6100
rect 9732 6060 9738 6072
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10686 6100 10692 6112
rect 10192 6072 10692 6100
rect 10192 6060 10198 6072
rect 10686 6060 10692 6072
rect 10744 6100 10750 6112
rect 11348 6109 11376 6140
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10744 6072 10885 6100
rect 10744 6060 10750 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 11333 6103 11391 6109
rect 11333 6069 11345 6103
rect 11379 6100 11391 6103
rect 11882 6100 11888 6112
rect 11379 6072 11888 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 1104 6010 16008 6032
rect 1104 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 10976 6010
rect 11028 5958 11040 6010
rect 11092 5958 11104 6010
rect 11156 5958 11168 6010
rect 11220 5958 16008 6010
rect 1104 5936 16008 5958
rect 2041 5899 2099 5905
rect 2041 5865 2053 5899
rect 2087 5896 2099 5899
rect 2590 5896 2596 5908
rect 2087 5868 2596 5896
rect 2087 5865 2099 5868
rect 2041 5859 2099 5865
rect 2590 5856 2596 5868
rect 2648 5856 2654 5908
rect 2866 5896 2872 5908
rect 2827 5868 2872 5896
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 4154 5896 4160 5908
rect 3835 5868 4160 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 1762 5828 1768 5840
rect 1723 5800 1768 5828
rect 1762 5788 1768 5800
rect 1820 5788 1826 5840
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5828 2467 5831
rect 3804 5828 3832 5859
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 5592 5868 5641 5896
rect 5592 5856 5598 5868
rect 5629 5865 5641 5868
rect 5675 5865 5687 5899
rect 5629 5859 5687 5865
rect 6365 5899 6423 5905
rect 6365 5865 6377 5899
rect 6411 5896 6423 5899
rect 7006 5896 7012 5908
rect 6411 5868 7012 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 11514 5896 11520 5908
rect 7432 5868 11520 5896
rect 7432 5856 7438 5868
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 2455 5800 3832 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 4062 5788 4068 5840
rect 4120 5788 4126 5840
rect 4246 5828 4252 5840
rect 4159 5800 4252 5828
rect 1486 5760 1492 5772
rect 1447 5732 1492 5760
rect 1486 5720 1492 5732
rect 1544 5720 1550 5772
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 4080 5760 4108 5788
rect 3283 5732 4108 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 2498 5692 2504 5704
rect 2459 5664 2504 5692
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 3326 5692 3332 5704
rect 3287 5664 3332 5692
rect 2685 5655 2743 5661
rect 2700 5624 2728 5655
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 4065 5695 4123 5701
rect 3476 5664 3569 5692
rect 3476 5652 3482 5664
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4172 5692 4200 5800
rect 4246 5788 4252 5800
rect 4304 5828 4310 5840
rect 5258 5828 5264 5840
rect 4304 5800 5264 5828
rect 4304 5788 4310 5800
rect 5258 5788 5264 5800
rect 5316 5788 5322 5840
rect 6638 5788 6644 5840
rect 6696 5828 6702 5840
rect 7392 5828 7420 5856
rect 6696 5800 7420 5828
rect 6696 5788 6702 5800
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 8757 5831 8815 5837
rect 8757 5828 8769 5831
rect 7892 5800 8769 5828
rect 7892 5788 7898 5800
rect 8757 5797 8769 5800
rect 8803 5828 8815 5831
rect 9030 5828 9036 5840
rect 8803 5800 9036 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 9030 5788 9036 5800
rect 9088 5828 9094 5840
rect 9493 5831 9551 5837
rect 9493 5828 9505 5831
rect 9088 5800 9505 5828
rect 9088 5788 9094 5800
rect 9493 5797 9505 5800
rect 9539 5797 9551 5831
rect 9493 5791 9551 5797
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 9858 5828 9864 5840
rect 9732 5800 9777 5828
rect 9819 5800 9864 5828
rect 9732 5788 9738 5800
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 10686 5828 10692 5840
rect 10647 5800 10692 5828
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 14918 5828 14924 5840
rect 14879 5800 14924 5828
rect 14918 5788 14924 5800
rect 14976 5788 14982 5840
rect 4338 5769 4344 5772
rect 4332 5760 4344 5769
rect 4299 5732 4344 5760
rect 4332 5723 4344 5732
rect 4338 5720 4344 5723
rect 4396 5720 4402 5772
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6914 5760 6920 5772
rect 6503 5732 6920 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7092 5763 7150 5769
rect 7092 5729 7104 5763
rect 7138 5760 7150 5763
rect 7466 5760 7472 5772
rect 7138 5732 7472 5760
rect 7138 5729 7150 5732
rect 7092 5723 7150 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 8665 5763 8723 5769
rect 8665 5760 8677 5763
rect 8352 5732 8677 5760
rect 8352 5720 8358 5732
rect 8665 5729 8677 5732
rect 8711 5760 8723 5763
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 8711 5732 9229 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 9217 5729 9229 5732
rect 9263 5760 9275 5763
rect 9263 5732 9720 5760
rect 9263 5729 9275 5732
rect 9217 5723 9275 5729
rect 4111 5664 4200 5692
rect 6641 5695 6699 5701
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 6641 5661 6653 5695
rect 6687 5692 6699 5695
rect 6730 5692 6736 5704
rect 6687 5664 6736 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 8846 5692 8852 5704
rect 8807 5664 8852 5692
rect 6825 5655 6883 5661
rect 3436 5624 3464 5652
rect 2700 5596 4108 5624
rect 4080 5556 4108 5596
rect 5258 5584 5264 5636
rect 5316 5624 5322 5636
rect 6840 5624 6868 5655
rect 8846 5652 8852 5664
rect 8904 5692 8910 5704
rect 9582 5692 9588 5704
rect 8904 5664 9588 5692
rect 8904 5652 8910 5664
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9692 5692 9720 5732
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 10008 5732 10333 5760
rect 10008 5720 10014 5732
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 14642 5760 14648 5772
rect 14603 5732 14648 5760
rect 10321 5723 10379 5729
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 11514 5692 11520 5704
rect 9692 5664 11520 5692
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 5316 5596 6868 5624
rect 5316 5584 5322 5596
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 10137 5627 10195 5633
rect 10137 5624 10149 5627
rect 8168 5596 10149 5624
rect 8168 5584 8174 5596
rect 10137 5593 10149 5596
rect 10183 5624 10195 5627
rect 10778 5624 10784 5636
rect 10183 5596 10784 5624
rect 10183 5593 10195 5596
rect 10137 5587 10195 5593
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 5445 5559 5503 5565
rect 5445 5556 5457 5559
rect 4080 5528 5457 5556
rect 5445 5525 5457 5528
rect 5491 5525 5503 5559
rect 5445 5519 5503 5525
rect 5997 5559 6055 5565
rect 5997 5525 6009 5559
rect 6043 5556 6055 5559
rect 6362 5556 6368 5568
rect 6043 5528 6368 5556
rect 6043 5525 6055 5528
rect 5997 5519 6055 5525
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 8202 5556 8208 5568
rect 6788 5528 8208 5556
rect 6788 5516 6794 5528
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 9306 5556 9312 5568
rect 8352 5528 8397 5556
rect 9267 5528 9312 5556
rect 8352 5516 8358 5528
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 9493 5559 9551 5565
rect 9493 5525 9505 5559
rect 9539 5556 9551 5559
rect 10505 5559 10563 5565
rect 10505 5556 10517 5559
rect 9539 5528 10517 5556
rect 9539 5525 9551 5528
rect 9493 5519 9551 5525
rect 10505 5525 10517 5528
rect 10551 5556 10563 5559
rect 12710 5556 12716 5568
rect 10551 5528 12716 5556
rect 10551 5525 10563 5528
rect 10505 5519 10563 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 1104 5466 16008 5488
rect 1104 5414 3480 5466
rect 3532 5414 3544 5466
rect 3596 5414 3608 5466
rect 3660 5414 3672 5466
rect 3724 5414 8478 5466
rect 8530 5414 8542 5466
rect 8594 5414 8606 5466
rect 8658 5414 8670 5466
rect 8722 5414 13475 5466
rect 13527 5414 13539 5466
rect 13591 5414 13603 5466
rect 13655 5414 13667 5466
rect 13719 5414 16008 5466
rect 1104 5392 16008 5414
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2556 5324 2605 5352
rect 2556 5312 2562 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 3421 5355 3479 5361
rect 3421 5352 3433 5355
rect 3384 5324 3433 5352
rect 3384 5312 3390 5324
rect 3421 5321 3433 5324
rect 3467 5321 3479 5355
rect 3421 5315 3479 5321
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 4212 5324 4261 5352
rect 4212 5312 4218 5324
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 4249 5315 4307 5321
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 6914 5352 6920 5364
rect 5224 5324 6776 5352
rect 6875 5324 6920 5352
rect 5224 5312 5230 5324
rect 6748 5284 6776 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 8076 5324 8217 5352
rect 8076 5312 8082 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 9769 5355 9827 5361
rect 9769 5352 9781 5355
rect 9640 5324 9781 5352
rect 9640 5312 9646 5324
rect 9769 5321 9781 5324
rect 9815 5321 9827 5355
rect 9769 5315 9827 5321
rect 9953 5355 10011 5361
rect 9953 5321 9965 5355
rect 9999 5352 10011 5355
rect 11422 5352 11428 5364
rect 9999 5324 11428 5352
rect 9999 5321 10011 5324
rect 9953 5315 10011 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 11756 5324 15301 5352
rect 11756 5312 11762 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 7834 5284 7840 5296
rect 6748 5256 7840 5284
rect 7834 5244 7840 5256
rect 7892 5244 7898 5296
rect 8110 5244 8116 5296
rect 8168 5284 8174 5296
rect 12161 5287 12219 5293
rect 8168 5256 8432 5284
rect 8168 5244 8174 5256
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3283 5188 4077 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 4065 5185 4077 5188
rect 4111 5216 4123 5219
rect 4338 5216 4344 5228
rect 4111 5188 4344 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4338 5176 4344 5188
rect 4396 5216 4402 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4396 5188 4813 5216
rect 4396 5176 4402 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 4801 5179 4859 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 8404 5225 8432 5256
rect 12161 5253 12173 5287
rect 12207 5253 12219 5287
rect 12161 5247 12219 5253
rect 13817 5287 13875 5293
rect 13817 5253 13829 5287
rect 13863 5253 13875 5287
rect 13817 5247 13875 5253
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 10686 5216 10692 5228
rect 10643 5188 10692 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 3326 5108 3332 5160
rect 3384 5148 3390 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3384 5120 3801 5148
rect 3384 5108 3390 5120
rect 3789 5117 3801 5120
rect 3835 5148 3847 5151
rect 4982 5148 4988 5160
rect 3835 5120 4988 5148
rect 3835 5117 3847 5120
rect 3789 5111 3847 5117
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5148 5227 5151
rect 5258 5148 5264 5160
rect 5215 5120 5264 5148
rect 5215 5117 5227 5120
rect 5169 5111 5227 5117
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5436 5151 5494 5157
rect 5436 5117 5448 5151
rect 5482 5148 5494 5151
rect 6730 5148 6736 5160
rect 5482 5120 6736 5148
rect 5482 5117 5494 5120
rect 5436 5111 5494 5117
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 7285 5151 7343 5157
rect 7285 5148 7297 5151
rect 7248 5120 7297 5148
rect 7248 5108 7254 5120
rect 7285 5117 7297 5120
rect 7331 5148 7343 5151
rect 7742 5148 7748 5160
rect 7331 5120 7748 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7742 5108 7748 5120
rect 7800 5148 7806 5160
rect 8021 5151 8079 5157
rect 8021 5148 8033 5151
rect 7800 5120 8033 5148
rect 7800 5108 7806 5120
rect 8021 5117 8033 5120
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 10778 5148 10784 5160
rect 8536 5120 10640 5148
rect 10739 5120 10784 5148
rect 8536 5108 8542 5120
rect 2406 5040 2412 5092
rect 2464 5080 2470 5092
rect 3970 5080 3976 5092
rect 2464 5052 3976 5080
rect 2464 5040 2470 5052
rect 3970 5040 3976 5052
rect 4028 5080 4034 5092
rect 4617 5083 4675 5089
rect 4617 5080 4629 5083
rect 4028 5052 4629 5080
rect 4028 5040 4034 5052
rect 4617 5049 4629 5052
rect 4663 5080 4675 5083
rect 4663 5052 5028 5080
rect 4663 5049 4675 5052
rect 4617 5043 4675 5049
rect 2958 5012 2964 5024
rect 2919 4984 2964 5012
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 5012 3111 5015
rect 3602 5012 3608 5024
rect 3099 4984 3608 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 3881 5015 3939 5021
rect 3881 4981 3893 5015
rect 3927 5012 3939 5015
rect 4246 5012 4252 5024
rect 3927 4984 4252 5012
rect 3927 4981 3939 4984
rect 3881 4975 3939 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5000 5012 5028 5052
rect 5074 5040 5080 5092
rect 5132 5080 5138 5092
rect 5132 5052 6684 5080
rect 5132 5040 5138 5052
rect 5166 5012 5172 5024
rect 5000 4984 5172 5012
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 6656 5012 6684 5052
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 7377 5083 7435 5089
rect 7377 5080 7389 5083
rect 6972 5052 7389 5080
rect 6972 5040 6978 5052
rect 7377 5049 7389 5052
rect 7423 5049 7435 5083
rect 8656 5083 8714 5089
rect 7377 5043 7435 5049
rect 7484 5052 7880 5080
rect 7484 5012 7512 5052
rect 7742 5012 7748 5024
rect 6656 4984 7512 5012
rect 7703 4984 7748 5012
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 7852 5012 7880 5052
rect 8656 5049 8668 5083
rect 8702 5080 8714 5083
rect 9398 5080 9404 5092
rect 8702 5052 9404 5080
rect 8702 5049 8714 5052
rect 8656 5043 8714 5049
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 10321 5083 10379 5089
rect 10321 5049 10333 5083
rect 10367 5080 10379 5083
rect 10502 5080 10508 5092
rect 10367 5052 10508 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 10502 5040 10508 5052
rect 10560 5040 10566 5092
rect 10226 5012 10232 5024
rect 7852 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 10410 4972 10416 5024
rect 10468 5012 10474 5024
rect 10612 5012 10640 5120
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 12176 5148 12204 5247
rect 13832 5216 13860 5247
rect 13832 5188 14044 5216
rect 10888 5120 12204 5148
rect 12437 5151 12495 5157
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 10888 5080 10916 5120
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 13909 5151 13967 5157
rect 13909 5148 13921 5151
rect 12483 5120 13921 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12912 5092 12940 5120
rect 13909 5117 13921 5120
rect 13955 5117 13967 5151
rect 13909 5111 13967 5117
rect 10744 5052 10916 5080
rect 11048 5083 11106 5089
rect 10744 5040 10750 5052
rect 11048 5049 11060 5083
rect 11094 5080 11106 5083
rect 11698 5080 11704 5092
rect 11094 5052 11704 5080
rect 11094 5049 11106 5052
rect 11048 5043 11106 5049
rect 11698 5040 11704 5052
rect 11756 5040 11762 5092
rect 12618 5040 12624 5092
rect 12676 5089 12682 5092
rect 12676 5083 12740 5089
rect 12676 5049 12694 5083
rect 12728 5049 12740 5083
rect 12676 5043 12740 5049
rect 12676 5040 12682 5043
rect 12894 5040 12900 5092
rect 12952 5040 12958 5092
rect 14016 5080 14044 5188
rect 14176 5083 14234 5089
rect 14176 5080 14188 5083
rect 14016 5052 14188 5080
rect 14176 5049 14188 5052
rect 14222 5080 14234 5083
rect 14918 5080 14924 5092
rect 14222 5052 14924 5080
rect 14222 5049 14234 5052
rect 14176 5043 14234 5049
rect 14918 5040 14924 5052
rect 14976 5040 14982 5092
rect 14274 5012 14280 5024
rect 10468 4984 10513 5012
rect 10612 4984 14280 5012
rect 10468 4972 10474 4984
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 1104 4922 16008 4944
rect 1104 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 10976 4922
rect 11028 4870 11040 4922
rect 11092 4870 11104 4922
rect 11156 4870 11168 4922
rect 11220 4870 16008 4922
rect 1104 4848 16008 4870
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 1504 4780 6009 4808
rect 1504 4681 1532 4780
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 5997 4771 6055 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 6825 4811 6883 4817
rect 6825 4808 6837 4811
rect 6696 4780 6837 4808
rect 6696 4768 6702 4780
rect 6825 4777 6837 4780
rect 6871 4777 6883 4811
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 6825 4771 6883 4777
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 7742 4808 7748 4820
rect 7423 4780 7748 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 8297 4811 8355 4817
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8343 4780 8677 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8665 4777 8677 4780
rect 8711 4777 8723 4811
rect 9122 4808 9128 4820
rect 8665 4771 8723 4777
rect 8956 4780 9128 4808
rect 2314 4740 2320 4752
rect 2275 4712 2320 4740
rect 2314 4700 2320 4712
rect 2372 4700 2378 4752
rect 3602 4740 3608 4752
rect 3515 4712 3608 4740
rect 3602 4700 3608 4712
rect 3660 4740 3666 4752
rect 4890 4740 4896 4752
rect 3660 4712 4896 4740
rect 3660 4700 3666 4712
rect 4890 4700 4896 4712
rect 4948 4740 4954 4752
rect 5074 4740 5080 4752
rect 4948 4712 5080 4740
rect 4948 4700 4954 4712
rect 5074 4700 5080 4712
rect 5132 4700 5138 4752
rect 5166 4700 5172 4752
rect 5224 4740 5230 4752
rect 5261 4743 5319 4749
rect 5261 4740 5273 4743
rect 5224 4712 5273 4740
rect 5224 4700 5230 4712
rect 5261 4709 5273 4712
rect 5307 4709 5319 4743
rect 5261 4703 5319 4709
rect 5350 4700 5356 4752
rect 5408 4740 5414 4752
rect 5813 4743 5871 4749
rect 5813 4740 5825 4743
rect 5408 4712 5825 4740
rect 5408 4700 5414 4712
rect 5813 4709 5825 4712
rect 5859 4740 5871 4743
rect 6730 4740 6736 4752
rect 5859 4712 6736 4740
rect 5859 4709 5871 4712
rect 5813 4703 5871 4709
rect 6730 4700 6736 4712
rect 6788 4700 6794 4752
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 7469 4743 7527 4749
rect 7469 4740 7481 4743
rect 7340 4712 7481 4740
rect 7340 4700 7346 4712
rect 7469 4709 7481 4712
rect 7515 4740 7527 4743
rect 8018 4740 8024 4752
rect 7515 4712 8024 4740
rect 7515 4709 7527 4712
rect 7469 4703 7527 4709
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 8205 4743 8263 4749
rect 8205 4709 8217 4743
rect 8251 4740 8263 4743
rect 8956 4740 8984 4780
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10410 4808 10416 4820
rect 10183 4780 10416 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 10965 4811 11023 4817
rect 10965 4808 10977 4811
rect 10704 4780 10977 4808
rect 8251 4712 8984 4740
rect 9033 4743 9091 4749
rect 8251 4709 8263 4712
rect 8205 4703 8263 4709
rect 9033 4709 9045 4743
rect 9079 4740 9091 4743
rect 9079 4712 9628 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 2041 4675 2099 4681
rect 2041 4641 2053 4675
rect 2087 4641 2099 4675
rect 3050 4672 3056 4684
rect 3011 4644 3056 4672
rect 2041 4635 2099 4641
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 2056 4536 2084 4635
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 4614 4672 4620 4684
rect 3191 4644 4620 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 5442 4672 5448 4684
rect 4755 4644 5448 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 7650 4672 7656 4684
rect 6503 4644 7656 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 8220 4672 8248 4703
rect 8846 4672 8852 4684
rect 7800 4644 8248 4672
rect 8404 4644 8852 4672
rect 7800 4632 7806 4644
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 4246 4604 4252 4616
rect 3292 4576 3337 4604
rect 4207 4576 4252 4604
rect 3292 4564 3298 4576
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 5258 4604 5264 4616
rect 4540 4576 5264 4604
rect 2685 4539 2743 4545
rect 2685 4536 2697 4539
rect 2056 4508 2697 4536
rect 2685 4505 2697 4508
rect 2731 4505 2743 4539
rect 2685 4499 2743 4505
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3789 4539 3847 4545
rect 3789 4536 3801 4539
rect 3016 4508 3801 4536
rect 3016 4496 3022 4508
rect 3789 4505 3801 4508
rect 3835 4536 3847 4539
rect 3970 4536 3976 4548
rect 3835 4508 3976 4536
rect 3835 4505 3847 4508
rect 3789 4499 3847 4505
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 3326 4468 3332 4480
rect 1636 4440 3332 4468
rect 1636 4428 1642 4440
rect 3326 4428 3332 4440
rect 3384 4428 3390 4480
rect 4264 4468 4292 4564
rect 4540 4545 4568 4576
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6604 4576 6649 4604
rect 6604 4564 6610 4576
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 8404 4613 8432 4644
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 9600 4672 9628 4712
rect 9858 4700 9864 4752
rect 9916 4740 9922 4752
rect 10505 4743 10563 4749
rect 10505 4740 10517 4743
rect 9916 4712 10517 4740
rect 9916 4700 9922 4712
rect 10505 4709 10517 4712
rect 10551 4709 10563 4743
rect 10505 4703 10563 4709
rect 9766 4672 9772 4684
rect 9600 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10704 4672 10732 4780
rect 10965 4777 10977 4780
rect 11011 4777 11023 4811
rect 10965 4771 11023 4777
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4777 13599 4811
rect 13541 4771 13599 4777
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 14642 4808 14648 4820
rect 14415 4780 14648 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 12152 4743 12210 4749
rect 10836 4712 11928 4740
rect 10836 4700 10842 4712
rect 10520 4644 10732 4672
rect 10520 4616 10548 4644
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 11900 4681 11928 4712
rect 12152 4709 12164 4743
rect 12198 4740 12210 4743
rect 12250 4740 12256 4752
rect 12198 4712 12256 4740
rect 12198 4709 12210 4712
rect 12152 4703 12210 4709
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 13556 4740 13584 4771
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 14737 4743 14795 4749
rect 14737 4740 14749 4743
rect 13556 4712 14749 4740
rect 14737 4709 14749 4712
rect 14783 4709 14795 4743
rect 14737 4703 14795 4709
rect 11333 4675 11391 4681
rect 11333 4672 11345 4675
rect 10928 4644 11345 4672
rect 10928 4632 10934 4644
rect 11333 4641 11345 4644
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4672 11943 4675
rect 12894 4672 12900 4684
rect 11931 4644 12900 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 13909 4675 13967 4681
rect 13909 4641 13921 4675
rect 13955 4672 13967 4675
rect 14642 4672 14648 4684
rect 13955 4644 14648 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 14826 4672 14832 4684
rect 14787 4644 14832 4672
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7524 4576 7573 4604
rect 7524 4564 7530 4576
rect 7561 4573 7573 4576
rect 7607 4604 7619 4607
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 7607 4576 8401 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8938 4604 8944 4616
rect 8389 4567 8447 4573
rect 8496 4576 8944 4604
rect 4525 4539 4583 4545
rect 4525 4505 4537 4539
rect 4571 4505 4583 4539
rect 5537 4539 5595 4545
rect 4525 4499 4583 4505
rect 4816 4508 5488 4536
rect 4816 4468 4844 4508
rect 4264 4440 4844 4468
rect 4893 4471 4951 4477
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 4982 4468 4988 4480
rect 4939 4440 4988 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5166 4468 5172 4480
rect 5127 4440 5172 4468
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5460 4468 5488 4508
rect 5537 4505 5549 4539
rect 5583 4536 5595 4539
rect 5626 4536 5632 4548
rect 5583 4508 5632 4536
rect 5583 4505 5595 4508
rect 5537 4499 5595 4505
rect 5626 4496 5632 4508
rect 5684 4536 5690 4548
rect 6454 4536 6460 4548
rect 5684 4508 6460 4536
rect 5684 4496 5690 4508
rect 6454 4496 6460 4508
rect 6512 4496 6518 4548
rect 8496 4536 8524 4576
rect 7668 4508 8524 4536
rect 7668 4468 7696 4508
rect 7834 4468 7840 4480
rect 5460 4440 7696 4468
rect 7795 4440 7840 4468
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 8772 4468 8800 4576
rect 8938 4564 8944 4576
rect 8996 4604 9002 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8996 4576 9137 4604
rect 8996 4564 9002 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4604 9367 4607
rect 9398 4604 9404 4616
rect 9355 4576 9404 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 10502 4564 10508 4616
rect 10560 4564 10566 4616
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 9214 4536 9220 4548
rect 8904 4508 9220 4536
rect 8904 4496 8910 4508
rect 9214 4496 9220 4508
rect 9272 4536 9278 4548
rect 9953 4539 10011 4545
rect 9953 4536 9965 4539
rect 9272 4508 9965 4536
rect 9272 4496 9278 4508
rect 9953 4505 9965 4508
rect 9999 4536 10011 4539
rect 10612 4536 10640 4567
rect 9999 4508 10640 4536
rect 10796 4536 10824 4567
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 11204 4576 11437 4604
rect 11204 4564 11210 4576
rect 11425 4573 11437 4576
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4604 11667 4607
rect 11698 4604 11704 4616
rect 11655 4576 11704 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 10962 4536 10968 4548
rect 10796 4508 10968 4536
rect 9999 4505 10011 4508
rect 9953 4499 10011 4505
rect 10962 4496 10968 4508
rect 11020 4536 11026 4548
rect 11624 4536 11652 4567
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 13998 4604 14004 4616
rect 13959 4576 14004 4604
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14093 4607 14151 4613
rect 14093 4573 14105 4607
rect 14139 4573 14151 4607
rect 14918 4604 14924 4616
rect 14879 4576 14924 4604
rect 14093 4567 14151 4573
rect 11020 4508 11652 4536
rect 13265 4539 13323 4545
rect 11020 4496 11026 4508
rect 13265 4505 13277 4539
rect 13311 4536 13323 4539
rect 14108 4536 14136 4567
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 15286 4604 15292 4616
rect 15247 4576 15292 4604
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 13311 4508 14136 4536
rect 13311 4505 13323 4508
rect 13265 4499 13323 4505
rect 9769 4471 9827 4477
rect 9769 4468 9781 4471
rect 8772 4440 9781 4468
rect 9769 4437 9781 4440
rect 9815 4468 9827 4471
rect 9858 4468 9864 4480
rect 9815 4440 9864 4468
rect 9815 4437 9827 4440
rect 9769 4431 9827 4437
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 12158 4428 12164 4480
rect 12216 4468 12222 4480
rect 12618 4468 12624 4480
rect 12216 4440 12624 4468
rect 12216 4428 12222 4440
rect 12618 4428 12624 4440
rect 12676 4468 12682 4480
rect 13280 4468 13308 4499
rect 12676 4440 13308 4468
rect 12676 4428 12682 4440
rect 1104 4378 16008 4400
rect 1104 4326 3480 4378
rect 3532 4326 3544 4378
rect 3596 4326 3608 4378
rect 3660 4326 3672 4378
rect 3724 4326 8478 4378
rect 8530 4326 8542 4378
rect 8594 4326 8606 4378
rect 8658 4326 8670 4378
rect 8722 4326 13475 4378
rect 13527 4326 13539 4378
rect 13591 4326 13603 4378
rect 13655 4326 13667 4378
rect 13719 4326 16008 4378
rect 1104 4304 16008 4326
rect 2869 4267 2927 4273
rect 2869 4233 2881 4267
rect 2915 4264 2927 4267
rect 3234 4264 3240 4276
rect 2915 4236 3240 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 4338 4264 4344 4276
rect 4299 4236 4344 4264
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 4893 4267 4951 4273
rect 4893 4264 4905 4267
rect 4672 4236 4905 4264
rect 4672 4224 4678 4236
rect 4893 4233 4905 4236
rect 4939 4233 4951 4267
rect 4893 4227 4951 4233
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 5040 4236 5764 4264
rect 5040 4224 5046 4236
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 4801 4199 4859 4205
rect 4801 4196 4813 4199
rect 4764 4168 4813 4196
rect 4764 4156 4770 4168
rect 4801 4165 4813 4168
rect 4847 4196 4859 4199
rect 5626 4196 5632 4208
rect 4847 4168 5632 4196
rect 4847 4165 4859 4168
rect 4801 4159 4859 4165
rect 5626 4156 5632 4168
rect 5684 4156 5690 4208
rect 5736 4196 5764 4236
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 7282 4264 7288 4276
rect 5868 4236 5913 4264
rect 7243 4236 7288 4264
rect 5868 4224 5874 4236
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 9766 4264 9772 4276
rect 7392 4236 9772 4264
rect 7392 4196 7420 4236
rect 9766 4224 9772 4236
rect 9824 4264 9830 4276
rect 10410 4264 10416 4276
rect 9824 4236 10416 4264
rect 9824 4224 9830 4236
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 11517 4267 11575 4273
rect 10836 4236 11468 4264
rect 10836 4224 10842 4236
rect 5736 4168 7420 4196
rect 7561 4199 7619 4205
rect 7561 4165 7573 4199
rect 7607 4196 7619 4199
rect 8386 4196 8392 4208
rect 7607 4168 8392 4196
rect 7607 4165 7619 4168
rect 7561 4159 7619 4165
rect 8386 4156 8392 4168
rect 8444 4196 8450 4208
rect 9490 4196 9496 4208
rect 8444 4168 9496 4196
rect 8444 4156 8450 4168
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 10134 4156 10140 4208
rect 10192 4196 10198 4208
rect 11146 4196 11152 4208
rect 10192 4168 11152 4196
rect 10192 4156 10198 4168
rect 11146 4156 11152 4168
rect 11204 4196 11210 4208
rect 11333 4199 11391 4205
rect 11333 4196 11345 4199
rect 11204 4168 11345 4196
rect 11204 4156 11210 4168
rect 11333 4165 11345 4168
rect 11379 4165 11391 4199
rect 11333 4159 11391 4165
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1489 4131 1547 4137
rect 1489 4128 1501 4131
rect 1452 4100 1501 4128
rect 1452 4088 1458 4100
rect 1489 4097 1501 4100
rect 1535 4097 1547 4131
rect 1489 4091 1547 4097
rect 1504 4060 1532 4091
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5500 4100 5549 4128
rect 5500 4088 5506 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5960 4100 6009 4128
rect 5960 4088 5966 4100
rect 5997 4097 6009 4100
rect 6043 4128 6055 4131
rect 6454 4128 6460 4140
rect 6043 4100 6460 4128
rect 6043 4097 6055 4100
rect 5997 4091 6055 4097
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 7098 4128 7104 4140
rect 7059 4100 7104 4128
rect 7098 4088 7104 4100
rect 7156 4128 7162 4140
rect 7466 4128 7472 4140
rect 7156 4100 7472 4128
rect 7156 4088 7162 4100
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 7892 4100 8125 4128
rect 7892 4088 7898 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 9306 4128 9312 4140
rect 8260 4100 8305 4128
rect 8496 4100 9312 4128
rect 8260 4088 8266 4100
rect 2130 4060 2136 4072
rect 1504 4032 2136 4060
rect 2130 4020 2136 4032
rect 2188 4060 2194 4072
rect 2682 4060 2688 4072
rect 2188 4032 2688 4060
rect 2188 4020 2194 4032
rect 2682 4020 2688 4032
rect 2740 4060 2746 4072
rect 3234 4069 3240 4072
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 2740 4032 2973 4060
rect 2740 4020 2746 4032
rect 2961 4029 2973 4032
rect 3007 4029 3019 4063
rect 3228 4060 3240 4069
rect 3195 4032 3240 4060
rect 2961 4023 3019 4029
rect 3228 4023 3240 4032
rect 3234 4020 3240 4023
rect 3292 4020 3298 4072
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 5776 4032 6193 4060
rect 5776 4020 5782 4032
rect 6181 4029 6193 4032
rect 6227 4060 6239 4063
rect 7926 4060 7932 4072
rect 6227 4032 7932 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8294 4060 8300 4072
rect 8067 4032 8300 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8496 4069 8524 4100
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9824 4100 10057 4128
rect 9824 4088 9830 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10962 4128 10968 4140
rect 10923 4100 10968 4128
rect 10045 4091 10103 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 11241 4131 11299 4137
rect 11241 4097 11253 4131
rect 11287 4128 11299 4131
rect 11440 4128 11468 4236
rect 11517 4233 11529 4267
rect 11563 4264 11575 4267
rect 13262 4264 13268 4276
rect 11563 4236 12296 4264
rect 13223 4236 13268 4264
rect 11563 4233 11575 4236
rect 11517 4227 11575 4233
rect 12158 4196 12164 4208
rect 12084 4168 12164 4196
rect 11287 4100 11468 4128
rect 11287 4097 11299 4100
rect 11241 4091 11299 4097
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4029 8539 4063
rect 8481 4023 8539 4029
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4060 8907 4063
rect 9674 4060 9680 4072
rect 8895 4032 9680 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 11330 4060 11336 4072
rect 9999 4032 11336 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 11440 4060 11468 4100
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 12084 4137 12112 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 12268 4196 12296 4236
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 13998 4264 14004 4276
rect 13959 4236 14004 4264
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 14826 4196 14832 4208
rect 12268 4168 14832 4196
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 12069 4131 12127 4137
rect 12069 4097 12081 4131
rect 12115 4097 12127 4131
rect 12069 4091 12127 4097
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12308 4100 13001 4128
rect 12308 4088 12314 4100
rect 12989 4097 13001 4100
rect 13035 4128 13047 4131
rect 14366 4128 14372 4140
rect 13035 4100 14372 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 14366 4088 14372 4100
rect 14424 4128 14430 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14424 4100 14565 4128
rect 14424 4088 14430 4100
rect 14553 4097 14565 4100
rect 14599 4128 14611 4131
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 14599 4100 15393 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 11900 4060 11928 4088
rect 13262 4060 13268 4072
rect 11440 4032 13268 4060
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13814 4060 13820 4072
rect 13775 4032 13820 4060
rect 13814 4020 13820 4032
rect 13872 4060 13878 4072
rect 14461 4063 14519 4069
rect 14461 4060 14473 4063
rect 13872 4032 14473 4060
rect 13872 4020 13878 4032
rect 14461 4029 14473 4032
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 15197 4063 15255 4069
rect 15197 4029 15209 4063
rect 15243 4060 15255 4063
rect 15286 4060 15292 4072
rect 15243 4032 15292 4060
rect 15243 4029 15255 4032
rect 15197 4023 15255 4029
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 1756 3995 1814 4001
rect 1756 3961 1768 3995
rect 1802 3992 1814 3995
rect 3694 3992 3700 4004
rect 1802 3964 3700 3992
rect 1802 3961 1814 3964
rect 1756 3955 1814 3961
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 6914 3992 6920 4004
rect 4448 3964 6920 3992
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4448 3933 4476 3964
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3992 7067 3995
rect 7558 3992 7564 4004
rect 7055 3964 7564 3992
rect 7055 3961 7067 3964
rect 7009 3955 7067 3961
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 8168 3964 9076 3992
rect 8168 3952 8174 3964
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 4396 3896 4445 3924
rect 4396 3884 4402 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5261 3927 5319 3933
rect 5261 3924 5273 3927
rect 5132 3896 5273 3924
rect 5132 3884 5138 3896
rect 5261 3893 5273 3896
rect 5307 3893 5319 3927
rect 5261 3887 5319 3893
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 5626 3924 5632 3936
rect 5399 3896 5632 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 6270 3924 6276 3936
rect 6231 3896 6276 3924
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6362 3884 6368 3936
rect 6420 3924 6426 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 6420 3896 6469 3924
rect 6420 3884 6426 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 7650 3924 7656 3936
rect 7611 3896 7656 3924
rect 6457 3887 6515 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 9048 3933 9076 3964
rect 9122 3952 9128 4004
rect 9180 3992 9186 4004
rect 10042 3992 10048 4004
rect 9180 3964 10048 3992
rect 9180 3952 9186 3964
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10689 3995 10747 4001
rect 10689 3961 10701 3995
rect 10735 3992 10747 3995
rect 10870 3992 10876 4004
rect 10735 3964 10876 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 10870 3952 10876 3964
rect 10928 3992 10934 4004
rect 13449 3995 13507 4001
rect 13449 3992 13461 3995
rect 10928 3964 13461 3992
rect 10928 3952 10934 3964
rect 13449 3961 13461 3964
rect 13495 3961 13507 3995
rect 16482 3992 16488 4004
rect 13449 3955 13507 3961
rect 13648 3964 16488 3992
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 7800 3896 8677 3924
rect 7800 3884 7806 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 8665 3887 8723 3893
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3893 9091 3927
rect 9306 3924 9312 3936
rect 9267 3896 9312 3924
rect 9033 3887 9091 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9490 3924 9496 3936
rect 9451 3896 9496 3924
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 9858 3924 9864 3936
rect 9819 3896 9864 3924
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10321 3927 10379 3933
rect 10321 3893 10333 3927
rect 10367 3924 10379 3927
rect 10502 3924 10508 3936
rect 10367 3896 10508 3924
rect 10367 3893 10379 3896
rect 10321 3887 10379 3893
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 10781 3927 10839 3933
rect 10781 3924 10793 3927
rect 10652 3896 10793 3924
rect 10652 3884 10658 3896
rect 10781 3893 10793 3896
rect 10827 3893 10839 3927
rect 10781 3887 10839 3893
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 11756 3896 11897 3924
rect 11756 3884 11762 3896
rect 11885 3893 11897 3896
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 11977 3927 12035 3933
rect 11977 3893 11989 3927
rect 12023 3924 12035 3927
rect 12437 3927 12495 3933
rect 12437 3924 12449 3927
rect 12023 3896 12449 3924
rect 12023 3893 12035 3896
rect 11977 3887 12035 3893
rect 12437 3893 12449 3896
rect 12483 3893 12495 3927
rect 12802 3924 12808 3936
rect 12763 3896 12808 3924
rect 12437 3887 12495 3893
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13078 3924 13084 3936
rect 12943 3896 13084 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13078 3884 13084 3896
rect 13136 3884 13142 3936
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13648 3924 13676 3964
rect 16482 3952 16488 3964
rect 16540 3952 16546 4004
rect 13228 3896 13676 3924
rect 14369 3927 14427 3933
rect 13228 3884 13234 3896
rect 14369 3893 14381 3927
rect 14415 3924 14427 3927
rect 14458 3924 14464 3936
rect 14415 3896 14464 3924
rect 14415 3893 14427 3896
rect 14369 3887 14427 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 14829 3927 14887 3933
rect 14829 3924 14841 3927
rect 14700 3896 14841 3924
rect 14700 3884 14706 3896
rect 14829 3893 14841 3896
rect 14875 3893 14887 3927
rect 14829 3887 14887 3893
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15252 3896 15301 3924
rect 15252 3884 15258 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15289 3887 15347 3893
rect 1104 3834 16008 3856
rect 1104 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 10976 3834
rect 11028 3782 11040 3834
rect 11092 3782 11104 3834
rect 11156 3782 11168 3834
rect 11220 3782 16008 3834
rect 1104 3760 16008 3782
rect 2038 3720 2044 3732
rect 1999 3692 2044 3720
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3145 3723 3203 3729
rect 3145 3720 3157 3723
rect 3108 3692 3157 3720
rect 3108 3680 3114 3692
rect 3145 3689 3157 3692
rect 3191 3689 3203 3723
rect 3145 3683 3203 3689
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 5442 3720 5448 3732
rect 3752 3692 5448 3720
rect 3752 3680 3758 3692
rect 5442 3680 5448 3692
rect 5500 3720 5506 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5500 3692 5549 3720
rect 5500 3680 5506 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 5537 3683 5595 3689
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 6880 3692 7665 3720
rect 6880 3680 6886 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 7653 3683 7711 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3689 10103 3723
rect 10502 3720 10508 3732
rect 10463 3692 10508 3720
rect 10045 3683 10103 3689
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 2056 3584 2084 3680
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3652 3571 3655
rect 4154 3652 4160 3664
rect 3559 3624 4160 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 4154 3612 4160 3624
rect 4212 3612 4218 3664
rect 6264 3655 6322 3661
rect 6264 3621 6276 3655
rect 6310 3652 6322 3655
rect 6546 3652 6552 3664
rect 6310 3624 6552 3652
rect 6310 3621 6322 3624
rect 6264 3615 6322 3621
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 10060 3652 10088 3683
rect 10502 3680 10508 3692
rect 10560 3680 10566 3732
rect 11333 3723 11391 3729
rect 11333 3689 11345 3723
rect 11379 3720 11391 3723
rect 11422 3720 11428 3732
rect 11379 3692 11428 3720
rect 11379 3689 11391 3692
rect 11333 3683 11391 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11698 3720 11704 3732
rect 11659 3692 11704 3720
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 12529 3723 12587 3729
rect 12529 3689 12541 3723
rect 12575 3720 12587 3723
rect 13078 3720 13084 3732
rect 12575 3692 13084 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 14458 3680 14464 3732
rect 14516 3720 14522 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14516 3692 14841 3720
rect 14516 3680 14522 3692
rect 14829 3689 14841 3692
rect 14875 3720 14887 3723
rect 15194 3720 15200 3732
rect 14875 3692 15200 3720
rect 14875 3689 14887 3692
rect 14829 3683 14887 3689
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15344 3692 15577 3720
rect 15344 3680 15350 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 15565 3683 15623 3689
rect 11241 3655 11299 3661
rect 11241 3652 11253 3655
rect 10060 3624 11253 3652
rect 11241 3621 11253 3624
rect 11287 3621 11299 3655
rect 12066 3652 12072 3664
rect 12027 3624 12072 3652
rect 11241 3615 11299 3621
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 12250 3612 12256 3664
rect 12308 3652 12314 3664
rect 12308 3624 12388 3652
rect 12308 3612 12314 3624
rect 1627 3556 2084 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 2406 3544 2412 3596
rect 2464 3584 2470 3596
rect 2777 3587 2835 3593
rect 2777 3584 2789 3587
rect 2464 3556 2789 3584
rect 2464 3544 2470 3556
rect 2777 3553 2789 3556
rect 2823 3553 2835 3587
rect 2777 3547 2835 3553
rect 3605 3587 3663 3593
rect 3605 3553 3617 3587
rect 3651 3584 3663 3587
rect 4062 3584 4068 3596
rect 3651 3556 4068 3584
rect 3651 3553 3663 3556
rect 3605 3547 3663 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4430 3593 4436 3596
rect 4424 3584 4436 3593
rect 4391 3556 4436 3584
rect 4424 3547 4436 3556
rect 4430 3544 4436 3547
rect 4488 3544 4494 3596
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5718 3584 5724 3596
rect 5675 3556 5724 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 7469 3587 7527 3593
rect 7469 3553 7481 3587
rect 7515 3584 7527 3587
rect 7558 3584 7564 3596
rect 7515 3556 7564 3584
rect 7515 3553 7527 3556
rect 7469 3547 7527 3553
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 8018 3584 8024 3596
rect 7979 3556 8024 3584
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8288 3587 8346 3593
rect 8288 3553 8300 3587
rect 8334 3584 8346 3587
rect 9398 3584 9404 3596
rect 8334 3556 9404 3584
rect 8334 3553 8346 3556
rect 8288 3547 8346 3553
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3584 10471 3587
rect 10778 3584 10784 3596
rect 10459 3556 10784 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 12084 3584 12112 3612
rect 11992 3556 12112 3584
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 3694 3516 3700 3528
rect 2740 3488 3464 3516
rect 3655 3488 3700 3516
rect 2740 3476 2746 3488
rect 3050 3448 3056 3460
rect 3011 3420 3056 3448
rect 3050 3408 3056 3420
rect 3108 3408 3114 3460
rect 3436 3448 3464 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 4172 3448 4200 3479
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5994 3516 6000 3528
rect 5316 3488 6000 3516
rect 5316 3476 5322 3488
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 9953 3519 10011 3525
rect 9732 3488 9777 3516
rect 9732 3476 9738 3488
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10226 3516 10232 3528
rect 9999 3488 10232 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10686 3516 10692 3528
rect 10647 3488 10692 3516
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10928 3488 11437 3516
rect 10928 3476 10934 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 3436 3420 4200 3448
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5813 3451 5871 3457
rect 5813 3448 5825 3451
rect 5224 3420 5825 3448
rect 5224 3408 5230 3420
rect 5813 3417 5825 3420
rect 5859 3417 5871 3451
rect 5813 3411 5871 3417
rect 9122 3408 9128 3460
rect 9180 3448 9186 3460
rect 9180 3420 9352 3448
rect 9180 3408 9186 3420
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 1765 3383 1823 3389
rect 1765 3380 1777 3383
rect 1452 3352 1777 3380
rect 1452 3340 1458 3352
rect 1765 3349 1777 3352
rect 1811 3349 1823 3383
rect 1765 3343 1823 3349
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2409 3383 2467 3389
rect 2409 3380 2421 3383
rect 2096 3352 2421 3380
rect 2096 3340 2102 3352
rect 2409 3349 2421 3352
rect 2455 3380 2467 3383
rect 6270 3380 6276 3392
rect 2455 3352 6276 3380
rect 2455 3349 2467 3352
rect 2409 3343 2467 3349
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 7374 3380 7380 3392
rect 7335 3352 7380 3380
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7926 3380 7932 3392
rect 7887 3352 7932 3380
rect 7926 3340 7932 3352
rect 7984 3380 7990 3392
rect 8938 3380 8944 3392
rect 7984 3352 8944 3380
rect 7984 3340 7990 3352
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9324 3380 9352 3420
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 11992 3448 12020 3556
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 12360 3525 12388 3624
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 12989 3655 13047 3661
rect 12989 3652 13001 3655
rect 12676 3624 13001 3652
rect 12676 3612 12682 3624
rect 12989 3621 13001 3624
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 12897 3587 12955 3593
rect 12897 3553 12909 3587
rect 12943 3584 12955 3587
rect 13541 3587 13599 3593
rect 13541 3584 13553 3587
rect 12943 3556 13553 3584
rect 12943 3553 12955 3556
rect 12897 3547 12955 3553
rect 13541 3553 13553 3556
rect 13587 3553 13599 3587
rect 13541 3547 13599 3553
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 12124 3488 12173 3516
rect 12124 3476 12130 3488
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3485 12403 3519
rect 12345 3479 12403 3485
rect 12912 3448 12940 3547
rect 13170 3516 13176 3528
rect 13131 3488 13176 3516
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 9640 3420 12020 3448
rect 12268 3420 12940 3448
rect 9640 3408 9646 3420
rect 12268 3392 12296 3420
rect 10318 3380 10324 3392
rect 9324 3352 10324 3380
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10410 3340 10416 3392
rect 10468 3380 10474 3392
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10468 3352 10885 3380
rect 10468 3340 10474 3352
rect 10873 3349 10885 3352
rect 10919 3349 10931 3383
rect 10873 3343 10931 3349
rect 12250 3340 12256 3392
rect 12308 3340 12314 3392
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 13044 3352 13369 3380
rect 13044 3340 13050 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13814 3380 13820 3392
rect 13775 3352 13820 3380
rect 13357 3343 13415 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 1104 3290 16008 3312
rect 1104 3238 3480 3290
rect 3532 3238 3544 3290
rect 3596 3238 3608 3290
rect 3660 3238 3672 3290
rect 3724 3238 8478 3290
rect 8530 3238 8542 3290
rect 8594 3238 8606 3290
rect 8658 3238 8670 3290
rect 8722 3238 13475 3290
rect 13527 3238 13539 3290
rect 13591 3238 13603 3290
rect 13655 3238 13667 3290
rect 13719 3238 16008 3290
rect 1104 3216 16008 3238
rect 2222 3136 2228 3188
rect 2280 3176 2286 3188
rect 3329 3179 3387 3185
rect 3329 3176 3341 3179
rect 2280 3148 3341 3176
rect 2280 3136 2286 3148
rect 3329 3145 3341 3148
rect 3375 3145 3387 3179
rect 4062 3176 4068 3188
rect 4023 3148 4068 3176
rect 3329 3139 3387 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 5074 3176 5080 3188
rect 5035 3148 5080 3176
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 6380 3148 8309 3176
rect 1026 3068 1032 3120
rect 1084 3108 1090 3120
rect 2593 3111 2651 3117
rect 2593 3108 2605 3111
rect 1084 3080 2605 3108
rect 1084 3068 1090 3080
rect 2593 3077 2605 3080
rect 2639 3077 2651 3111
rect 2961 3111 3019 3117
rect 2961 3108 2973 3111
rect 2593 3071 2651 3077
rect 2700 3080 2973 3108
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 1486 2972 1492 2984
rect 1447 2944 1492 2972
rect 1486 2932 1492 2944
rect 1544 2932 1550 2984
rect 2038 2972 2044 2984
rect 1999 2944 2044 2972
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2406 2972 2412 2984
rect 2367 2944 2412 2972
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2498 2932 2504 2984
rect 2556 2972 2562 2984
rect 2700 2972 2728 3080
rect 2961 3077 2973 3080
rect 3007 3077 3019 3111
rect 3970 3108 3976 3120
rect 3931 3080 3976 3108
rect 2961 3071 3019 3077
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 4982 3108 4988 3120
rect 4672 3080 4988 3108
rect 4672 3068 4678 3080
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 6380 3049 6408 3148
rect 8297 3145 8309 3148
rect 8343 3176 8355 3179
rect 8846 3176 8852 3188
rect 8343 3148 8852 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9582 3176 9588 3188
rect 9456 3148 9588 3176
rect 9456 3136 9462 3148
rect 9582 3136 9588 3148
rect 9640 3176 9646 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9640 3148 9873 3176
rect 9640 3136 9646 3148
rect 9861 3145 9873 3148
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 11517 3179 11575 3185
rect 10192 3148 10916 3176
rect 10192 3136 10198 3148
rect 10888 3108 10916 3148
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 12066 3176 12072 3188
rect 11563 3148 12072 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 13170 3176 13176 3188
rect 12584 3148 13176 3176
rect 12584 3136 12590 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 14826 3176 14832 3188
rect 14787 3148 14832 3176
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 12897 3111 12955 3117
rect 12897 3108 12909 3111
rect 10888 3080 12909 3108
rect 12897 3077 12909 3080
rect 12943 3077 12955 3111
rect 12897 3071 12955 3077
rect 4709 3043 4767 3049
rect 4709 3040 4721 3043
rect 4488 3012 4721 3040
rect 4488 3000 4494 3012
rect 4709 3009 4721 3012
rect 4755 3040 4767 3043
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 4755 3012 5641 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 5629 3009 5641 3012
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6595 3012 6960 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 2556 2944 2728 2972
rect 2777 2975 2835 2981
rect 2556 2932 2562 2944
rect 2777 2941 2789 2975
rect 2823 2972 2835 2975
rect 2823 2941 2845 2972
rect 2777 2935 2845 2941
rect 2817 2904 2845 2935
rect 3050 2932 3056 2984
rect 3108 2972 3114 2984
rect 3145 2975 3203 2981
rect 3145 2972 3157 2975
rect 3108 2944 3157 2972
rect 3108 2932 3114 2944
rect 3145 2941 3157 2944
rect 3191 2941 3203 2975
rect 3145 2935 3203 2941
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 4338 2972 4344 2984
rect 3559 2944 4344 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2972 5503 2975
rect 5810 2972 5816 2984
rect 5491 2944 5816 2972
rect 5491 2941 5503 2944
rect 5445 2935 5503 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6052 2944 6837 2972
rect 6052 2932 6058 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6932 2972 6960 3012
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 8076 3012 8493 3040
rect 8076 3000 8082 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 7092 2975 7150 2981
rect 7092 2972 7104 2975
rect 6932 2944 7104 2972
rect 6825 2935 6883 2941
rect 7092 2941 7104 2944
rect 7138 2972 7150 2975
rect 7374 2972 7380 2984
rect 7138 2944 7380 2972
rect 7138 2941 7150 2944
rect 7092 2935 7150 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 8294 2932 8300 2984
rect 8352 2932 8358 2984
rect 3970 2904 3976 2916
rect 2817 2876 3976 2904
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 4433 2907 4491 2913
rect 4433 2873 4445 2907
rect 4479 2904 4491 2907
rect 4614 2904 4620 2916
rect 4479 2876 4620 2904
rect 4479 2873 4491 2876
rect 4433 2867 4491 2873
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 5534 2904 5540 2916
rect 5495 2876 5540 2904
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 8312 2904 8340 2932
rect 5776 2876 8340 2904
rect 8496 2904 8524 3003
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9732 3012 9965 3040
rect 9732 3000 9738 3012
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 9953 3003 10011 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12526 3040 12532 3052
rect 12207 3012 12532 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12676 3012 12725 3040
rect 12676 3000 12682 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 8748 2975 8806 2981
rect 8748 2941 8760 2975
rect 8794 2972 8806 2975
rect 9766 2972 9772 2984
rect 8794 2944 9772 2972
rect 8794 2941 8806 2944
rect 8748 2935 8806 2941
rect 9766 2932 9772 2944
rect 9824 2972 9830 2984
rect 10220 2975 10278 2981
rect 9824 2944 10180 2972
rect 9824 2932 9830 2944
rect 9674 2904 9680 2916
rect 8496 2876 9680 2904
rect 5776 2864 5782 2876
rect 9674 2864 9680 2876
rect 9732 2864 9738 2916
rect 566 2796 572 2848
rect 624 2836 630 2848
rect 2225 2839 2283 2845
rect 2225 2836 2237 2839
rect 624 2808 2237 2836
rect 624 2796 630 2808
rect 2225 2805 2237 2808
rect 2271 2805 2283 2839
rect 2225 2799 2283 2805
rect 2682 2796 2688 2848
rect 2740 2836 2746 2848
rect 3697 2839 3755 2845
rect 3697 2836 3709 2839
rect 2740 2808 3709 2836
rect 2740 2796 2746 2808
rect 3697 2805 3709 2808
rect 3743 2805 3755 2839
rect 3697 2799 3755 2805
rect 4525 2839 4583 2845
rect 4525 2805 4537 2839
rect 4571 2836 4583 2839
rect 4706 2836 4712 2848
rect 4571 2808 4712 2836
rect 4571 2805 4583 2808
rect 4525 2799 4583 2805
rect 4706 2796 4712 2808
rect 4764 2836 4770 2848
rect 4982 2836 4988 2848
rect 4764 2808 4988 2836
rect 4764 2796 4770 2808
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5868 2808 5917 2836
rect 5868 2796 5874 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 6270 2836 6276 2848
rect 6231 2808 6276 2836
rect 5905 2799 5963 2805
rect 6270 2796 6276 2808
rect 6328 2796 6334 2848
rect 6546 2796 6552 2848
rect 6604 2836 6610 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 6604 2808 8217 2836
rect 6604 2796 6610 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 9950 2836 9956 2848
rect 9180 2808 9956 2836
rect 9180 2796 9186 2808
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10152 2836 10180 2944
rect 10220 2941 10232 2975
rect 10266 2972 10278 2975
rect 10686 2972 10692 2984
rect 10266 2944 10692 2972
rect 10266 2941 10278 2944
rect 10220 2935 10278 2941
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 11606 2932 11612 2984
rect 11664 2972 11670 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11664 2944 11897 2972
rect 11664 2932 11670 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11885 2935 11943 2941
rect 11900 2904 11928 2935
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12308 2944 12449 2972
rect 12308 2932 12314 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12894 2932 12900 2984
rect 12952 2972 12958 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12952 2944 13001 2972
rect 12952 2932 12958 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 13814 2972 13820 2984
rect 12989 2935 13047 2941
rect 13096 2944 13820 2972
rect 13096 2904 13124 2944
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14884 2944 15025 2972
rect 14884 2932 14890 2944
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 11900 2876 13124 2904
rect 13170 2864 13176 2916
rect 13228 2913 13234 2916
rect 13228 2907 13292 2913
rect 13228 2873 13246 2907
rect 13280 2873 13292 2907
rect 13228 2867 13292 2873
rect 15289 2907 15347 2913
rect 15289 2873 15301 2907
rect 15335 2904 15347 2907
rect 16942 2904 16948 2916
rect 15335 2876 16948 2904
rect 15335 2873 15347 2876
rect 15289 2867 15347 2873
rect 13228 2864 13234 2867
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 10870 2836 10876 2848
rect 10152 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2836 10934 2848
rect 11333 2839 11391 2845
rect 11333 2836 11345 2839
rect 10928 2808 11345 2836
rect 10928 2796 10934 2808
rect 11333 2805 11345 2808
rect 11379 2805 11391 2839
rect 11333 2799 11391 2805
rect 12897 2839 12955 2845
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 14826 2836 14832 2848
rect 12943 2808 14832 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 14826 2796 14832 2808
rect 14884 2796 14890 2848
rect 1104 2746 16008 2768
rect 1104 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 10976 2746
rect 11028 2694 11040 2746
rect 11092 2694 11104 2746
rect 11156 2694 11168 2746
rect 11220 2694 16008 2746
rect 1104 2672 16008 2694
rect 1489 2635 1547 2641
rect 1489 2601 1501 2635
rect 1535 2632 1547 2635
rect 1578 2632 1584 2644
rect 1535 2604 1584 2632
rect 1535 2601 1547 2604
rect 1489 2595 1547 2601
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 4154 2632 4160 2644
rect 4115 2604 4160 2632
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4430 2592 4436 2644
rect 4488 2632 4494 2644
rect 4706 2632 4712 2644
rect 4488 2604 4712 2632
rect 4488 2592 4494 2604
rect 4706 2592 4712 2604
rect 4764 2632 4770 2644
rect 5626 2632 5632 2644
rect 4764 2604 5488 2632
rect 5587 2604 5632 2632
rect 4764 2592 4770 2604
rect 1596 2505 1624 2592
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 4617 2567 4675 2573
rect 4617 2564 4629 2567
rect 3927 2536 4629 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4617 2533 4629 2536
rect 4663 2564 4675 2567
rect 4890 2564 4896 2576
rect 4663 2536 4896 2564
rect 4663 2533 4675 2536
rect 4617 2527 4675 2533
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2465 1639 2499
rect 2481 2499 2539 2505
rect 2481 2496 2493 2499
rect 1581 2459 1639 2465
rect 2056 2468 2493 2496
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 256 2332 1777 2360
rect 256 2320 262 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 2056 2304 2084 2468
rect 2481 2465 2493 2468
rect 2527 2465 2539 2499
rect 2481 2459 2539 2465
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4571 2468 4936 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 2130 2388 2136 2440
rect 2188 2428 2194 2440
rect 2225 2431 2283 2437
rect 2225 2428 2237 2431
rect 2188 2400 2237 2428
rect 2188 2388 2194 2400
rect 2225 2397 2237 2400
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4908 2428 4936 2468
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 5460 2496 5488 2604
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5997 2635 6055 2641
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 6362 2632 6368 2644
rect 6043 2604 6368 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 6641 2635 6699 2641
rect 6641 2601 6653 2635
rect 6687 2601 6699 2635
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 6641 2595 6699 2601
rect 7944 2604 8217 2632
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 6089 2567 6147 2573
rect 6089 2564 6101 2567
rect 5868 2536 6101 2564
rect 5868 2524 5874 2536
rect 6089 2533 6101 2536
rect 6135 2533 6147 2567
rect 6089 2527 6147 2533
rect 6178 2524 6184 2576
rect 6236 2564 6242 2576
rect 6656 2564 6684 2595
rect 6236 2536 6684 2564
rect 6236 2524 6242 2536
rect 6730 2524 6736 2576
rect 6788 2564 6794 2576
rect 7944 2564 7972 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 8352 2604 8585 2632
rect 8352 2592 8358 2604
rect 8573 2601 8585 2604
rect 8619 2601 8631 2635
rect 8846 2632 8852 2644
rect 8807 2604 8852 2632
rect 8573 2595 8631 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 9217 2635 9275 2641
rect 9217 2601 9229 2635
rect 9263 2632 9275 2635
rect 9490 2632 9496 2644
rect 9263 2604 9496 2632
rect 9263 2601 9275 2604
rect 9217 2595 9275 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 9916 2604 10241 2632
rect 9916 2592 9922 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10229 2595 10287 2601
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11330 2632 11336 2644
rect 11103 2604 11336 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12066 2632 12072 2644
rect 12027 2604 12072 2632
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12621 2635 12679 2641
rect 12216 2604 12388 2632
rect 12216 2592 12222 2604
rect 6788 2536 7972 2564
rect 9309 2567 9367 2573
rect 6788 2524 6794 2536
rect 9309 2533 9321 2567
rect 9355 2564 9367 2567
rect 10410 2564 10416 2576
rect 9355 2536 10416 2564
rect 9355 2533 9367 2536
rect 9309 2527 9367 2533
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 11425 2567 11483 2573
rect 10520 2536 10732 2564
rect 6457 2499 6515 2505
rect 5040 2468 5085 2496
rect 5460 2468 6316 2496
rect 5040 2456 5046 2468
rect 6288 2437 6316 2468
rect 6457 2465 6469 2499
rect 6503 2496 6515 2499
rect 6638 2496 6644 2508
rect 6503 2468 6644 2496
rect 6503 2465 6515 2468
rect 6457 2459 6515 2465
rect 6638 2456 6644 2468
rect 6696 2456 6702 2508
rect 6914 2496 6920 2508
rect 6875 2468 6920 2496
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7282 2496 7288 2508
rect 7243 2468 7288 2496
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 7650 2496 7656 2508
rect 7611 2468 7656 2496
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7984 2468 8033 2496
rect 7984 2456 7990 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8386 2496 8392 2508
rect 8347 2468 8392 2496
rect 8021 2459 8079 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10520 2496 10548 2536
rect 10704 2505 10732 2536
rect 11425 2533 11437 2567
rect 11471 2564 11483 2567
rect 11698 2564 11704 2576
rect 11471 2536 11704 2564
rect 11471 2533 11483 2536
rect 11425 2527 11483 2533
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 12360 2564 12388 2604
rect 12621 2601 12633 2635
rect 12667 2632 12679 2635
rect 12802 2632 12808 2644
rect 12667 2604 12808 2632
rect 12667 2601 12679 2604
rect 12621 2595 12679 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12952 2604 13001 2632
rect 12952 2592 12958 2604
rect 12989 2601 13001 2604
rect 13035 2632 13047 2635
rect 14369 2635 14427 2641
rect 14369 2632 14381 2635
rect 13035 2604 14381 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 14369 2601 14381 2604
rect 14415 2601 14427 2635
rect 14369 2595 14427 2601
rect 12526 2564 12532 2576
rect 12360 2536 12532 2564
rect 12526 2524 12532 2536
rect 12584 2564 12590 2576
rect 13262 2564 13268 2576
rect 12584 2536 13268 2564
rect 12584 2524 12590 2536
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 13725 2567 13783 2573
rect 13725 2533 13737 2567
rect 13771 2564 13783 2567
rect 13906 2564 13912 2576
rect 13771 2536 13912 2564
rect 13771 2533 13783 2536
rect 13725 2527 13783 2533
rect 9815 2468 10548 2496
rect 10597 2499 10655 2505
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 10689 2499 10747 2505
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 10962 2496 10968 2508
rect 10735 2468 10968 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 4764 2400 4809 2428
rect 4908 2400 5365 2428
rect 4764 2388 4770 2400
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2428 6331 2431
rect 6546 2428 6552 2440
rect 6319 2400 6552 2428
rect 6319 2397 6331 2400
rect 6273 2391 6331 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9582 2428 9588 2440
rect 9539 2400 9588 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 5169 2363 5227 2369
rect 5169 2360 5181 2363
rect 3292 2332 5181 2360
rect 3292 2320 3298 2332
rect 5169 2329 5181 2332
rect 5215 2329 5227 2363
rect 5169 2323 5227 2329
rect 5994 2320 6000 2372
rect 6052 2360 6058 2372
rect 7469 2363 7527 2369
rect 7469 2360 7481 2363
rect 6052 2332 7481 2360
rect 6052 2320 6058 2332
rect 7469 2329 7481 2332
rect 7515 2329 7527 2363
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 7469 2323 7527 2329
rect 7668 2332 9965 2360
rect 2038 2292 2044 2304
rect 1999 2264 2044 2292
rect 2038 2252 2044 2264
rect 2096 2252 2102 2304
rect 3605 2295 3663 2301
rect 3605 2261 3617 2295
rect 3651 2292 3663 2295
rect 3878 2292 3884 2304
rect 3651 2264 3884 2292
rect 3651 2261 3663 2264
rect 3605 2255 3663 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 3970 2252 3976 2304
rect 4028 2292 4034 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 4028 2264 7113 2292
rect 4028 2252 4034 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 7282 2252 7288 2304
rect 7340 2292 7346 2304
rect 7668 2292 7696 2332
rect 9953 2329 9965 2332
rect 9999 2329 10011 2363
rect 10612 2360 10640 2459
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2496 11575 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11563 2468 11897 2496
rect 11563 2465 11575 2468
rect 11517 2459 11575 2465
rect 11885 2465 11897 2468
rect 11931 2496 11943 2499
rect 13740 2496 13768 2527
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 11931 2468 13768 2496
rect 11931 2465 11943 2468
rect 11885 2459 11943 2465
rect 10778 2428 10784 2440
rect 10739 2400 10784 2428
rect 10778 2388 10784 2400
rect 10836 2428 10842 2440
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 10836 2400 11621 2428
rect 10836 2388 10842 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 11756 2400 12357 2428
rect 11756 2388 11762 2400
rect 12345 2397 12357 2400
rect 12391 2428 12403 2431
rect 12434 2428 12440 2440
rect 12391 2400 12440 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13262 2428 13268 2440
rect 13223 2400 13268 2428
rect 13081 2391 13139 2397
rect 12158 2360 12164 2372
rect 10612 2332 12164 2360
rect 9953 2323 10011 2329
rect 12158 2320 12164 2332
rect 12216 2320 12222 2372
rect 13096 2360 13124 2391
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 13449 2363 13507 2369
rect 13449 2360 13461 2363
rect 13096 2332 13461 2360
rect 7834 2292 7840 2304
rect 7340 2264 7696 2292
rect 7795 2264 7840 2292
rect 7340 2252 7346 2264
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 9398 2252 9404 2304
rect 9456 2292 9462 2304
rect 13096 2292 13124 2332
rect 13449 2329 13461 2332
rect 13495 2329 13507 2363
rect 13449 2323 13507 2329
rect 14090 2292 14096 2304
rect 9456 2264 13124 2292
rect 14051 2264 14096 2292
rect 9456 2252 9462 2264
rect 14090 2252 14096 2264
rect 14148 2292 14154 2304
rect 14185 2295 14243 2301
rect 14185 2292 14197 2295
rect 14148 2264 14197 2292
rect 14148 2252 14154 2264
rect 14185 2261 14197 2264
rect 14231 2261 14243 2295
rect 14185 2255 14243 2261
rect 1104 2202 16008 2224
rect 1104 2150 3480 2202
rect 3532 2150 3544 2202
rect 3596 2150 3608 2202
rect 3660 2150 3672 2202
rect 3724 2150 8478 2202
rect 8530 2150 8542 2202
rect 8594 2150 8606 2202
rect 8658 2150 8670 2202
rect 8722 2150 13475 2202
rect 13527 2150 13539 2202
rect 13591 2150 13603 2202
rect 13655 2150 13667 2202
rect 13719 2150 16008 2202
rect 1104 2128 16008 2150
rect 4890 2048 4896 2100
rect 4948 2088 4954 2100
rect 7650 2088 7656 2100
rect 4948 2060 7656 2088
rect 4948 2048 4954 2060
rect 7650 2048 7656 2060
rect 7708 2048 7714 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 14090 2088 14096 2100
rect 11020 2060 14096 2088
rect 11020 2048 11026 2060
rect 14090 2048 14096 2060
rect 14148 2048 14154 2100
rect 3878 1980 3884 2032
rect 3936 2020 3942 2032
rect 12066 2020 12072 2032
rect 3936 1992 12072 2020
rect 3936 1980 3942 1992
rect 12066 1980 12072 1992
rect 12124 1980 12130 2032
rect 4982 1776 4988 1828
rect 5040 1816 5046 1828
rect 14734 1816 14740 1828
rect 5040 1788 14740 1816
rect 5040 1776 5046 1788
rect 14734 1776 14740 1788
rect 14792 1776 14798 1828
rect 10318 1504 10324 1556
rect 10376 1544 10382 1556
rect 11514 1544 11520 1556
rect 10376 1516 11520 1544
rect 10376 1504 10382 1516
rect 11514 1504 11520 1516
rect 11572 1504 11578 1556
rect 4338 1436 4344 1488
rect 4396 1476 4402 1488
rect 6730 1476 6736 1488
rect 4396 1448 6736 1476
rect 4396 1436 4402 1448
rect 6730 1436 6736 1448
rect 6788 1436 6794 1488
rect 3510 1368 3516 1420
rect 3568 1408 3574 1420
rect 6178 1408 6184 1420
rect 3568 1380 6184 1408
rect 3568 1368 3574 1380
rect 6178 1368 6184 1380
rect 6236 1368 6242 1420
rect 6454 1368 6460 1420
rect 6512 1408 6518 1420
rect 7834 1408 7840 1420
rect 6512 1380 7840 1408
rect 6512 1368 6518 1380
rect 7834 1368 7840 1380
rect 7892 1368 7898 1420
rect 12434 1368 12440 1420
rect 12492 1408 12498 1420
rect 15654 1408 15660 1420
rect 12492 1380 15660 1408
rect 12492 1368 12498 1380
rect 15654 1368 15660 1380
rect 15712 1368 15718 1420
rect 1854 1300 1860 1352
rect 1912 1340 1918 1352
rect 2498 1340 2504 1352
rect 1912 1312 2504 1340
rect 1912 1300 1918 1312
rect 2498 1300 2504 1312
rect 2556 1300 2562 1352
rect 8570 1096 8576 1148
rect 8628 1136 8634 1148
rect 9122 1136 9128 1148
rect 8628 1108 9128 1136
rect 8628 1096 8634 1108
rect 9122 1096 9128 1108
rect 9180 1096 9186 1148
<< via1 >>
rect 9680 18096 9732 18148
rect 12900 18096 12952 18148
rect 14280 18096 14332 18148
rect 4068 17960 4120 18012
rect 12900 17960 12952 18012
rect 2228 17620 2280 17672
rect 2964 17620 3016 17672
rect 12532 17620 12584 17672
rect 13268 17620 13320 17672
rect 12992 17552 13044 17604
rect 13636 17552 13688 17604
rect 204 17484 256 17536
rect 14372 17484 14424 17536
rect 3480 17382 3532 17434
rect 3544 17382 3596 17434
rect 3608 17382 3660 17434
rect 3672 17382 3724 17434
rect 8478 17382 8530 17434
rect 8542 17382 8594 17434
rect 8606 17382 8658 17434
rect 8670 17382 8722 17434
rect 13475 17382 13527 17434
rect 13539 17382 13591 17434
rect 13603 17382 13655 17434
rect 13667 17382 13719 17434
rect 2780 17280 2832 17332
rect 7104 17280 7156 17332
rect 7564 17280 7616 17332
rect 8208 17280 8260 17332
rect 12808 17280 12860 17332
rect 14372 17323 14424 17332
rect 14372 17289 14381 17323
rect 14381 17289 14415 17323
rect 14415 17289 14424 17323
rect 14372 17280 14424 17289
rect 1492 17212 1544 17264
rect 12624 17212 12676 17264
rect 2504 17144 2556 17196
rect 10140 17144 10192 17196
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11244 17144 11296 17196
rect 11428 17187 11480 17196
rect 11428 17153 11437 17187
rect 11437 17153 11471 17187
rect 11471 17153 11480 17187
rect 11428 17144 11480 17153
rect 4068 17076 4120 17128
rect 3240 17008 3292 17060
rect 6552 17008 6604 17060
rect 6644 17008 6696 17060
rect 8208 17076 8260 17128
rect 7840 17008 7892 17060
rect 14924 17119 14976 17128
rect 2780 16940 2832 16992
rect 4988 16940 5040 16992
rect 5724 16940 5776 16992
rect 6368 16940 6420 16992
rect 7564 16940 7616 16992
rect 8852 16940 8904 16992
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 10508 16983 10560 16992
rect 10508 16949 10517 16983
rect 10517 16949 10551 16983
rect 10551 16949 10560 16983
rect 12440 17008 12492 17060
rect 10508 16940 10560 16949
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 13360 17008 13412 17060
rect 11336 16940 11388 16949
rect 13084 16940 13136 16992
rect 14004 16983 14056 16992
rect 14004 16949 14013 16983
rect 14013 16949 14047 16983
rect 14047 16949 14056 16983
rect 14004 16940 14056 16949
rect 14740 16940 14792 16992
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 10976 16838 11028 16890
rect 11040 16838 11092 16890
rect 11104 16838 11156 16890
rect 11168 16838 11220 16890
rect 1860 16736 1912 16788
rect 2964 16779 3016 16788
rect 2964 16745 2973 16779
rect 2973 16745 3007 16779
rect 3007 16745 3016 16779
rect 2964 16736 3016 16745
rect 3332 16736 3384 16788
rect 4252 16736 4304 16788
rect 5080 16736 5132 16788
rect 5816 16736 5868 16788
rect 6276 16736 6328 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 8300 16736 8352 16788
rect 10140 16779 10192 16788
rect 10140 16745 10149 16779
rect 10149 16745 10183 16779
rect 10183 16745 10192 16779
rect 10140 16736 10192 16745
rect 10324 16736 10376 16788
rect 1768 16711 1820 16720
rect 1768 16677 1777 16711
rect 1777 16677 1811 16711
rect 1811 16677 1820 16711
rect 1768 16668 1820 16677
rect 1492 16643 1544 16652
rect 1492 16609 1501 16643
rect 1501 16609 1535 16643
rect 1535 16609 1544 16643
rect 1492 16600 1544 16609
rect 2320 16600 2372 16652
rect 2872 16668 2924 16720
rect 2780 16643 2832 16652
rect 2780 16609 2789 16643
rect 2789 16609 2823 16643
rect 2823 16609 2832 16643
rect 2780 16600 2832 16609
rect 3240 16600 3292 16652
rect 3332 16600 3384 16652
rect 4804 16600 4856 16652
rect 5172 16600 5224 16652
rect 5540 16600 5592 16652
rect 5816 16600 5868 16652
rect 8760 16668 8812 16720
rect 9128 16668 9180 16720
rect 9496 16668 9548 16720
rect 11428 16736 11480 16788
rect 12624 16736 12676 16788
rect 11152 16668 11204 16720
rect 11244 16668 11296 16720
rect 13176 16711 13228 16720
rect 13176 16677 13185 16711
rect 13185 16677 13219 16711
rect 13219 16677 13228 16711
rect 13176 16668 13228 16677
rect 6368 16643 6420 16652
rect 6368 16609 6377 16643
rect 6377 16609 6411 16643
rect 6411 16609 6420 16643
rect 6368 16600 6420 16609
rect 6736 16643 6788 16652
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 8208 16600 8260 16652
rect 8852 16643 8904 16652
rect 8852 16609 8861 16643
rect 8861 16609 8895 16643
rect 8895 16609 8904 16643
rect 8852 16600 8904 16609
rect 9864 16600 9916 16652
rect 5448 16532 5500 16584
rect 6828 16532 6880 16584
rect 9404 16532 9456 16584
rect 13268 16643 13320 16652
rect 940 16464 992 16516
rect 2596 16396 2648 16448
rect 3884 16464 3936 16516
rect 4528 16464 4580 16516
rect 4620 16464 4672 16516
rect 8944 16464 8996 16516
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 14004 16668 14056 16720
rect 13084 16464 13136 16516
rect 8024 16396 8076 16448
rect 10140 16396 10192 16448
rect 10324 16396 10376 16448
rect 14924 16396 14976 16448
rect 3480 16294 3532 16346
rect 3544 16294 3596 16346
rect 3608 16294 3660 16346
rect 3672 16294 3724 16346
rect 8478 16294 8530 16346
rect 8542 16294 8594 16346
rect 8606 16294 8658 16346
rect 8670 16294 8722 16346
rect 13475 16294 13527 16346
rect 13539 16294 13591 16346
rect 13603 16294 13655 16346
rect 13667 16294 13719 16346
rect 3056 16192 3108 16244
rect 8208 16235 8260 16244
rect 5540 16124 5592 16176
rect 6644 16124 6696 16176
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 3884 15988 3936 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 10048 16192 10100 16244
rect 10416 16192 10468 16244
rect 11612 16192 11664 16244
rect 11888 16192 11940 16244
rect 12440 16235 12492 16244
rect 12440 16201 12449 16235
rect 12449 16201 12483 16235
rect 12483 16201 12492 16235
rect 12440 16192 12492 16201
rect 13176 16192 13228 16244
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 10140 16056 10192 16108
rect 12900 16124 12952 16176
rect 11244 16056 11296 16108
rect 11520 16056 11572 16108
rect 13360 16056 13412 16108
rect 13728 16056 13780 16108
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 7104 15963 7156 15972
rect 7104 15929 7138 15963
rect 7138 15929 7156 15963
rect 7104 15920 7156 15929
rect 8116 15920 8168 15972
rect 2504 15895 2556 15904
rect 2504 15861 2513 15895
rect 2513 15861 2547 15895
rect 2547 15861 2556 15895
rect 2504 15852 2556 15861
rect 2872 15895 2924 15904
rect 2872 15861 2881 15895
rect 2881 15861 2915 15895
rect 2915 15861 2924 15895
rect 2872 15852 2924 15861
rect 3148 15852 3200 15904
rect 3240 15852 3292 15904
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 4804 15852 4856 15904
rect 5172 15852 5224 15904
rect 5448 15852 5500 15904
rect 5724 15852 5776 15904
rect 6276 15895 6328 15904
rect 6276 15861 6285 15895
rect 6285 15861 6319 15895
rect 6319 15861 6328 15895
rect 6276 15852 6328 15861
rect 7196 15852 7248 15904
rect 12164 15988 12216 16040
rect 8944 15920 8996 15972
rect 9128 15920 9180 15972
rect 9220 15920 9272 15972
rect 9680 15920 9732 15972
rect 9404 15852 9456 15904
rect 10232 15895 10284 15904
rect 10232 15861 10241 15895
rect 10241 15861 10275 15895
rect 10275 15861 10284 15895
rect 10232 15852 10284 15861
rect 10416 15852 10468 15904
rect 10692 15852 10744 15904
rect 11152 15920 11204 15972
rect 11796 15920 11848 15972
rect 12716 15852 12768 15904
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 14188 15895 14240 15904
rect 14188 15861 14197 15895
rect 14197 15861 14231 15895
rect 14231 15861 14240 15895
rect 14740 15963 14792 15972
rect 14740 15929 14749 15963
rect 14749 15929 14783 15963
rect 14783 15929 14792 15963
rect 14740 15920 14792 15929
rect 14188 15852 14240 15861
rect 16580 15852 16632 15904
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 10976 15750 11028 15802
rect 11040 15750 11092 15802
rect 11104 15750 11156 15802
rect 11168 15750 11220 15802
rect 5724 15648 5776 15700
rect 7196 15691 7248 15700
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 8024 15691 8076 15700
rect 8024 15657 8033 15691
rect 8033 15657 8067 15691
rect 8067 15657 8076 15691
rect 8024 15648 8076 15657
rect 1768 15623 1820 15632
rect 1768 15589 1777 15623
rect 1777 15589 1811 15623
rect 1811 15589 1820 15623
rect 1768 15580 1820 15589
rect 3976 15580 4028 15632
rect 8208 15580 8260 15632
rect 8576 15648 8628 15700
rect 10508 15691 10560 15700
rect 10508 15657 10517 15691
rect 10517 15657 10551 15691
rect 10551 15657 10560 15691
rect 10508 15648 10560 15657
rect 10692 15648 10744 15700
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 12532 15648 12584 15700
rect 8852 15580 8904 15632
rect 9588 15580 9640 15632
rect 9864 15580 9916 15632
rect 4160 15512 4212 15564
rect 7380 15512 7432 15564
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 8300 15512 8352 15564
rect 8668 15512 8720 15564
rect 3056 15444 3108 15496
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 8852 15487 8904 15496
rect 7104 15376 7156 15428
rect 8484 15376 8536 15428
rect 2964 15308 3016 15360
rect 5448 15308 5500 15360
rect 7656 15308 7708 15360
rect 8208 15308 8260 15360
rect 8852 15453 8861 15487
rect 8861 15453 8895 15487
rect 8895 15453 8904 15487
rect 8852 15444 8904 15453
rect 9036 15512 9088 15564
rect 10232 15580 10284 15632
rect 12164 15580 12216 15632
rect 13084 15580 13136 15632
rect 14096 15648 14148 15700
rect 14832 15648 14884 15700
rect 15292 15691 15344 15700
rect 15292 15657 15301 15691
rect 15301 15657 15335 15691
rect 15335 15657 15344 15691
rect 15292 15648 15344 15657
rect 16120 15580 16172 15632
rect 11060 15487 11112 15496
rect 11060 15453 11069 15487
rect 11069 15453 11103 15487
rect 11103 15453 11112 15487
rect 11060 15444 11112 15453
rect 11428 15444 11480 15496
rect 11520 15444 11572 15496
rect 13176 15555 13228 15564
rect 13176 15521 13210 15555
rect 13210 15521 13228 15555
rect 13176 15512 13228 15521
rect 13728 15512 13780 15564
rect 12624 15444 12676 15496
rect 8760 15376 8812 15428
rect 10048 15376 10100 15428
rect 10416 15376 10468 15428
rect 10876 15376 10928 15428
rect 8944 15308 8996 15360
rect 9588 15308 9640 15360
rect 10324 15308 10376 15360
rect 10784 15308 10836 15360
rect 12164 15376 12216 15428
rect 15016 15512 15068 15564
rect 14096 15444 14148 15496
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 12716 15308 12768 15360
rect 14464 15308 14516 15360
rect 14832 15308 14884 15360
rect 3480 15206 3532 15258
rect 3544 15206 3596 15258
rect 3608 15206 3660 15258
rect 3672 15206 3724 15258
rect 8478 15206 8530 15258
rect 8542 15206 8594 15258
rect 8606 15206 8658 15258
rect 8670 15206 8722 15258
rect 13475 15206 13527 15258
rect 13539 15206 13591 15258
rect 13603 15206 13655 15258
rect 13667 15206 13719 15258
rect 1400 15104 1452 15156
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 6828 15104 6880 15156
rect 572 15036 624 15088
rect 3700 15036 3752 15088
rect 4068 15036 4120 15088
rect 5264 15079 5316 15088
rect 2688 14943 2740 14952
rect 2688 14909 2697 14943
rect 2697 14909 2731 14943
rect 2731 14909 2740 14943
rect 2688 14900 2740 14909
rect 4252 14900 4304 14952
rect 2596 14875 2648 14884
rect 2596 14841 2605 14875
rect 2605 14841 2639 14875
rect 2639 14841 2648 14875
rect 2596 14832 2648 14841
rect 3056 14832 3108 14884
rect 4160 14832 4212 14884
rect 5264 15045 5273 15079
rect 5273 15045 5307 15079
rect 5307 15045 5316 15079
rect 5264 15036 5316 15045
rect 6276 15036 6328 15088
rect 9404 15104 9456 15156
rect 9680 15104 9732 15156
rect 9772 15104 9824 15156
rect 10416 15104 10468 15156
rect 10600 15104 10652 15156
rect 13268 15147 13320 15156
rect 13268 15113 13277 15147
rect 13277 15113 13311 15147
rect 13311 15113 13320 15147
rect 13268 15104 13320 15113
rect 14188 15147 14240 15156
rect 14188 15113 14197 15147
rect 14197 15113 14231 15147
rect 14231 15113 14240 15147
rect 14188 15104 14240 15113
rect 9036 15036 9088 15088
rect 4620 14968 4672 15020
rect 6736 14968 6788 15020
rect 7380 14968 7432 15020
rect 8208 14968 8260 15020
rect 9772 15011 9824 15020
rect 9772 14977 9781 15011
rect 9781 14977 9815 15011
rect 9815 14977 9824 15011
rect 9772 14968 9824 14977
rect 11336 14968 11388 15020
rect 14648 15036 14700 15088
rect 4896 14900 4948 14952
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 8852 14900 8904 14952
rect 9036 14900 9088 14952
rect 6736 14832 6788 14884
rect 9128 14832 9180 14884
rect 9404 14900 9456 14952
rect 11060 14900 11112 14952
rect 11704 14900 11756 14952
rect 12256 14900 12308 14952
rect 13360 14968 13412 15020
rect 14832 15011 14884 15020
rect 14832 14977 14841 15011
rect 14841 14977 14875 15011
rect 14875 14977 14884 15011
rect 14832 14968 14884 14977
rect 15016 15011 15068 15020
rect 15016 14977 15025 15011
rect 15025 14977 15059 15011
rect 15059 14977 15068 15011
rect 15016 14968 15068 14977
rect 13176 14900 13228 14952
rect 12164 14875 12216 14884
rect 3332 14764 3384 14816
rect 4436 14764 4488 14816
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 7932 14764 7984 14816
rect 8300 14764 8352 14816
rect 8760 14807 8812 14816
rect 8760 14773 8769 14807
rect 8769 14773 8803 14807
rect 8803 14773 8812 14807
rect 8760 14764 8812 14773
rect 9312 14764 9364 14816
rect 10140 14807 10192 14816
rect 10140 14773 10149 14807
rect 10149 14773 10183 14807
rect 10183 14773 10192 14807
rect 10140 14764 10192 14773
rect 12164 14841 12173 14875
rect 12173 14841 12207 14875
rect 12207 14841 12216 14875
rect 12164 14832 12216 14841
rect 14464 14832 14516 14884
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 12900 14764 12952 14816
rect 14280 14764 14332 14816
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 10976 14662 11028 14714
rect 11040 14662 11092 14714
rect 11104 14662 11156 14714
rect 11168 14662 11220 14714
rect 3792 14560 3844 14612
rect 3884 14560 3936 14612
rect 5264 14560 5316 14612
rect 5724 14560 5776 14612
rect 6276 14560 6328 14612
rect 7380 14560 7432 14612
rect 7564 14560 7616 14612
rect 7656 14560 7708 14612
rect 9404 14560 9456 14612
rect 12808 14560 12860 14612
rect 2688 14492 2740 14544
rect 4068 14492 4120 14544
rect 4252 14492 4304 14544
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 2872 14356 2924 14408
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 4436 14467 4488 14476
rect 4436 14433 4470 14467
rect 4470 14433 4488 14467
rect 4436 14424 4488 14433
rect 5172 14492 5224 14544
rect 6644 14424 6696 14476
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 8760 14467 8812 14476
rect 8760 14433 8769 14467
rect 8769 14433 8803 14467
rect 8803 14433 8812 14467
rect 8760 14424 8812 14433
rect 8944 14424 8996 14476
rect 6184 14399 6236 14408
rect 2780 14288 2832 14340
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 8208 14356 8260 14408
rect 8852 14399 8904 14408
rect 8852 14365 8861 14399
rect 8861 14365 8895 14399
rect 8895 14365 8904 14399
rect 8852 14356 8904 14365
rect 9128 14424 9180 14476
rect 9312 14424 9364 14476
rect 10508 14492 10560 14544
rect 10600 14492 10652 14544
rect 12164 14492 12216 14544
rect 15016 14492 15068 14544
rect 10416 14424 10468 14476
rect 11244 14424 11296 14476
rect 13176 14467 13228 14476
rect 13176 14433 13185 14467
rect 13185 14433 13219 14467
rect 13219 14433 13228 14467
rect 13176 14424 13228 14433
rect 14372 14399 14424 14408
rect 4160 14220 4212 14272
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 5816 14220 5868 14272
rect 6644 14220 6696 14272
rect 9036 14220 9088 14272
rect 9404 14288 9456 14340
rect 9680 14288 9732 14340
rect 13084 14288 13136 14340
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 15384 14263 15436 14272
rect 15384 14229 15393 14263
rect 15393 14229 15427 14263
rect 15427 14229 15436 14263
rect 15384 14220 15436 14229
rect 3480 14118 3532 14170
rect 3544 14118 3596 14170
rect 3608 14118 3660 14170
rect 3672 14118 3724 14170
rect 8478 14118 8530 14170
rect 8542 14118 8594 14170
rect 8606 14118 8658 14170
rect 8670 14118 8722 14170
rect 13475 14118 13527 14170
rect 13539 14118 13591 14170
rect 13603 14118 13655 14170
rect 13667 14118 13719 14170
rect 3148 14059 3200 14068
rect 3148 14025 3157 14059
rect 3157 14025 3191 14059
rect 3191 14025 3200 14059
rect 3148 14016 3200 14025
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 5540 14016 5592 14068
rect 6368 14016 6420 14068
rect 9772 14059 9824 14068
rect 5172 13948 5224 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 3332 13880 3384 13932
rect 4160 13880 4212 13932
rect 4620 13923 4672 13932
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 5632 13948 5684 14000
rect 6460 13948 6512 14000
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 11336 14016 11388 14068
rect 11520 14016 11572 14068
rect 14372 14016 14424 14068
rect 15016 14016 15068 14068
rect 10140 13948 10192 14000
rect 13176 13948 13228 14000
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 4252 13812 4304 13864
rect 4988 13812 5040 13864
rect 5724 13812 5776 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 9680 13880 9732 13932
rect 12164 13880 12216 13932
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 7564 13812 7616 13864
rect 8116 13812 8168 13864
rect 8392 13855 8444 13864
rect 8392 13821 8401 13855
rect 8401 13821 8435 13855
rect 8435 13821 8444 13855
rect 8392 13812 8444 13821
rect 8944 13812 8996 13864
rect 9036 13812 9088 13864
rect 13268 13812 13320 13864
rect 14832 13948 14884 14000
rect 14740 13812 14792 13864
rect 15016 13855 15068 13864
rect 15016 13821 15034 13855
rect 15034 13821 15068 13855
rect 15016 13812 15068 13821
rect 2964 13744 3016 13796
rect 5816 13744 5868 13796
rect 5908 13744 5960 13796
rect 6644 13744 6696 13796
rect 1492 13676 1544 13728
rect 3240 13676 3292 13728
rect 3608 13676 3660 13728
rect 4528 13676 4580 13728
rect 5632 13719 5684 13728
rect 5632 13685 5641 13719
rect 5641 13685 5675 13719
rect 5675 13685 5684 13719
rect 5632 13676 5684 13685
rect 5724 13676 5776 13728
rect 6828 13676 6880 13728
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 9036 13676 9088 13728
rect 10784 13676 10836 13728
rect 12164 13744 12216 13796
rect 13728 13744 13780 13796
rect 12348 13676 12400 13728
rect 13360 13676 13412 13728
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 10976 13574 11028 13626
rect 11040 13574 11092 13626
rect 11104 13574 11156 13626
rect 11168 13574 11220 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 5540 13472 5592 13524
rect 8944 13515 8996 13524
rect 3056 13404 3108 13456
rect 3976 13404 4028 13456
rect 4528 13404 4580 13456
rect 6368 13404 6420 13456
rect 6828 13404 6880 13456
rect 7932 13404 7984 13456
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 11612 13472 11664 13524
rect 12716 13472 12768 13524
rect 13360 13515 13412 13524
rect 13360 13481 13369 13515
rect 13369 13481 13403 13515
rect 13403 13481 13412 13515
rect 13360 13472 13412 13481
rect 9680 13404 9732 13456
rect 1492 13379 1544 13388
rect 1492 13345 1501 13379
rect 1501 13345 1535 13379
rect 1535 13345 1544 13379
rect 1492 13336 1544 13345
rect 5356 13336 5408 13388
rect 9128 13336 9180 13388
rect 11336 13404 11388 13456
rect 11520 13404 11572 13456
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2412 13268 2464 13320
rect 4160 13268 4212 13320
rect 4252 13268 4304 13320
rect 4528 13268 4580 13320
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 3608 13200 3660 13252
rect 10600 13336 10652 13388
rect 11520 13268 11572 13320
rect 12532 13268 12584 13320
rect 13084 13268 13136 13320
rect 13728 13268 13780 13320
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 7288 13175 7340 13184
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7932 13132 7984 13184
rect 12256 13200 12308 13252
rect 12900 13243 12952 13252
rect 12900 13209 12909 13243
rect 12909 13209 12943 13243
rect 12943 13209 12952 13243
rect 12900 13200 12952 13209
rect 8944 13132 8996 13184
rect 9128 13132 9180 13184
rect 11704 13132 11756 13184
rect 3480 13030 3532 13082
rect 3544 13030 3596 13082
rect 3608 13030 3660 13082
rect 3672 13030 3724 13082
rect 8478 13030 8530 13082
rect 8542 13030 8594 13082
rect 8606 13030 8658 13082
rect 8670 13030 8722 13082
rect 13475 13030 13527 13082
rect 13539 13030 13591 13082
rect 13603 13030 13655 13082
rect 13667 13030 13719 13082
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 2412 12928 2464 12937
rect 2780 12928 2832 12980
rect 3884 12928 3936 12980
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 6644 12928 6696 12980
rect 8852 12928 8904 12980
rect 9956 12928 10008 12980
rect 10416 12928 10468 12980
rect 10508 12928 10560 12980
rect 6184 12903 6236 12912
rect 1584 12792 1636 12844
rect 6184 12869 6193 12903
rect 6193 12869 6227 12903
rect 6227 12869 6236 12903
rect 6184 12860 6236 12869
rect 7196 12860 7248 12912
rect 7472 12860 7524 12912
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 5632 12792 5684 12844
rect 4988 12724 5040 12776
rect 5356 12724 5408 12776
rect 6460 12792 6512 12844
rect 7012 12792 7064 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 10508 12792 10560 12844
rect 10784 12792 10836 12844
rect 12440 12860 12492 12912
rect 13176 12860 13228 12912
rect 14004 12928 14056 12980
rect 14464 12860 14516 12912
rect 11612 12835 11664 12844
rect 11612 12801 11621 12835
rect 11621 12801 11655 12835
rect 11655 12801 11664 12835
rect 11612 12792 11664 12801
rect 12348 12792 12400 12844
rect 16948 12792 17000 12844
rect 3516 12699 3568 12708
rect 3516 12665 3550 12699
rect 3550 12665 3568 12699
rect 3516 12656 3568 12665
rect 4712 12656 4764 12708
rect 5448 12656 5500 12708
rect 6184 12656 6236 12708
rect 10600 12724 10652 12776
rect 12440 12724 12492 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 14004 12724 14056 12776
rect 7932 12656 7984 12708
rect 2504 12588 2556 12640
rect 3608 12588 3660 12640
rect 4160 12588 4212 12640
rect 6644 12588 6696 12640
rect 6920 12588 6972 12640
rect 7196 12631 7248 12640
rect 7196 12597 7205 12631
rect 7205 12597 7239 12631
rect 7239 12597 7248 12631
rect 7196 12588 7248 12597
rect 7472 12588 7524 12640
rect 8024 12631 8076 12640
rect 8024 12597 8033 12631
rect 8033 12597 8067 12631
rect 8067 12597 8076 12631
rect 8024 12588 8076 12597
rect 8852 12588 8904 12640
rect 9864 12631 9916 12640
rect 9864 12597 9873 12631
rect 9873 12597 9907 12631
rect 9907 12597 9916 12631
rect 9864 12588 9916 12597
rect 10416 12588 10468 12640
rect 10692 12631 10744 12640
rect 10692 12597 10701 12631
rect 10701 12597 10735 12631
rect 10735 12597 10744 12631
rect 12532 12656 12584 12708
rect 12808 12699 12860 12708
rect 12808 12665 12817 12699
rect 12817 12665 12851 12699
rect 12851 12665 12860 12699
rect 12808 12656 12860 12665
rect 10692 12588 10744 12597
rect 12624 12588 12676 12640
rect 12900 12588 12952 12640
rect 14832 12631 14884 12640
rect 14832 12597 14841 12631
rect 14841 12597 14875 12631
rect 14875 12597 14884 12631
rect 14832 12588 14884 12597
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 10976 12486 11028 12538
rect 11040 12486 11092 12538
rect 11104 12486 11156 12538
rect 11168 12486 11220 12538
rect 3608 12427 3660 12436
rect 3608 12393 3617 12427
rect 3617 12393 3651 12427
rect 3651 12393 3660 12427
rect 3608 12384 3660 12393
rect 6736 12384 6788 12436
rect 2044 12248 2096 12300
rect 2872 12316 2924 12368
rect 3240 12316 3292 12368
rect 5356 12316 5408 12368
rect 6276 12316 6328 12368
rect 6460 12316 6512 12368
rect 2780 12248 2832 12300
rect 4712 12248 4764 12300
rect 5816 12248 5868 12300
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 3240 12180 3292 12232
rect 3516 12155 3568 12164
rect 3516 12121 3525 12155
rect 3525 12121 3559 12155
rect 3559 12121 3568 12155
rect 3516 12112 3568 12121
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4068 12044 4120 12096
rect 7104 12248 7156 12300
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 10692 12384 10744 12436
rect 12348 12384 12400 12436
rect 9036 12316 9088 12368
rect 9956 12316 10008 12368
rect 11980 12316 12032 12368
rect 6276 12180 6328 12189
rect 6092 12044 6144 12096
rect 6276 12044 6328 12096
rect 9680 12180 9732 12232
rect 9956 12180 10008 12232
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 9680 12044 9732 12096
rect 10140 12044 10192 12096
rect 10416 12044 10468 12096
rect 10968 12291 11020 12300
rect 10968 12257 11002 12291
rect 11002 12257 11020 12291
rect 10968 12248 11020 12257
rect 13820 12248 13872 12300
rect 14832 12248 14884 12300
rect 12624 12180 12676 12232
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 11336 12044 11388 12096
rect 12256 12044 12308 12096
rect 3480 11942 3532 11994
rect 3544 11942 3596 11994
rect 3608 11942 3660 11994
rect 3672 11942 3724 11994
rect 8478 11942 8530 11994
rect 8542 11942 8594 11994
rect 8606 11942 8658 11994
rect 8670 11942 8722 11994
rect 13475 11942 13527 11994
rect 13539 11942 13591 11994
rect 13603 11942 13655 11994
rect 13667 11942 13719 11994
rect 2780 11883 2832 11892
rect 2780 11849 2789 11883
rect 2789 11849 2823 11883
rect 2823 11849 2832 11883
rect 2780 11840 2832 11849
rect 3792 11840 3844 11892
rect 4344 11840 4396 11892
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 7932 11883 7984 11892
rect 3884 11772 3936 11824
rect 5724 11772 5776 11824
rect 4712 11747 4764 11756
rect 2872 11636 2924 11688
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 5172 11704 5224 11756
rect 6276 11704 6328 11756
rect 7104 11772 7156 11824
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 9680 11883 9732 11892
rect 9680 11849 9689 11883
rect 9689 11849 9723 11883
rect 9723 11849 9732 11883
rect 10600 11883 10652 11892
rect 9680 11840 9732 11849
rect 10600 11849 10609 11883
rect 10609 11849 10643 11883
rect 10643 11849 10652 11883
rect 10600 11840 10652 11849
rect 11428 11840 11480 11892
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 13820 11840 13872 11892
rect 6920 11704 6972 11756
rect 9496 11772 9548 11824
rect 8024 11704 8076 11756
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 9864 11772 9916 11824
rect 10232 11747 10284 11756
rect 10232 11713 10241 11747
rect 10241 11713 10275 11747
rect 10275 11713 10284 11747
rect 10232 11704 10284 11713
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 10968 11704 11020 11756
rect 12348 11704 12400 11756
rect 2964 11568 3016 11620
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 5632 11568 5684 11620
rect 4620 11500 4672 11509
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 7472 11636 7524 11688
rect 8116 11679 8168 11688
rect 8116 11645 8125 11679
rect 8125 11645 8159 11679
rect 8159 11645 8168 11679
rect 8116 11636 8168 11645
rect 10048 11636 10100 11688
rect 10784 11636 10836 11688
rect 11428 11636 11480 11688
rect 11704 11636 11756 11688
rect 12624 11636 12676 11688
rect 9680 11568 9732 11620
rect 6920 11500 6972 11552
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 9496 11500 9548 11552
rect 9864 11500 9916 11552
rect 11336 11500 11388 11552
rect 12072 11500 12124 11552
rect 12348 11500 12400 11552
rect 14188 11500 14240 11552
rect 15752 11500 15804 11552
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 10976 11398 11028 11450
rect 11040 11398 11092 11450
rect 11104 11398 11156 11450
rect 11168 11398 11220 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 4160 11296 4212 11348
rect 4712 11296 4764 11348
rect 5632 11339 5684 11348
rect 5632 11305 5641 11339
rect 5641 11305 5675 11339
rect 5675 11305 5684 11339
rect 5632 11296 5684 11305
rect 6276 11296 6328 11348
rect 7012 11296 7064 11348
rect 7748 11296 7800 11348
rect 9772 11296 9824 11348
rect 10416 11296 10468 11348
rect 11520 11296 11572 11348
rect 3792 11228 3844 11280
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 2780 11092 2832 11144
rect 3332 11092 3384 11144
rect 5724 11160 5776 11212
rect 6460 11228 6512 11280
rect 6552 11228 6604 11280
rect 6828 11228 6880 11280
rect 9036 11228 9088 11280
rect 7564 11160 7616 11212
rect 8852 11160 8904 11212
rect 10876 11228 10928 11280
rect 4068 11135 4120 11144
rect 3240 11024 3292 11076
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 3056 10956 3108 11008
rect 6644 10956 6696 11008
rect 9772 11092 9824 11144
rect 12072 11228 12124 11280
rect 11336 11160 11388 11212
rect 12256 11160 12308 11212
rect 10048 11092 10100 11144
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 10876 11092 10928 11144
rect 11428 11092 11480 11144
rect 7656 10956 7708 11008
rect 8024 10956 8076 11008
rect 10140 11067 10192 11076
rect 9772 10956 9824 11008
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 10784 11024 10836 11076
rect 12440 10956 12492 11008
rect 12624 10956 12676 11008
rect 16120 10999 16172 11008
rect 16120 10965 16129 10999
rect 16129 10965 16163 10999
rect 16163 10965 16172 10999
rect 16120 10956 16172 10965
rect 3480 10854 3532 10906
rect 3544 10854 3596 10906
rect 3608 10854 3660 10906
rect 3672 10854 3724 10906
rect 8478 10854 8530 10906
rect 8542 10854 8594 10906
rect 8606 10854 8658 10906
rect 8670 10854 8722 10906
rect 13475 10854 13527 10906
rect 13539 10854 13591 10906
rect 13603 10854 13655 10906
rect 13667 10854 13719 10906
rect 3332 10752 3384 10804
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 5724 10684 5776 10736
rect 5816 10684 5868 10736
rect 12256 10752 12308 10804
rect 9220 10727 9272 10736
rect 3516 10480 3568 10532
rect 4160 10616 4212 10668
rect 6644 10616 6696 10668
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 6920 10548 6972 10600
rect 7656 10548 7708 10600
rect 7840 10591 7892 10600
rect 7840 10557 7849 10591
rect 7849 10557 7883 10591
rect 7883 10557 7892 10591
rect 7840 10548 7892 10557
rect 9220 10693 9229 10727
rect 9229 10693 9263 10727
rect 9263 10693 9272 10727
rect 9220 10684 9272 10693
rect 9036 10616 9088 10668
rect 9496 10616 9548 10668
rect 12624 10616 12676 10668
rect 9864 10548 9916 10600
rect 5172 10480 5224 10532
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 3608 10412 3660 10464
rect 4344 10412 4396 10464
rect 7932 10412 7984 10464
rect 8760 10480 8812 10532
rect 11336 10548 11388 10600
rect 10692 10480 10744 10532
rect 12808 10480 12860 10532
rect 12992 10523 13044 10532
rect 12992 10489 13026 10523
rect 13026 10489 13044 10523
rect 12992 10480 13044 10489
rect 9772 10412 9824 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 12440 10412 12492 10464
rect 12900 10412 12952 10464
rect 14740 10412 14792 10464
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 10976 10310 11028 10362
rect 11040 10310 11092 10362
rect 11104 10310 11156 10362
rect 11168 10310 11220 10362
rect 2596 10208 2648 10260
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3608 10251 3660 10260
rect 3056 10208 3108 10217
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 3976 10208 4028 10260
rect 4620 10208 4672 10260
rect 5172 10208 5224 10260
rect 8852 10208 8904 10260
rect 13084 10208 13136 10260
rect 14740 10251 14792 10260
rect 5816 10140 5868 10192
rect 6644 10140 6696 10192
rect 3884 10072 3936 10124
rect 4344 10072 4396 10124
rect 5172 10072 5224 10124
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 5632 10072 5684 10124
rect 6460 10072 6512 10124
rect 7104 10072 7156 10124
rect 7932 10072 7984 10124
rect 9864 10072 9916 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 12624 10140 12676 10192
rect 14740 10217 14749 10251
rect 14749 10217 14783 10251
rect 14783 10217 14792 10251
rect 14740 10208 14792 10217
rect 13268 10072 13320 10124
rect 13820 10072 13872 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2964 10004 3016 10056
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 2504 9936 2556 9988
rect 3516 9979 3568 9988
rect 3516 9945 3525 9979
rect 3525 9945 3559 9979
rect 3559 9945 3568 9979
rect 3516 9936 3568 9945
rect 5264 9936 5316 9988
rect 8208 9936 8260 9988
rect 10232 9936 10284 9988
rect 7564 9868 7616 9920
rect 8116 9868 8168 9920
rect 9956 9911 10008 9920
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 9956 9868 10008 9877
rect 11336 10004 11388 10056
rect 12624 10004 12676 10056
rect 12992 9936 13044 9988
rect 13912 9936 13964 9988
rect 10692 9868 10744 9920
rect 13360 9868 13412 9920
rect 14372 9911 14424 9920
rect 14372 9877 14381 9911
rect 14381 9877 14415 9911
rect 14415 9877 14424 9911
rect 14372 9868 14424 9877
rect 3480 9766 3532 9818
rect 3544 9766 3596 9818
rect 3608 9766 3660 9818
rect 3672 9766 3724 9818
rect 8478 9766 8530 9818
rect 8542 9766 8594 9818
rect 8606 9766 8658 9818
rect 8670 9766 8722 9818
rect 13475 9766 13527 9818
rect 13539 9766 13591 9818
rect 13603 9766 13655 9818
rect 13667 9766 13719 9818
rect 3884 9664 3936 9716
rect 7656 9664 7708 9716
rect 4160 9596 4212 9648
rect 4528 9596 4580 9648
rect 5356 9528 5408 9580
rect 5632 9528 5684 9580
rect 4436 9460 4488 9512
rect 4804 9460 4856 9512
rect 5264 9460 5316 9512
rect 5816 9503 5868 9512
rect 5816 9469 5825 9503
rect 5825 9469 5859 9503
rect 5859 9469 5868 9503
rect 5816 9460 5868 9469
rect 8300 9528 8352 9580
rect 9128 9596 9180 9648
rect 9220 9596 9272 9648
rect 9312 9596 9364 9648
rect 9036 9528 9088 9580
rect 9772 9528 9824 9580
rect 4620 9392 4672 9444
rect 5540 9392 5592 9444
rect 3792 9324 3844 9376
rect 5816 9324 5868 9376
rect 8852 9392 8904 9444
rect 6828 9324 6880 9376
rect 8576 9367 8628 9376
rect 8576 9333 8585 9367
rect 8585 9333 8619 9367
rect 8619 9333 8628 9367
rect 8576 9324 8628 9333
rect 9128 9460 9180 9512
rect 9956 9460 10008 9512
rect 9956 9324 10008 9376
rect 10784 9596 10836 9648
rect 11980 9664 12032 9716
rect 12256 9664 12308 9716
rect 12072 9596 12124 9648
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 10876 9460 10928 9512
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 12808 9596 12860 9648
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 13360 9528 13412 9580
rect 13084 9460 13136 9512
rect 14372 9460 14424 9512
rect 12808 9435 12860 9444
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 10508 9324 10560 9333
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13820 9324 13872 9376
rect 16120 9324 16172 9376
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 10976 9222 11028 9274
rect 11040 9222 11092 9274
rect 11104 9222 11156 9274
rect 11168 9222 11220 9274
rect 2044 9120 2096 9172
rect 3792 9052 3844 9104
rect 5172 9120 5224 9172
rect 8576 9163 8628 9172
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 9128 9120 9180 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 9864 9052 9916 9104
rect 10692 9120 10744 9172
rect 12164 9163 12216 9172
rect 11152 9052 11204 9104
rect 12164 9129 12173 9163
rect 12173 9129 12207 9163
rect 12207 9129 12216 9163
rect 12164 9120 12216 9129
rect 12900 9120 12952 9172
rect 13084 9120 13136 9172
rect 14096 9052 14148 9104
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 6184 9027 6236 9036
rect 6184 8993 6218 9027
rect 6218 8993 6236 9027
rect 6184 8984 6236 8993
rect 7656 8984 7708 9036
rect 5816 8916 5868 8968
rect 7104 8848 7156 8900
rect 5724 8780 5776 8832
rect 6184 8780 6236 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 9588 8984 9640 9036
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9772 8916 9824 8968
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 9680 8848 9732 8900
rect 9956 8848 10008 8900
rect 9220 8780 9272 8832
rect 9772 8780 9824 8832
rect 10692 8780 10744 8832
rect 12164 8984 12216 9036
rect 13360 8984 13412 9036
rect 11796 8916 11848 8968
rect 12072 8891 12124 8900
rect 12072 8857 12081 8891
rect 12081 8857 12115 8891
rect 12115 8857 12124 8891
rect 13176 8916 13228 8968
rect 13912 8959 13964 8968
rect 13912 8925 13921 8959
rect 13921 8925 13955 8959
rect 13955 8925 13964 8959
rect 13912 8916 13964 8925
rect 12072 8848 12124 8857
rect 13820 8780 13872 8832
rect 3480 8678 3532 8730
rect 3544 8678 3596 8730
rect 3608 8678 3660 8730
rect 3672 8678 3724 8730
rect 8478 8678 8530 8730
rect 8542 8678 8594 8730
rect 8606 8678 8658 8730
rect 8670 8678 8722 8730
rect 13475 8678 13527 8730
rect 13539 8678 13591 8730
rect 13603 8678 13655 8730
rect 13667 8678 13719 8730
rect 8944 8576 8996 8628
rect 9588 8576 9640 8628
rect 10416 8576 10468 8628
rect 10692 8576 10744 8628
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11428 8576 11480 8628
rect 13176 8576 13228 8628
rect 13912 8576 13964 8628
rect 2780 8440 2832 8492
rect 2044 8415 2096 8424
rect 2044 8381 2053 8415
rect 2053 8381 2087 8415
rect 2087 8381 2096 8415
rect 2044 8372 2096 8381
rect 5816 8508 5868 8560
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 11336 8508 11388 8560
rect 4620 8440 4672 8449
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 4712 8372 4764 8424
rect 5080 8304 5132 8356
rect 3240 8279 3292 8288
rect 3240 8245 3249 8279
rect 3249 8245 3283 8279
rect 3283 8245 3292 8279
rect 3240 8236 3292 8245
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 5264 8415 5316 8424
rect 5264 8381 5273 8415
rect 5273 8381 5307 8415
rect 5307 8381 5316 8415
rect 5264 8372 5316 8381
rect 6000 8372 6052 8424
rect 6368 8372 6420 8424
rect 7104 8415 7156 8424
rect 7104 8381 7138 8415
rect 7138 8381 7156 8415
rect 7104 8372 7156 8381
rect 5816 8304 5868 8356
rect 7472 8236 7524 8288
rect 9128 8440 9180 8492
rect 9220 8440 9272 8492
rect 9404 8372 9456 8424
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 11796 8440 11848 8492
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 11520 8372 11572 8424
rect 12348 8372 12400 8424
rect 13084 8372 13136 8424
rect 10692 8304 10744 8356
rect 11796 8304 11848 8356
rect 8392 8279 8444 8288
rect 8392 8245 8401 8279
rect 8401 8245 8435 8279
rect 8435 8245 8444 8279
rect 8392 8236 8444 8245
rect 8484 8236 8536 8288
rect 8760 8236 8812 8288
rect 9220 8279 9272 8288
rect 9220 8245 9229 8279
rect 9229 8245 9263 8279
rect 9263 8245 9272 8279
rect 9220 8236 9272 8245
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 9864 8236 9916 8288
rect 10876 8236 10928 8288
rect 12256 8236 12308 8288
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 10976 8134 11028 8186
rect 11040 8134 11092 8186
rect 11104 8134 11156 8186
rect 11168 8134 11220 8186
rect 3240 8032 3292 8084
rect 6368 8032 6420 8084
rect 7104 8032 7156 8084
rect 7380 8032 7432 8084
rect 8392 8032 8444 8084
rect 8852 8032 8904 8084
rect 9220 8032 9272 8084
rect 9496 8032 9548 8084
rect 9772 8075 9824 8084
rect 9772 8041 9781 8075
rect 9781 8041 9815 8075
rect 9815 8041 9824 8075
rect 9772 8032 9824 8041
rect 9956 8032 10008 8084
rect 12808 8032 12860 8084
rect 4896 7964 4948 8016
rect 5264 8007 5316 8016
rect 5264 7973 5273 8007
rect 5273 7973 5307 8007
rect 5307 7973 5316 8007
rect 5264 7964 5316 7973
rect 5448 7896 5500 7948
rect 5632 7896 5684 7948
rect 6920 7964 6972 8016
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4620 7828 4672 7880
rect 5724 7760 5776 7812
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 7380 7871 7432 7880
rect 6184 7828 6236 7837
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 8668 7828 8720 7880
rect 9496 7896 9548 7948
rect 12256 8007 12308 8016
rect 12256 7973 12265 8007
rect 12265 7973 12299 8007
rect 12299 7973 12308 8007
rect 12256 7964 12308 7973
rect 10416 7939 10468 7948
rect 10416 7905 10425 7939
rect 10425 7905 10459 7939
rect 10459 7905 10468 7939
rect 10416 7896 10468 7905
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 11704 7939 11756 7948
rect 11704 7905 11713 7939
rect 11713 7905 11747 7939
rect 11747 7905 11756 7939
rect 11704 7896 11756 7905
rect 12624 7896 12676 7948
rect 12808 7896 12860 7948
rect 10140 7828 10192 7880
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 7564 7692 7616 7744
rect 9312 7760 9364 7812
rect 10876 7803 10928 7812
rect 10876 7769 10885 7803
rect 10885 7769 10919 7803
rect 10919 7769 10928 7803
rect 10876 7760 10928 7769
rect 9588 7692 9640 7744
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 3480 7590 3532 7642
rect 3544 7590 3596 7642
rect 3608 7590 3660 7642
rect 3672 7590 3724 7642
rect 8478 7590 8530 7642
rect 8542 7590 8594 7642
rect 8606 7590 8658 7642
rect 8670 7590 8722 7642
rect 13475 7590 13527 7642
rect 13539 7590 13591 7642
rect 13603 7590 13655 7642
rect 13667 7590 13719 7642
rect 4620 7488 4672 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5264 7488 5316 7540
rect 4528 7284 4580 7336
rect 8944 7531 8996 7540
rect 8944 7497 8953 7531
rect 8953 7497 8987 7531
rect 8987 7497 8996 7531
rect 8944 7488 8996 7497
rect 9864 7488 9916 7540
rect 10324 7488 10376 7540
rect 10508 7488 10560 7540
rect 11244 7488 11296 7540
rect 6920 7420 6972 7472
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 2044 7216 2096 7268
rect 7472 7420 7524 7472
rect 8576 7420 8628 7472
rect 7472 7327 7524 7336
rect 7472 7293 7481 7327
rect 7481 7293 7515 7327
rect 7515 7293 7524 7327
rect 7472 7284 7524 7293
rect 8300 7284 8352 7336
rect 8668 7284 8720 7336
rect 9128 7420 9180 7472
rect 9312 7352 9364 7404
rect 10692 7420 10744 7472
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 10876 7352 10928 7404
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 12716 7352 12768 7404
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 13912 7284 13964 7336
rect 6552 7216 6604 7268
rect 6276 7148 6328 7200
rect 8760 7216 8812 7268
rect 9036 7216 9088 7268
rect 7288 7148 7340 7200
rect 7656 7148 7708 7200
rect 9680 7148 9732 7200
rect 12624 7216 12676 7268
rect 9864 7148 9916 7200
rect 10692 7148 10744 7200
rect 13084 7148 13136 7200
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 10976 7046 11028 7098
rect 11040 7046 11092 7098
rect 11104 7046 11156 7098
rect 11168 7046 11220 7098
rect 7656 6944 7708 6996
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 6644 6876 6696 6928
rect 7380 6876 7432 6928
rect 7564 6876 7616 6928
rect 10692 6944 10744 6996
rect 10876 6944 10928 6996
rect 8668 6876 8720 6928
rect 8852 6876 8904 6928
rect 9128 6876 9180 6928
rect 9588 6876 9640 6928
rect 9680 6876 9732 6928
rect 10324 6876 10376 6928
rect 2596 6851 2648 6860
rect 2596 6817 2605 6851
rect 2605 6817 2639 6851
rect 2639 6817 2648 6851
rect 2596 6808 2648 6817
rect 2872 6808 2924 6860
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 6092 6808 6144 6860
rect 6736 6808 6788 6860
rect 7472 6808 7524 6860
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 1676 6672 1728 6724
rect 2504 6672 2556 6724
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 4620 6672 4672 6724
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 9220 6740 9272 6792
rect 9772 6808 9824 6860
rect 12624 6944 12676 6996
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 5816 6672 5868 6724
rect 8576 6672 8628 6724
rect 8760 6672 8812 6724
rect 1492 6604 1544 6656
rect 9220 6604 9272 6656
rect 9864 6604 9916 6656
rect 11336 6740 11388 6792
rect 12992 6740 13044 6792
rect 11336 6604 11388 6656
rect 12072 6604 12124 6656
rect 3480 6502 3532 6554
rect 3544 6502 3596 6554
rect 3608 6502 3660 6554
rect 3672 6502 3724 6554
rect 8478 6502 8530 6554
rect 8542 6502 8594 6554
rect 8606 6502 8658 6554
rect 8670 6502 8722 6554
rect 13475 6502 13527 6554
rect 13539 6502 13591 6554
rect 13603 6502 13655 6554
rect 13667 6502 13719 6554
rect 2044 6400 2096 6452
rect 4620 6443 4672 6452
rect 2504 6332 2556 6384
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 4804 6400 4856 6452
rect 5448 6400 5500 6452
rect 6092 6400 6144 6452
rect 7012 6400 7064 6452
rect 8024 6400 8076 6452
rect 9680 6443 9732 6452
rect 6736 6332 6788 6384
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 9956 6400 10008 6452
rect 10140 6400 10192 6452
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 10600 6332 10652 6384
rect 5724 6307 5776 6316
rect 1400 6128 1452 6180
rect 1676 6239 1728 6248
rect 1676 6205 1699 6239
rect 1699 6205 1728 6239
rect 1676 6196 1728 6205
rect 4252 6196 4304 6248
rect 3424 6128 3476 6180
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 5356 6196 5408 6248
rect 7196 6264 7248 6316
rect 10876 6264 10928 6316
rect 13268 6264 13320 6316
rect 6828 6196 6880 6248
rect 8116 6196 8168 6248
rect 8852 6196 8904 6248
rect 7288 6128 7340 6180
rect 6644 6060 6696 6112
rect 6736 6060 6788 6112
rect 7380 6060 7432 6112
rect 9680 6060 9732 6112
rect 10048 6060 10100 6112
rect 10140 6060 10192 6112
rect 10692 6060 10744 6112
rect 11888 6060 11940 6112
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 10976 5958 11028 6010
rect 11040 5958 11092 6010
rect 11104 5958 11156 6010
rect 11168 5958 11220 6010
rect 2596 5856 2648 5908
rect 2872 5899 2924 5908
rect 2872 5865 2881 5899
rect 2881 5865 2915 5899
rect 2915 5865 2924 5899
rect 2872 5856 2924 5865
rect 1768 5831 1820 5840
rect 1768 5797 1777 5831
rect 1777 5797 1811 5831
rect 1811 5797 1820 5831
rect 1768 5788 1820 5797
rect 4160 5856 4212 5908
rect 5540 5856 5592 5908
rect 7012 5856 7064 5908
rect 7380 5856 7432 5908
rect 11520 5856 11572 5908
rect 4068 5788 4120 5840
rect 1492 5763 1544 5772
rect 1492 5729 1501 5763
rect 1501 5729 1535 5763
rect 1535 5729 1544 5763
rect 1492 5720 1544 5729
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 4252 5788 4304 5840
rect 5264 5788 5316 5840
rect 6644 5788 6696 5840
rect 7840 5788 7892 5840
rect 9036 5788 9088 5840
rect 9680 5831 9732 5840
rect 9680 5797 9689 5831
rect 9689 5797 9723 5831
rect 9723 5797 9732 5831
rect 9864 5831 9916 5840
rect 9680 5788 9732 5797
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 10692 5831 10744 5840
rect 10692 5797 10701 5831
rect 10701 5797 10735 5831
rect 10735 5797 10744 5831
rect 10692 5788 10744 5797
rect 14924 5831 14976 5840
rect 14924 5797 14933 5831
rect 14933 5797 14967 5831
rect 14967 5797 14976 5831
rect 14924 5788 14976 5797
rect 4344 5763 4396 5772
rect 4344 5729 4378 5763
rect 4378 5729 4396 5763
rect 4344 5720 4396 5729
rect 6920 5720 6972 5772
rect 7472 5720 7524 5772
rect 8300 5720 8352 5772
rect 6736 5652 6788 5704
rect 8852 5695 8904 5704
rect 5264 5584 5316 5636
rect 8852 5661 8861 5695
rect 8861 5661 8895 5695
rect 8895 5661 8904 5695
rect 8852 5652 8904 5661
rect 9588 5652 9640 5704
rect 9956 5720 10008 5772
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 11520 5652 11572 5704
rect 8116 5584 8168 5636
rect 10784 5584 10836 5636
rect 6368 5516 6420 5568
rect 6736 5516 6788 5568
rect 8208 5559 8260 5568
rect 8208 5525 8217 5559
rect 8217 5525 8251 5559
rect 8251 5525 8260 5559
rect 8208 5516 8260 5525
rect 8300 5559 8352 5568
rect 8300 5525 8309 5559
rect 8309 5525 8343 5559
rect 8343 5525 8352 5559
rect 9312 5559 9364 5568
rect 8300 5516 8352 5525
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 12716 5516 12768 5568
rect 3480 5414 3532 5466
rect 3544 5414 3596 5466
rect 3608 5414 3660 5466
rect 3672 5414 3724 5466
rect 8478 5414 8530 5466
rect 8542 5414 8594 5466
rect 8606 5414 8658 5466
rect 8670 5414 8722 5466
rect 13475 5414 13527 5466
rect 13539 5414 13591 5466
rect 13603 5414 13655 5466
rect 13667 5414 13719 5466
rect 2504 5312 2556 5364
rect 3332 5312 3384 5364
rect 4160 5312 4212 5364
rect 5172 5312 5224 5364
rect 6920 5355 6972 5364
rect 6920 5321 6929 5355
rect 6929 5321 6963 5355
rect 6963 5321 6972 5355
rect 6920 5312 6972 5321
rect 8024 5312 8076 5364
rect 9588 5312 9640 5364
rect 11428 5312 11480 5364
rect 11704 5312 11756 5364
rect 7840 5244 7892 5296
rect 8116 5244 8168 5296
rect 4344 5176 4396 5228
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 10692 5176 10744 5228
rect 3332 5108 3384 5160
rect 4988 5108 5040 5160
rect 5264 5108 5316 5160
rect 6736 5108 6788 5160
rect 7196 5108 7248 5160
rect 7748 5108 7800 5160
rect 8484 5108 8536 5160
rect 10784 5151 10836 5160
rect 2412 5040 2464 5092
rect 3976 5040 4028 5092
rect 2964 5015 3016 5024
rect 2964 4981 2973 5015
rect 2973 4981 3007 5015
rect 3007 4981 3016 5015
rect 2964 4972 3016 4981
rect 3608 4972 3660 5024
rect 4252 4972 4304 5024
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 5080 5040 5132 5092
rect 5172 4972 5224 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 6920 5040 6972 5092
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 9404 5040 9456 5092
rect 10508 5040 10560 5092
rect 10232 4972 10284 5024
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 10692 5040 10744 5092
rect 11704 5040 11756 5092
rect 12624 5040 12676 5092
rect 12900 5040 12952 5092
rect 14924 5040 14976 5092
rect 10416 4972 10468 4981
rect 14280 4972 14332 5024
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 10976 4870 11028 4922
rect 11040 4870 11092 4922
rect 11104 4870 11156 4922
rect 11168 4870 11220 4922
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 6644 4768 6696 4820
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7748 4768 7800 4820
rect 2320 4743 2372 4752
rect 2320 4709 2329 4743
rect 2329 4709 2363 4743
rect 2363 4709 2372 4743
rect 2320 4700 2372 4709
rect 3608 4743 3660 4752
rect 3608 4709 3617 4743
rect 3617 4709 3651 4743
rect 3651 4709 3660 4743
rect 3608 4700 3660 4709
rect 4896 4700 4948 4752
rect 5080 4700 5132 4752
rect 5172 4700 5224 4752
rect 5356 4700 5408 4752
rect 6736 4700 6788 4752
rect 7288 4700 7340 4752
rect 8024 4700 8076 4752
rect 9128 4768 9180 4820
rect 10416 4768 10468 4820
rect 3056 4675 3108 4684
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 3056 4641 3065 4675
rect 3065 4641 3099 4675
rect 3099 4641 3108 4675
rect 3056 4632 3108 4641
rect 4620 4632 4672 4684
rect 5448 4632 5500 4684
rect 7656 4632 7708 4684
rect 7748 4632 7800 4684
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 4252 4607 4304 4616
rect 3240 4564 3292 4573
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 2964 4496 3016 4548
rect 3976 4496 4028 4548
rect 1584 4428 1636 4480
rect 3332 4428 3384 4480
rect 5264 4564 5316 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7472 4564 7524 4616
rect 8852 4632 8904 4684
rect 9864 4700 9916 4752
rect 9772 4632 9824 4684
rect 10784 4700 10836 4752
rect 10876 4632 10928 4684
rect 12256 4700 12308 4752
rect 14648 4768 14700 4820
rect 12900 4632 12952 4684
rect 14648 4632 14700 4684
rect 14832 4675 14884 4684
rect 14832 4641 14841 4675
rect 14841 4641 14875 4675
rect 14875 4641 14884 4675
rect 14832 4632 14884 4641
rect 4988 4428 5040 4480
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 5632 4496 5684 4548
rect 6460 4496 6512 4548
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 8944 4564 8996 4616
rect 9404 4564 9456 4616
rect 10508 4564 10560 4616
rect 8852 4496 8904 4548
rect 9220 4496 9272 4548
rect 11152 4564 11204 4616
rect 10968 4496 11020 4548
rect 11704 4564 11756 4616
rect 14004 4607 14056 4616
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 9864 4428 9916 4480
rect 12164 4428 12216 4480
rect 12624 4428 12676 4480
rect 3480 4326 3532 4378
rect 3544 4326 3596 4378
rect 3608 4326 3660 4378
rect 3672 4326 3724 4378
rect 8478 4326 8530 4378
rect 8542 4326 8594 4378
rect 8606 4326 8658 4378
rect 8670 4326 8722 4378
rect 13475 4326 13527 4378
rect 13539 4326 13591 4378
rect 13603 4326 13655 4378
rect 13667 4326 13719 4378
rect 3240 4224 3292 4276
rect 4344 4267 4396 4276
rect 4344 4233 4353 4267
rect 4353 4233 4387 4267
rect 4387 4233 4396 4267
rect 4344 4224 4396 4233
rect 4620 4224 4672 4276
rect 4988 4224 5040 4276
rect 4712 4156 4764 4208
rect 5632 4156 5684 4208
rect 5816 4267 5868 4276
rect 5816 4233 5825 4267
rect 5825 4233 5859 4267
rect 5859 4233 5868 4267
rect 7288 4267 7340 4276
rect 5816 4224 5868 4233
rect 7288 4233 7297 4267
rect 7297 4233 7331 4267
rect 7331 4233 7340 4267
rect 7288 4224 7340 4233
rect 9772 4224 9824 4276
rect 10416 4224 10468 4276
rect 10784 4224 10836 4276
rect 8392 4156 8444 4208
rect 9496 4156 9548 4208
rect 10140 4156 10192 4208
rect 11152 4156 11204 4208
rect 1400 4088 1452 4140
rect 5448 4088 5500 4140
rect 5908 4088 5960 4140
rect 6460 4088 6512 4140
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 7472 4088 7524 4140
rect 7840 4088 7892 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 2136 4020 2188 4072
rect 2688 4020 2740 4072
rect 3240 4063 3292 4072
rect 3240 4029 3274 4063
rect 3274 4029 3292 4063
rect 3240 4020 3292 4029
rect 5724 4020 5776 4072
rect 7932 4020 7984 4072
rect 8300 4020 8352 4072
rect 9312 4088 9364 4140
rect 9772 4088 9824 4140
rect 10968 4131 11020 4140
rect 10968 4097 10977 4131
rect 10977 4097 11011 4131
rect 11011 4097 11020 4131
rect 10968 4088 11020 4097
rect 13268 4267 13320 4276
rect 9680 4020 9732 4072
rect 11336 4020 11388 4072
rect 11888 4088 11940 4140
rect 12164 4156 12216 4208
rect 13268 4233 13277 4267
rect 13277 4233 13311 4267
rect 13311 4233 13320 4267
rect 13268 4224 13320 4233
rect 14004 4267 14056 4276
rect 14004 4233 14013 4267
rect 14013 4233 14047 4267
rect 14047 4233 14056 4267
rect 14004 4224 14056 4233
rect 14832 4156 14884 4208
rect 12256 4088 12308 4140
rect 14372 4088 14424 4140
rect 13268 4020 13320 4072
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 13820 4020 13872 4029
rect 15292 4020 15344 4072
rect 3700 3952 3752 4004
rect 4344 3884 4396 3936
rect 6920 3952 6972 4004
rect 7564 3952 7616 4004
rect 8116 3952 8168 4004
rect 5080 3884 5132 3936
rect 5632 3884 5684 3936
rect 6276 3927 6328 3936
rect 6276 3893 6285 3927
rect 6285 3893 6319 3927
rect 6319 3893 6328 3927
rect 6276 3884 6328 3893
rect 6368 3884 6420 3936
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 7748 3884 7800 3936
rect 9128 3952 9180 4004
rect 10048 3952 10100 4004
rect 10876 3952 10928 4004
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 9864 3884 9916 3893
rect 10508 3884 10560 3936
rect 10600 3884 10652 3936
rect 11704 3884 11756 3936
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 13084 3884 13136 3936
rect 13176 3884 13228 3936
rect 16488 3952 16540 4004
rect 14464 3884 14516 3936
rect 14648 3884 14700 3936
rect 15200 3884 15252 3936
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 10976 3782 11028 3834
rect 11040 3782 11092 3834
rect 11104 3782 11156 3834
rect 11168 3782 11220 3834
rect 2044 3723 2096 3732
rect 2044 3689 2053 3723
rect 2053 3689 2087 3723
rect 2087 3689 2096 3723
rect 2044 3680 2096 3689
rect 3056 3680 3108 3732
rect 3700 3680 3752 3732
rect 5448 3680 5500 3732
rect 6828 3680 6880 3732
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 10508 3723 10560 3732
rect 4160 3612 4212 3664
rect 6552 3612 6604 3664
rect 10508 3689 10517 3723
rect 10517 3689 10551 3723
rect 10551 3689 10560 3723
rect 10508 3680 10560 3689
rect 11428 3680 11480 3732
rect 11704 3723 11756 3732
rect 11704 3689 11713 3723
rect 11713 3689 11747 3723
rect 11747 3689 11756 3723
rect 11704 3680 11756 3689
rect 13084 3680 13136 3732
rect 14464 3680 14516 3732
rect 15200 3680 15252 3732
rect 15292 3680 15344 3732
rect 12072 3655 12124 3664
rect 12072 3621 12081 3655
rect 12081 3621 12115 3655
rect 12115 3621 12124 3655
rect 12072 3612 12124 3621
rect 12256 3612 12308 3664
rect 2412 3544 2464 3596
rect 4068 3544 4120 3596
rect 4436 3587 4488 3596
rect 4436 3553 4470 3587
rect 4470 3553 4488 3587
rect 4436 3544 4488 3553
rect 5724 3544 5776 3596
rect 7564 3544 7616 3596
rect 8024 3587 8076 3596
rect 8024 3553 8033 3587
rect 8033 3553 8067 3587
rect 8067 3553 8076 3587
rect 8024 3544 8076 3553
rect 9404 3544 9456 3596
rect 10784 3544 10836 3596
rect 2688 3476 2740 3528
rect 3700 3519 3752 3528
rect 3056 3451 3108 3460
rect 3056 3417 3065 3451
rect 3065 3417 3099 3451
rect 3099 3417 3108 3451
rect 3056 3408 3108 3417
rect 3700 3485 3709 3519
rect 3709 3485 3743 3519
rect 3743 3485 3752 3519
rect 3700 3476 3752 3485
rect 5264 3476 5316 3528
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 10232 3476 10284 3528
rect 10692 3519 10744 3528
rect 10692 3485 10701 3519
rect 10701 3485 10735 3519
rect 10735 3485 10744 3519
rect 10692 3476 10744 3485
rect 10876 3476 10928 3528
rect 5172 3408 5224 3460
rect 9128 3408 9180 3460
rect 1400 3340 1452 3392
rect 2044 3340 2096 3392
rect 6276 3340 6328 3392
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 7932 3383 7984 3392
rect 7932 3349 7941 3383
rect 7941 3349 7975 3383
rect 7975 3349 7984 3383
rect 7932 3340 7984 3349
rect 8944 3340 8996 3392
rect 9588 3408 9640 3460
rect 12072 3476 12124 3528
rect 12624 3612 12676 3664
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 10324 3340 10376 3392
rect 10416 3340 10468 3392
rect 12256 3340 12308 3392
rect 12992 3340 13044 3392
rect 13820 3383 13872 3392
rect 13820 3349 13829 3383
rect 13829 3349 13863 3383
rect 13863 3349 13872 3383
rect 13820 3340 13872 3349
rect 3480 3238 3532 3290
rect 3544 3238 3596 3290
rect 3608 3238 3660 3290
rect 3672 3238 3724 3290
rect 8478 3238 8530 3290
rect 8542 3238 8594 3290
rect 8606 3238 8658 3290
rect 8670 3238 8722 3290
rect 13475 3238 13527 3290
rect 13539 3238 13591 3290
rect 13603 3238 13655 3290
rect 13667 3238 13719 3290
rect 2228 3136 2280 3188
rect 4068 3179 4120 3188
rect 4068 3145 4077 3179
rect 4077 3145 4111 3179
rect 4111 3145 4120 3179
rect 4068 3136 4120 3145
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 1032 3068 1084 3120
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 1492 2975 1544 2984
rect 1492 2941 1501 2975
rect 1501 2941 1535 2975
rect 1535 2941 1544 2975
rect 1492 2932 1544 2941
rect 2044 2975 2096 2984
rect 2044 2941 2053 2975
rect 2053 2941 2087 2975
rect 2087 2941 2096 2975
rect 2044 2932 2096 2941
rect 2412 2975 2464 2984
rect 2412 2941 2421 2975
rect 2421 2941 2455 2975
rect 2455 2941 2464 2975
rect 2412 2932 2464 2941
rect 2504 2932 2556 2984
rect 3976 3111 4028 3120
rect 3976 3077 3985 3111
rect 3985 3077 4019 3111
rect 4019 3077 4028 3111
rect 3976 3068 4028 3077
rect 4620 3068 4672 3120
rect 4988 3111 5040 3120
rect 4988 3077 4997 3111
rect 4997 3077 5031 3111
rect 5031 3077 5040 3111
rect 4988 3068 5040 3077
rect 4436 3000 4488 3052
rect 8852 3136 8904 3188
rect 9404 3136 9456 3188
rect 9588 3136 9640 3188
rect 10140 3136 10192 3188
rect 12072 3136 12124 3188
rect 12532 3136 12584 3188
rect 13176 3136 13228 3188
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 14832 3179 14884 3188
rect 14832 3145 14841 3179
rect 14841 3145 14875 3179
rect 14875 3145 14884 3179
rect 14832 3136 14884 3145
rect 3056 2932 3108 2984
rect 4344 2932 4396 2984
rect 5816 2932 5868 2984
rect 6000 2932 6052 2984
rect 8024 3000 8076 3052
rect 7380 2932 7432 2984
rect 8300 2932 8352 2984
rect 3976 2864 4028 2916
rect 4620 2864 4672 2916
rect 5540 2907 5592 2916
rect 5540 2873 5549 2907
rect 5549 2873 5583 2907
rect 5583 2873 5592 2907
rect 5540 2864 5592 2873
rect 5724 2864 5776 2916
rect 9680 3000 9732 3052
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 12532 3000 12584 3052
rect 12624 3000 12676 3052
rect 9772 2932 9824 2984
rect 9680 2864 9732 2916
rect 572 2796 624 2848
rect 2688 2796 2740 2848
rect 4712 2796 4764 2848
rect 4988 2796 5040 2848
rect 5816 2796 5868 2848
rect 6276 2839 6328 2848
rect 6276 2805 6285 2839
rect 6285 2805 6319 2839
rect 6319 2805 6328 2839
rect 6276 2796 6328 2805
rect 6552 2796 6604 2848
rect 9128 2796 9180 2848
rect 9956 2796 10008 2848
rect 10692 2932 10744 2984
rect 11612 2932 11664 2984
rect 12256 2932 12308 2984
rect 12900 2932 12952 2984
rect 13820 2932 13872 2984
rect 14832 2932 14884 2984
rect 13176 2864 13228 2916
rect 16948 2864 17000 2916
rect 10876 2796 10928 2848
rect 14832 2796 14884 2848
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 10976 2694 11028 2746
rect 11040 2694 11092 2746
rect 11104 2694 11156 2746
rect 11168 2694 11220 2746
rect 1584 2592 1636 2644
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 4436 2592 4488 2644
rect 4712 2592 4764 2644
rect 5632 2635 5684 2644
rect 4896 2524 4948 2576
rect 204 2320 256 2372
rect 2136 2388 2188 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4988 2499 5040 2508
rect 4988 2465 4997 2499
rect 4997 2465 5031 2499
rect 5031 2465 5040 2499
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 6368 2592 6420 2644
rect 5816 2524 5868 2576
rect 6184 2524 6236 2576
rect 6736 2524 6788 2576
rect 8300 2592 8352 2644
rect 8852 2635 8904 2644
rect 8852 2601 8861 2635
rect 8861 2601 8895 2635
rect 8895 2601 8904 2635
rect 8852 2592 8904 2601
rect 9496 2592 9548 2644
rect 9864 2592 9916 2644
rect 11336 2592 11388 2644
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 12164 2592 12216 2644
rect 10416 2524 10468 2576
rect 4988 2456 5040 2465
rect 6644 2456 6696 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 7288 2499 7340 2508
rect 7288 2465 7297 2499
rect 7297 2465 7331 2499
rect 7331 2465 7340 2499
rect 7288 2456 7340 2465
rect 7656 2499 7708 2508
rect 7656 2465 7665 2499
rect 7665 2465 7699 2499
rect 7699 2465 7708 2499
rect 7656 2456 7708 2465
rect 7932 2456 7984 2508
rect 8392 2499 8444 2508
rect 8392 2465 8401 2499
rect 8401 2465 8435 2499
rect 8435 2465 8444 2499
rect 8392 2456 8444 2465
rect 11704 2524 11756 2576
rect 12808 2592 12860 2644
rect 12900 2592 12952 2644
rect 12532 2524 12584 2576
rect 13268 2524 13320 2576
rect 13912 2567 13964 2576
rect 4712 2388 4764 2397
rect 6552 2388 6604 2440
rect 9588 2388 9640 2440
rect 3240 2320 3292 2372
rect 6000 2320 6052 2372
rect 2044 2295 2096 2304
rect 2044 2261 2053 2295
rect 2053 2261 2087 2295
rect 2087 2261 2096 2295
rect 2044 2252 2096 2261
rect 3884 2252 3936 2304
rect 3976 2252 4028 2304
rect 7288 2252 7340 2304
rect 10968 2456 11020 2508
rect 13912 2533 13921 2567
rect 13921 2533 13955 2567
rect 13955 2533 13964 2567
rect 13912 2524 13964 2533
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11704 2388 11756 2440
rect 12440 2388 12492 2440
rect 13268 2431 13320 2440
rect 12164 2320 12216 2372
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 7840 2295 7892 2304
rect 7840 2261 7849 2295
rect 7849 2261 7883 2295
rect 7883 2261 7892 2295
rect 7840 2252 7892 2261
rect 9404 2252 9456 2304
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 3480 2150 3532 2202
rect 3544 2150 3596 2202
rect 3608 2150 3660 2202
rect 3672 2150 3724 2202
rect 8478 2150 8530 2202
rect 8542 2150 8594 2202
rect 8606 2150 8658 2202
rect 8670 2150 8722 2202
rect 13475 2150 13527 2202
rect 13539 2150 13591 2202
rect 13603 2150 13655 2202
rect 13667 2150 13719 2202
rect 4896 2048 4948 2100
rect 7656 2048 7708 2100
rect 10968 2048 11020 2100
rect 14096 2048 14148 2100
rect 3884 1980 3936 2032
rect 12072 1980 12124 2032
rect 4988 1776 5040 1828
rect 14740 1776 14792 1828
rect 10324 1504 10376 1556
rect 11520 1504 11572 1556
rect 4344 1436 4396 1488
rect 6736 1436 6788 1488
rect 3516 1368 3568 1420
rect 6184 1368 6236 1420
rect 6460 1368 6512 1420
rect 7840 1368 7892 1420
rect 12440 1368 12492 1420
rect 15660 1368 15712 1420
rect 1860 1300 1912 1352
rect 2504 1300 2556 1352
rect 8576 1096 8628 1148
rect 9128 1096 9180 1148
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2226 19200 2282 20000
rect 2594 19200 2650 20000
rect 2778 19544 2834 19553
rect 2778 19479 2834 19488
rect 216 17542 244 19200
rect 204 17536 256 17542
rect 204 17478 256 17484
rect 584 15094 612 19200
rect 952 16522 980 19200
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 1412 15162 1440 19200
rect 1780 17762 1808 19200
rect 1780 17734 1900 17762
rect 1766 17640 1822 17649
rect 1766 17575 1822 17584
rect 1492 17264 1544 17270
rect 1492 17206 1544 17212
rect 1504 16658 1532 17206
rect 1780 16726 1808 17575
rect 1872 16794 1900 17734
rect 2240 17678 2268 19200
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1768 16720 1820 16726
rect 1674 16688 1730 16697
rect 1492 16652 1544 16658
rect 1768 16662 1820 16668
rect 1674 16623 1730 16632
rect 2320 16652 2372 16658
rect 1492 16594 1544 16600
rect 1688 16114 1716 16623
rect 2516 16640 2544 17138
rect 2372 16612 2544 16640
rect 2320 16594 2372 16600
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 2516 15910 2544 16612
rect 2608 16454 2636 19200
rect 2792 17338 2820 19479
rect 3054 19200 3110 20000
rect 3422 19200 3478 20000
rect 3882 19200 3938 20000
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5906 19200 5962 20000
rect 6274 19200 6330 20000
rect 6734 19200 6790 20000
rect 7102 19200 7158 20000
rect 7562 19200 7618 20000
rect 7930 19200 7986 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9586 19200 9642 20000
rect 9954 19200 10010 20000
rect 10414 19200 10470 20000
rect 10782 19200 10838 20000
rect 11242 19200 11298 20000
rect 11610 19200 11666 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12898 19200 12954 20000
rect 13266 19200 13322 20000
rect 13634 19200 13690 20000
rect 14094 19200 14150 20000
rect 14462 19200 14518 20000
rect 14922 19200 14978 20000
rect 15290 19200 15346 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 16578 19200 16634 20000
rect 16946 19200 17002 20000
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2792 16658 2820 16934
rect 2976 16794 3004 17614
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2884 15910 2912 16662
rect 3068 16250 3096 19200
rect 3436 17626 3464 19200
rect 3344 17598 3464 17626
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3252 16658 3280 17002
rect 3344 16794 3372 17598
rect 3454 17436 3750 17456
rect 3510 17434 3534 17436
rect 3590 17434 3614 17436
rect 3670 17434 3694 17436
rect 3532 17382 3534 17434
rect 3596 17382 3608 17434
rect 3670 17382 3672 17434
rect 3510 17380 3534 17382
rect 3590 17380 3614 17382
rect 3670 17380 3694 17382
rect 3454 17360 3750 17380
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3240 15904 3292 15910
rect 3344 15892 3372 16594
rect 3896 16522 3924 19200
rect 4066 18592 4122 18601
rect 4066 18527 4122 18536
rect 4080 18018 4108 18527
rect 4068 18012 4120 18018
rect 4068 17954 4120 17960
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3454 16348 3750 16368
rect 3510 16346 3534 16348
rect 3590 16346 3614 16348
rect 3670 16346 3694 16348
rect 3532 16294 3534 16346
rect 3596 16294 3608 16346
rect 3670 16294 3672 16346
rect 3510 16292 3534 16294
rect 3590 16292 3614 16294
rect 3670 16292 3694 16294
rect 3454 16272 3750 16292
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3292 15864 3372 15892
rect 3240 15846 3292 15852
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1780 15638 1808 15671
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 572 15088 624 15094
rect 572 15030 624 15036
rect 1674 14784 1730 14793
rect 1674 14719 1730 14728
rect 1688 13938 1716 14719
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1582 13832 1638 13841
rect 1582 13767 1638 13776
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13394 1532 13670
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1596 12850 1624 13767
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 1688 12889 1716 13262
rect 2424 12986 2452 13262
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 1674 12880 1730 12889
rect 1584 12844 1636 12850
rect 1674 12815 1730 12824
rect 1584 12786 1636 12792
rect 2516 12646 2544 15846
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2688 14952 2740 14958
rect 2594 14920 2650 14929
rect 2688 14894 2740 14900
rect 2594 14855 2596 14864
rect 2648 14855 2650 14864
rect 2596 14826 2648 14832
rect 2700 14550 2728 14894
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2780 14340 2832 14346
rect 2780 14282 2832 14288
rect 2792 13938 2820 14282
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2884 13530 2912 14350
rect 2976 13802 3004 15302
rect 3068 14890 3096 15438
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 3160 14770 3188 15846
rect 3068 14742 3188 14770
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3068 13462 3096 14742
rect 3146 14376 3202 14385
rect 3146 14311 3202 14320
rect 3160 14074 3188 14311
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3252 13734 3280 15846
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3454 15260 3750 15280
rect 3510 15258 3534 15260
rect 3590 15258 3614 15260
rect 3670 15258 3694 15260
rect 3532 15206 3534 15258
rect 3596 15206 3608 15258
rect 3670 15206 3672 15258
rect 3510 15204 3534 15206
rect 3590 15204 3614 15206
rect 3670 15204 3694 15206
rect 3454 15184 3750 15204
rect 3700 15088 3752 15094
rect 3700 15030 3752 15036
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3344 13938 3372 14758
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3528 14385 3556 14418
rect 3514 14376 3570 14385
rect 3514 14311 3570 14320
rect 3712 14260 3740 15030
rect 3804 14618 3832 15438
rect 3896 14618 3924 15982
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3804 14414 3832 14554
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3712 14232 3832 14260
rect 3454 14172 3750 14192
rect 3510 14170 3534 14172
rect 3590 14170 3614 14172
rect 3670 14170 3694 14172
rect 3532 14118 3534 14170
rect 3596 14118 3608 14170
rect 3670 14118 3672 14170
rect 3510 14116 3534 14118
rect 3590 14116 3614 14118
rect 3670 14116 3694 14118
rect 3454 14096 3750 14116
rect 3804 13977 3832 14232
rect 3988 14074 4016 15574
rect 4080 15094 4108 17070
rect 4264 16794 4292 19200
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4632 16522 4660 19200
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4804 16652 4856 16658
rect 5000 16640 5028 16934
rect 5092 16794 5120 19200
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5172 16652 5224 16658
rect 5000 16612 5120 16640
rect 4804 16594 4856 16600
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4540 15910 4568 16458
rect 4816 15910 4844 16594
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4172 15162 4200 15506
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4342 14920 4398 14929
rect 4160 14884 4212 14890
rect 4080 14844 4160 14872
rect 4080 14550 4108 14844
rect 4160 14826 4212 14832
rect 4264 14550 4292 14894
rect 4342 14855 4398 14864
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4264 14362 4292 14486
rect 4080 14334 4292 14362
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3422 13968 3478 13977
rect 3332 13932 3384 13938
rect 3422 13903 3478 13912
rect 3790 13968 3846 13977
rect 3790 13903 3846 13912
rect 3332 13874 3384 13880
rect 3436 13818 3464 13903
rect 3344 13790 3464 13818
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2792 12782 2820 12922
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 3252 12374 3280 12718
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11937 1716 12174
rect 1674 11928 1730 11937
rect 1674 11863 1730 11872
rect 2056 11354 2084 12242
rect 2792 11898 2820 12242
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2792 11150 2820 11834
rect 2884 11694 2912 12310
rect 3252 12238 3280 12310
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1688 10674 1716 10911
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1676 10056 1728 10062
rect 1674 10024 1676 10033
rect 1728 10024 1730 10033
rect 2516 9994 2544 11086
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 10266 2636 10406
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2976 10062 3004 11562
rect 3344 11234 3372 13790
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3620 13258 3648 13670
rect 3976 13456 4028 13462
rect 3974 13424 3976 13433
rect 4028 13424 4030 13433
rect 3974 13359 4030 13368
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3454 13084 3750 13104
rect 3510 13082 3534 13084
rect 3590 13082 3614 13084
rect 3670 13082 3694 13084
rect 3532 13030 3534 13082
rect 3596 13030 3608 13082
rect 3670 13030 3672 13082
rect 3510 13028 3534 13030
rect 3590 13028 3614 13030
rect 3670 13028 3694 13030
rect 3454 13008 3750 13028
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3528 12170 3556 12650
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3620 12442 3648 12582
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3896 12102 3924 12922
rect 4080 12186 4108 14334
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 13938 4200 14214
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4172 13326 4200 13874
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4264 13326 4292 13806
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4172 12646 4200 13262
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3988 12158 4108 12186
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3454 11996 3750 12016
rect 3510 11994 3534 11996
rect 3590 11994 3614 11996
rect 3670 11994 3694 11996
rect 3532 11942 3534 11994
rect 3596 11942 3608 11994
rect 3670 11942 3672 11994
rect 3510 11940 3534 11942
rect 3590 11940 3614 11942
rect 3670 11940 3694 11942
rect 3454 11920 3750 11940
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3804 11286 3832 11834
rect 3896 11830 3924 12038
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3160 11206 3372 11234
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3068 10266 3096 10950
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 1674 9959 1730 9968
rect 2504 9988 2556 9994
rect 2504 9930 2556 9936
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2056 8430 2084 9114
rect 2778 9072 2834 9081
rect 2778 9007 2834 9016
rect 2792 8498 2820 9007
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1780 8129 1808 8298
rect 1766 8120 1822 8129
rect 1766 8055 1822 8064
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1688 7177 1716 7822
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1674 7168 1730 7177
rect 1674 7103 1730 7112
rect 2056 6798 2084 7210
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 1676 6724 1728 6730
rect 1676 6666 1728 6672
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1400 6180 1452 6186
rect 1400 6122 1452 6128
rect 1412 4146 1440 6122
rect 1504 5778 1532 6598
rect 1688 6254 1716 6666
rect 2056 6458 2084 6734
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2516 6390 2544 6666
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1766 6216 1822 6225
rect 1766 6151 1822 6160
rect 1780 5846 1808 6151
rect 2608 5914 2636 6802
rect 2884 5914 2912 6802
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 2870 5808 2926 5817
rect 1492 5772 1544 5778
rect 2870 5743 2926 5752
rect 1492 5714 1544 5720
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 5370 2544 5646
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2318 5264 2374 5273
rect 2318 5199 2374 5208
rect 2332 4758 2360 5199
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 2320 4752 2372 4758
rect 2320 4694 2372 4700
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1032 3120 1084 3126
rect 1032 3062 1084 3068
rect 572 2848 624 2854
rect 572 2790 624 2796
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 800 244 2314
rect 584 800 612 2790
rect 1044 800 1072 3062
rect 1412 800 1440 3334
rect 1490 3088 1546 3097
rect 1490 3023 1546 3032
rect 1504 2990 1532 3023
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1596 2650 1624 4422
rect 1688 4321 1716 4558
rect 1674 4312 1730 4321
rect 1674 4247 1730 4256
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2042 3768 2098 3777
rect 2042 3703 2044 3712
rect 2096 3703 2098 3712
rect 2044 3674 2096 3680
rect 2044 3392 2096 3398
rect 1674 3360 1730 3369
rect 2044 3334 2096 3340
rect 1674 3295 1730 3304
rect 1688 3058 1716 3295
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 2056 2990 2084 3334
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2148 2446 2176 4014
rect 2424 3602 2452 5034
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 2056 1465 2084 2246
rect 2042 1456 2098 1465
rect 2042 1391 2098 1400
rect 1860 1352 1912 1358
rect 1860 1294 1912 1300
rect 1872 800 1900 1294
rect 2240 800 2268 3130
rect 2424 2990 2452 3538
rect 2700 3534 2728 4014
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2884 3448 2912 5743
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4554 3004 4966
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 3068 3738 3096 4626
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3056 3460 3108 3466
rect 2884 3420 3056 3448
rect 3056 3402 3108 3408
rect 3068 2990 3096 3402
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2516 1358 2544 2926
rect 2688 2848 2740 2854
rect 3160 2836 3188 11206
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 10674 3280 11018
rect 3344 10810 3372 11086
rect 3454 10908 3750 10928
rect 3510 10906 3534 10908
rect 3590 10906 3614 10908
rect 3670 10906 3694 10908
rect 3532 10854 3534 10906
rect 3596 10854 3608 10906
rect 3670 10854 3672 10906
rect 3510 10852 3534 10854
rect 3590 10852 3614 10854
rect 3670 10852 3694 10854
rect 3454 10832 3750 10852
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3884 10668 3936 10674
rect 3988 10656 4016 12158
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11150 4108 12038
rect 4356 11898 4384 14855
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14482 4476 14758
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4540 13818 4568 15846
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4632 13938 4660 14962
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4540 13790 4660 13818
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13462 4568 13670
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 4528 13320 4580 13326
rect 4526 13288 4528 13297
rect 4580 13288 4582 13297
rect 4526 13223 4582 13232
rect 4632 13172 4660 13790
rect 4540 13144 4660 13172
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4172 11354 4200 11494
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3936 10628 4016 10656
rect 4080 10656 4108 11086
rect 4160 10668 4212 10674
rect 4080 10628 4160 10656
rect 3884 10610 3936 10616
rect 4160 10610 4212 10616
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3528 9994 3556 10474
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 10266 3648 10406
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3896 10130 3924 10610
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3454 9820 3750 9840
rect 3510 9818 3534 9820
rect 3590 9818 3614 9820
rect 3670 9818 3694 9820
rect 3532 9766 3534 9818
rect 3596 9766 3608 9818
rect 3670 9766 3672 9818
rect 3510 9764 3534 9766
rect 3590 9764 3614 9766
rect 3670 9764 3694 9766
rect 3454 9744 3750 9764
rect 3896 9722 3924 10066
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 9110 3832 9318
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3454 8732 3750 8752
rect 3510 8730 3534 8732
rect 3590 8730 3614 8732
rect 3670 8730 3694 8732
rect 3532 8678 3534 8730
rect 3596 8678 3608 8730
rect 3670 8678 3672 8730
rect 3510 8676 3534 8678
rect 3590 8676 3614 8678
rect 3670 8676 3694 8678
rect 3454 8656 3750 8676
rect 3804 8498 3832 9046
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 8090 3280 8230
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3804 7886 3832 8434
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3454 7644 3750 7664
rect 3510 7642 3534 7644
rect 3590 7642 3614 7644
rect 3670 7642 3694 7644
rect 3532 7590 3534 7642
rect 3596 7590 3608 7642
rect 3670 7590 3672 7642
rect 3510 7588 3534 7590
rect 3590 7588 3614 7590
rect 3670 7588 3694 7590
rect 3454 7568 3750 7588
rect 3454 6556 3750 6576
rect 3510 6554 3534 6556
rect 3590 6554 3614 6556
rect 3670 6554 3694 6556
rect 3532 6502 3534 6554
rect 3596 6502 3608 6554
rect 3670 6502 3672 6554
rect 3510 6500 3534 6502
rect 3590 6500 3614 6502
rect 3670 6500 3694 6502
rect 3454 6480 3750 6500
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3436 5710 3464 6122
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3344 5370 3372 5646
rect 3454 5468 3750 5488
rect 3510 5466 3534 5468
rect 3590 5466 3614 5468
rect 3670 5466 3694 5468
rect 3532 5414 3534 5466
rect 3596 5414 3608 5466
rect 3670 5414 3672 5466
rect 3510 5412 3534 5414
rect 3590 5412 3614 5414
rect 3670 5412 3694 5414
rect 3454 5392 3750 5412
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4282 3280 4558
rect 3344 4486 3372 5102
rect 3988 5098 4016 10202
rect 4356 10130 4384 10406
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4540 9654 4568 13144
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12306 4752 12650
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4632 10266 4660 11494
rect 4724 11354 4752 11698
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4172 5914 4200 9590
rect 4816 9518 4844 15846
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4448 9042 4476 9454
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4436 9036 4488 9042
rect 4488 8996 4568 9024
rect 4436 8978 4488 8984
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4264 5846 4292 6190
rect 4448 5896 4476 8230
rect 4540 7750 4568 8996
rect 4632 8498 4660 9386
rect 4908 8786 4936 14894
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 13870 5028 14758
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5092 12889 5120 16612
rect 5172 16594 5224 16600
rect 5184 15910 5212 16594
rect 5460 16590 5488 19200
rect 5920 17898 5948 19200
rect 5828 17870 5948 17898
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5540 16652 5592 16658
rect 5736 16640 5764 16934
rect 5828 16794 5856 17870
rect 5953 16892 6249 16912
rect 6009 16890 6033 16892
rect 6089 16890 6113 16892
rect 6169 16890 6193 16892
rect 6031 16838 6033 16890
rect 6095 16838 6107 16890
rect 6169 16838 6171 16890
rect 6009 16836 6033 16838
rect 6089 16836 6113 16838
rect 6169 16836 6193 16838
rect 5953 16816 6249 16836
rect 6288 16794 6316 19200
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6380 16658 6408 16934
rect 5816 16652 5868 16658
rect 5736 16612 5816 16640
rect 5540 16594 5592 16600
rect 5816 16594 5868 16600
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5552 16182 5580 16594
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5276 15094 5304 15438
rect 5460 15366 5488 15846
rect 5736 15706 5764 15846
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 5184 14006 5212 14486
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5078 12880 5134 12889
rect 5078 12815 5134 12824
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5000 11898 5028 12718
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4724 8758 4936 8786
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4632 7886 4660 8434
rect 4724 8430 4752 8758
rect 5092 8616 5120 12815
rect 5184 11762 5212 13126
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5184 10266 5212 10474
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5170 10160 5226 10169
rect 5170 10095 5172 10104
rect 5224 10095 5226 10104
rect 5172 10066 5224 10072
rect 5184 9178 5212 10066
rect 5276 9994 5304 14554
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5368 12986 5396 13330
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5368 12374 5396 12718
rect 5460 12714 5488 14894
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5552 13530 5580 14010
rect 5644 14006 5672 14214
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5736 13870 5764 14554
rect 5828 14532 5856 16594
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 5953 15804 6249 15824
rect 6009 15802 6033 15804
rect 6089 15802 6113 15804
rect 6169 15802 6193 15804
rect 6031 15750 6033 15802
rect 6095 15750 6107 15802
rect 6169 15750 6171 15802
rect 6009 15748 6033 15750
rect 6089 15748 6113 15750
rect 6169 15748 6193 15750
rect 5953 15728 6249 15748
rect 6288 15609 6316 15846
rect 6274 15600 6330 15609
rect 6274 15535 6330 15544
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 5953 14716 6249 14736
rect 6009 14714 6033 14716
rect 6089 14714 6113 14716
rect 6169 14714 6193 14716
rect 6031 14662 6033 14714
rect 6095 14662 6107 14714
rect 6169 14662 6171 14714
rect 6009 14660 6033 14662
rect 6089 14660 6113 14662
rect 6169 14660 6193 14662
rect 5953 14640 6249 14660
rect 6288 14618 6316 15030
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 5828 14504 5948 14532
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5828 13802 5856 14214
rect 5920 13802 5948 14504
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13938 6224 14350
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5644 12850 5672 13670
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5356 12368 5408 12374
rect 5736 12356 5764 13670
rect 5953 13628 6249 13648
rect 6009 13626 6033 13628
rect 6089 13626 6113 13628
rect 6169 13626 6193 13628
rect 6031 13574 6033 13626
rect 6095 13574 6107 13626
rect 6169 13574 6171 13626
rect 6009 13572 6033 13574
rect 6089 13572 6113 13574
rect 6169 13572 6193 13574
rect 5953 13552 6249 13572
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5356 12310 5408 12316
rect 5552 12328 5764 12356
rect 5446 10160 5502 10169
rect 5446 10095 5448 10104
rect 5500 10095 5502 10104
rect 5448 10066 5500 10072
rect 5552 10062 5580 12328
rect 5828 12306 5856 13262
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6196 12714 6224 12854
rect 6288 12753 6316 14554
rect 6380 14249 6408 16594
rect 6366 14240 6422 14249
rect 6366 14175 6422 14184
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6380 13462 6408 14010
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6368 13456 6420 13462
rect 6368 13398 6420 13404
rect 6274 12744 6330 12753
rect 6184 12708 6236 12714
rect 6274 12679 6330 12688
rect 6184 12650 6236 12656
rect 5953 12540 6249 12560
rect 6009 12538 6033 12540
rect 6089 12538 6113 12540
rect 6169 12538 6193 12540
rect 6031 12486 6033 12538
rect 6095 12486 6107 12538
rect 6169 12486 6171 12538
rect 6009 12484 6033 12486
rect 6089 12484 6113 12486
rect 6169 12484 6193 12486
rect 5953 12464 6249 12484
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 6288 12238 6316 12310
rect 6276 12232 6328 12238
rect 6104 12192 6276 12220
rect 6104 12102 6132 12192
rect 6276 12174 6328 12180
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5644 11354 5672 11562
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5736 11218 5764 11766
rect 6288 11762 6316 12038
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 5953 11452 6249 11472
rect 6009 11450 6033 11452
rect 6089 11450 6113 11452
rect 6169 11450 6193 11452
rect 6031 11398 6033 11450
rect 6095 11398 6107 11450
rect 6169 11398 6171 11450
rect 6009 11396 6033 11398
rect 6089 11396 6113 11398
rect 6169 11396 6193 11398
rect 5953 11376 6249 11396
rect 6288 11354 6316 11494
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 10742 5764 11154
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4816 8588 5120 8616
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4620 7880 4672 7886
rect 4816 7868 4844 8588
rect 5184 8514 5212 9114
rect 5000 8486 5212 8514
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 8022 4936 8230
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4816 7840 4936 7868
rect 4620 7822 4672 7828
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4540 7342 4568 7686
rect 4632 7546 4660 7822
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4632 6458 4660 6666
rect 4816 6458 4844 6734
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4448 5868 4568 5896
rect 4068 5840 4120 5846
rect 4252 5840 4304 5846
rect 4120 5788 4200 5794
rect 4068 5782 4200 5788
rect 4252 5782 4304 5788
rect 4080 5766 4200 5782
rect 4172 5370 4200 5766
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4356 5234 4384 5714
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3620 4758 3648 4966
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 4264 4622 4292 4966
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3454 4380 3750 4400
rect 3510 4378 3534 4380
rect 3590 4378 3614 4380
rect 3670 4378 3694 4380
rect 3532 4326 3534 4378
rect 3596 4326 3608 4378
rect 3670 4326 3672 4378
rect 3510 4324 3534 4326
rect 3590 4324 3614 4326
rect 3670 4324 3694 4326
rect 3454 4304 3750 4324
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3252 4078 3280 4218
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3712 3738 3740 3946
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3712 3534 3740 3674
rect 3988 3641 4016 4490
rect 4356 4282 4384 5170
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4160 3664 4212 3670
rect 3974 3632 4030 3641
rect 4160 3606 4212 3612
rect 3974 3567 4030 3576
rect 4068 3596 4120 3602
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3454 3292 3750 3312
rect 3510 3290 3534 3292
rect 3590 3290 3614 3292
rect 3670 3290 3694 3292
rect 3532 3238 3534 3290
rect 3596 3238 3608 3290
rect 3670 3238 3672 3290
rect 3510 3236 3534 3238
rect 3590 3236 3614 3238
rect 3670 3236 3694 3238
rect 3454 3216 3750 3236
rect 3988 3126 4016 3567
rect 4068 3538 4120 3544
rect 4080 3194 4108 3538
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3988 2922 4016 3062
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 2688 2790 2740 2796
rect 2976 2808 3188 2836
rect 2504 1352 2556 1358
rect 2504 1294 2556 1300
rect 2700 800 2728 2790
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 2976 513 3004 2808
rect 4172 2650 4200 3606
rect 4356 2990 4384 3878
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4448 3058 4476 3538
rect 4540 3108 4568 5868
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4632 4282 4660 4626
rect 4724 4593 4752 4966
rect 4908 4758 4936 7840
rect 5000 5166 5028 8486
rect 5276 8430 5304 9454
rect 5264 8424 5316 8430
rect 5078 8392 5134 8401
rect 5264 8366 5316 8372
rect 5078 8327 5080 8336
rect 5132 8327 5134 8336
rect 5080 8298 5132 8304
rect 5092 7546 5120 8298
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5276 7546 5304 7958
rect 5080 7540 5132 7546
rect 5264 7540 5316 7546
rect 5132 7500 5212 7528
rect 5080 7482 5132 7488
rect 5184 5930 5212 7500
rect 5264 7482 5316 7488
rect 5368 6254 5396 9522
rect 5552 9450 5580 9998
rect 5644 9586 5672 10066
rect 5736 10062 5764 10678
rect 5828 10198 5856 10678
rect 5953 10364 6249 10384
rect 6009 10362 6033 10364
rect 6089 10362 6113 10364
rect 6169 10362 6193 10364
rect 6031 10310 6033 10362
rect 6095 10310 6107 10362
rect 6169 10310 6171 10362
rect 6009 10308 6033 10310
rect 6089 10308 6113 10310
rect 6169 10308 6193 10310
rect 5953 10288 6249 10308
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5816 9512 5868 9518
rect 5814 9480 5816 9489
rect 5868 9480 5870 9489
rect 5540 9444 5592 9450
rect 5814 9415 5870 9424
rect 5540 9386 5592 9392
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9058 5856 9318
rect 5953 9276 6249 9296
rect 6009 9274 6033 9276
rect 6089 9274 6113 9276
rect 6169 9274 6193 9276
rect 6031 9222 6033 9274
rect 6095 9222 6107 9274
rect 6169 9222 6171 9274
rect 6009 9220 6033 9222
rect 6089 9220 6113 9222
rect 6169 9220 6193 9222
rect 5953 9200 6249 9220
rect 5828 9030 6040 9058
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5460 6458 5488 7890
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5184 5902 5396 5930
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5276 5642 5304 5782
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4710 4584 4766 4593
rect 4710 4519 4766 4528
rect 5000 4486 5028 5102
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5092 4758 5120 5034
rect 5184 5030 5212 5306
rect 5276 5166 5304 5578
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4758 5212 4966
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5276 4622 5304 5102
rect 5368 4758 5396 5902
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5460 4690 5488 6394
rect 5552 5914 5580 6802
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5644 5250 5672 7890
rect 5736 7818 5764 8774
rect 5828 8566 5856 8910
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 6012 8430 6040 9030
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8838 6224 8978
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6380 8430 6408 13398
rect 6472 12850 6500 13942
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6472 11286 6500 12310
rect 6564 11370 6592 17002
rect 6656 16640 6684 17002
rect 6748 16776 6776 19200
rect 7116 17338 7144 19200
rect 7576 17338 7604 19200
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7564 16992 7616 16998
rect 7484 16940 7564 16946
rect 7484 16934 7616 16940
rect 7484 16918 7604 16934
rect 6920 16788 6972 16794
rect 6748 16748 6920 16776
rect 6920 16730 6972 16736
rect 6736 16652 6788 16658
rect 6656 16612 6736 16640
rect 6736 16594 6788 16600
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6656 16017 6684 16118
rect 6642 16008 6698 16017
rect 6642 15943 6698 15952
rect 6748 15026 6776 16594
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6840 16046 6868 16526
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6840 15162 6868 15982
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 7116 15434 7144 15914
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15706 7236 15846
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 14278 6684 14418
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6656 12986 6684 13738
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6656 12646 6684 12922
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6748 12442 6776 14826
rect 6840 13870 6868 15098
rect 7392 15026 7420 15506
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7380 14816 7432 14822
rect 7378 14784 7380 14793
rect 7432 14784 7434 14793
rect 7378 14719 7434 14728
rect 7392 14618 7420 14719
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13462 6868 13670
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6748 11506 6776 12378
rect 6932 11762 6960 12582
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6920 11552 6972 11558
rect 6748 11478 6868 11506
rect 6920 11494 6972 11500
rect 7024 11506 7052 12786
rect 7208 12646 7236 12854
rect 7300 12850 7328 13126
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7392 12730 7420 14554
rect 7484 13190 7512 16918
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7576 14618 7604 15506
rect 7746 15464 7802 15473
rect 7746 15399 7802 15408
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 14618 7696 15302
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 13326 7604 13806
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12918 7512 13126
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7300 12702 7420 12730
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7116 11830 7144 12242
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 6564 11342 6776 11370
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6472 10130 6500 11222
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6564 10010 6592 11222
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10674 6684 10950
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6656 10198 6684 10610
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6472 9982 6592 10010
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6322 5764 6734
rect 5828 6730 5856 8298
rect 5953 8188 6249 8208
rect 6009 8186 6033 8188
rect 6089 8186 6113 8188
rect 6169 8186 6193 8188
rect 6031 8134 6033 8186
rect 6095 8134 6107 8186
rect 6169 8134 6171 8186
rect 6009 8132 6033 8134
rect 6089 8132 6113 8134
rect 6169 8132 6193 8134
rect 5953 8112 6249 8132
rect 6380 8090 6408 8366
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6196 7410 6224 7822
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 5953 7100 6249 7120
rect 6009 7098 6033 7100
rect 6089 7098 6113 7100
rect 6169 7098 6193 7100
rect 6031 7046 6033 7098
rect 6095 7046 6107 7098
rect 6169 7046 6171 7098
rect 6009 7044 6033 7046
rect 6089 7044 6113 7046
rect 6169 7044 6193 7046
rect 5953 7024 6249 7044
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 6104 6458 6132 6802
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5953 6012 6249 6032
rect 6009 6010 6033 6012
rect 6089 6010 6113 6012
rect 6169 6010 6193 6012
rect 6031 5958 6033 6010
rect 6095 5958 6107 6010
rect 6169 5958 6171 6010
rect 6009 5956 6033 5958
rect 6089 5956 6113 5958
rect 6169 5956 6193 5958
rect 5953 5936 6249 5956
rect 5644 5222 5856 5250
rect 5448 4684 5500 4690
rect 5828 4672 5856 5222
rect 5953 4924 6249 4944
rect 6009 4922 6033 4924
rect 6089 4922 6113 4924
rect 6169 4922 6193 4924
rect 6031 4870 6033 4922
rect 6095 4870 6107 4922
rect 6169 4870 6171 4922
rect 6009 4868 6033 4870
rect 6089 4868 6113 4870
rect 6169 4868 6193 4870
rect 5953 4848 6249 4868
rect 5448 4626 5500 4632
rect 5552 4644 5856 4672
rect 5264 4616 5316 4622
rect 5170 4584 5226 4593
rect 5264 4558 5316 4564
rect 5170 4519 5226 4528
rect 5184 4486 5212 4519
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5000 4282 5028 4422
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4620 3120 4672 3126
rect 4540 3080 4620 3108
rect 4620 3062 4672 3068
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4448 2650 4476 2994
rect 4632 2922 4660 3062
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4724 2854 4752 4150
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4986 3496 5042 3505
rect 4986 3431 5042 3440
rect 5000 3126 5028 3431
rect 5092 3194 5120 3878
rect 5276 3534 5304 4558
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3738 5488 4082
rect 5552 3777 5580 4644
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5644 4214 5672 4490
rect 5828 4282 5856 4644
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5538 3768 5594 3777
rect 5448 3732 5500 3738
rect 5538 3703 5594 3712
rect 5448 3674 5500 3680
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4802 2952 4858 2961
rect 4802 2887 4858 2896
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4724 2446 4752 2586
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 3240 2372 3292 2378
rect 3068 2332 3240 2360
rect 3068 800 3096 2332
rect 3240 2314 3292 2320
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3454 2204 3750 2224
rect 3510 2202 3534 2204
rect 3590 2202 3614 2204
rect 3670 2202 3694 2204
rect 3532 2150 3534 2202
rect 3596 2150 3608 2202
rect 3670 2150 3672 2202
rect 3510 2148 3534 2150
rect 3590 2148 3614 2150
rect 3670 2148 3694 2150
rect 3454 2128 3750 2148
rect 3896 2038 3924 2246
rect 3884 2032 3936 2038
rect 3884 1974 3936 1980
rect 3516 1420 3568 1426
rect 3516 1362 3568 1368
rect 3528 800 3556 1362
rect 3988 800 4016 2246
rect 4344 1488 4396 1494
rect 4344 1430 4396 1436
rect 4356 800 4384 1430
rect 4816 800 4844 2887
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 4908 2106 4936 2518
rect 5000 2514 5028 2790
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 4986 2408 5042 2417
rect 4986 2343 5042 2352
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5000 1834 5028 2343
rect 4988 1828 5040 1834
rect 4988 1770 5040 1776
rect 5184 800 5212 3402
rect 5552 2922 5580 3703
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5644 2650 5672 3878
rect 5736 3602 5764 4014
rect 5920 3924 5948 4082
rect 6288 3942 6316 7142
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 4826 6408 5510
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6472 4554 6500 9982
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6564 6798 6592 7210
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6656 6236 6684 6870
rect 6748 6866 6776 11342
rect 6840 11286 6868 11478
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6932 10606 6960 11494
rect 7024 11478 7144 11506
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6390 6776 6802
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6840 6254 6868 9318
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6932 7478 6960 7958
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 7024 6458 7052 11290
rect 7116 10130 7144 11478
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7116 8430 7144 8842
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6828 6248 6880 6254
rect 6656 6208 6776 6236
rect 6748 6118 6776 6208
rect 6828 6190 6880 6196
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6656 5846 6684 6054
rect 6644 5840 6696 5846
rect 6748 5817 6776 6054
rect 6644 5782 6696 5788
rect 6734 5808 6790 5817
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4622 6592 4966
rect 6656 4826 6684 5782
rect 6734 5743 6790 5752
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5574 6776 5646
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5166 6776 5510
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6840 5080 6868 6190
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6932 5370 6960 5714
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6920 5092 6972 5098
rect 6840 5052 6920 5080
rect 6920 5034 6972 5040
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 5828 3896 5948 3924
rect 6276 3936 6328 3942
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5828 2990 5856 3896
rect 6276 3878 6328 3884
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 5953 3836 6249 3856
rect 6009 3834 6033 3836
rect 6089 3834 6113 3836
rect 6169 3834 6193 3836
rect 6031 3782 6033 3834
rect 6095 3782 6107 3834
rect 6169 3782 6171 3834
rect 6009 3780 6033 3782
rect 6089 3780 6113 3782
rect 6169 3780 6193 3782
rect 5953 3760 6249 3780
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6012 2990 6040 3470
rect 6288 3398 6316 3878
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5736 1442 5764 2858
rect 6288 2854 6316 3334
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 6276 2848 6328 2854
rect 6380 2825 6408 3878
rect 6472 3777 6500 4082
rect 6458 3768 6514 3777
rect 6458 3703 6514 3712
rect 6564 3670 6592 4558
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6552 2848 6604 2854
rect 6276 2790 6328 2796
rect 6366 2816 6422 2825
rect 5828 2582 5856 2790
rect 5953 2748 6249 2768
rect 6552 2790 6604 2796
rect 6366 2751 6422 2760
rect 6009 2746 6033 2748
rect 6089 2746 6113 2748
rect 6169 2746 6193 2748
rect 6031 2694 6033 2746
rect 6095 2694 6107 2746
rect 6169 2694 6171 2746
rect 6009 2692 6033 2694
rect 6089 2692 6113 2694
rect 6169 2692 6193 2694
rect 5953 2672 6249 2692
rect 6380 2650 6408 2751
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 5644 1414 5764 1442
rect 5644 800 5672 1414
rect 6012 800 6040 2314
rect 6196 1426 6224 2518
rect 6564 2446 6592 2790
rect 6656 2514 6684 4762
rect 6736 4752 6788 4758
rect 6788 4712 6868 4740
rect 6736 4694 6788 4700
rect 6840 3890 6868 4712
rect 6932 4010 6960 5034
rect 7024 4826 7052 5850
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7116 4146 7144 8026
rect 7196 7948 7248 7954
rect 7300 7936 7328 12702
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 11694 7512 12582
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7760 11354 7788 15399
rect 7852 13444 7880 17002
rect 7944 16436 7972 19200
rect 8404 17626 8432 19200
rect 8312 17598 8432 17626
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8220 17134 8248 17274
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8312 16794 8340 17598
rect 8772 17524 8800 19200
rect 8772 17496 9076 17524
rect 8452 17436 8748 17456
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8530 17382 8532 17434
rect 8594 17382 8606 17434
rect 8668 17382 8670 17434
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8452 17360 8748 17380
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8024 16448 8076 16454
rect 7944 16408 8024 16436
rect 8024 16390 8076 16396
rect 8220 16250 8248 16594
rect 8772 16561 8800 16662
rect 8864 16658 8892 16934
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8758 16552 8814 16561
rect 8758 16487 8814 16496
rect 8452 16348 8748 16368
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8530 16294 8532 16346
rect 8594 16294 8606 16346
rect 8668 16294 8670 16346
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8452 16272 8748 16292
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8206 16144 8262 16153
rect 8206 16079 8262 16088
rect 8666 16144 8722 16153
rect 8666 16079 8668 16088
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 8022 15736 8078 15745
rect 8022 15671 8024 15680
rect 8076 15671 8078 15680
rect 8024 15642 8076 15648
rect 7930 14920 7986 14929
rect 7930 14855 7986 14864
rect 7944 14822 7972 14855
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7944 14482 7972 14758
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8128 13870 8156 15914
rect 8220 15638 8248 16079
rect 8720 16079 8722 16088
rect 8668 16050 8720 16056
rect 8574 15736 8630 15745
rect 8574 15671 8576 15680
rect 8628 15671 8630 15680
rect 8576 15642 8628 15648
rect 8864 15638 8892 16594
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8956 15978 8984 16458
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 9048 15745 9076 17496
rect 9140 16726 9168 19200
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9218 16144 9274 16153
rect 9218 16079 9274 16088
rect 9232 15978 9260 16079
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9034 15736 9090 15745
rect 9034 15671 9090 15680
rect 8208 15632 8260 15638
rect 8852 15632 8904 15638
rect 8208 15574 8260 15580
rect 8758 15600 8814 15609
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8668 15564 8720 15570
rect 8852 15574 8904 15580
rect 8758 15535 8814 15544
rect 9036 15564 9088 15570
rect 8668 15506 8720 15512
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 15026 8248 15302
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8220 14414 8248 14962
rect 8312 14822 8340 15506
rect 8484 15428 8536 15434
rect 8680 15416 8708 15506
rect 8772 15434 8800 15535
rect 9036 15506 9088 15512
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8536 15388 8708 15416
rect 8760 15428 8812 15434
rect 8484 15370 8536 15376
rect 8760 15370 8812 15376
rect 8452 15260 8748 15280
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8530 15206 8532 15258
rect 8594 15206 8606 15258
rect 8668 15206 8670 15258
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8452 15184 8748 15204
rect 8864 14958 8892 15438
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8852 14952 8904 14958
rect 8956 14940 8984 15302
rect 9048 15094 9076 15506
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 9036 14952 9088 14958
rect 8956 14912 9036 14940
rect 8852 14894 8904 14900
rect 9036 14894 9088 14900
rect 8300 14816 8352 14822
rect 8760 14816 8812 14822
rect 8300 14758 8352 14764
rect 8758 14784 8760 14793
rect 8812 14784 8814 14793
rect 8758 14719 8814 14728
rect 8758 14512 8814 14521
rect 8758 14447 8760 14456
rect 8812 14447 8814 14456
rect 8944 14476 8996 14482
rect 8760 14418 8812 14424
rect 8944 14418 8996 14424
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8452 14172 8748 14192
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8530 14118 8532 14170
rect 8594 14118 8606 14170
rect 8668 14118 8670 14170
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8452 14096 8748 14116
rect 8116 13864 8168 13870
rect 8392 13864 8444 13870
rect 8116 13806 8168 13812
rect 8390 13832 8392 13841
rect 8444 13832 8446 13841
rect 8390 13767 8446 13776
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 7932 13456 7984 13462
rect 7852 13416 7932 13444
rect 7932 13398 7984 13404
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12714 7972 13126
rect 8220 12850 8248 13670
rect 8452 13084 8748 13104
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8530 13030 8532 13082
rect 8594 13030 8606 13082
rect 8668 13030 8670 13082
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8452 13008 8748 13028
rect 8864 12986 8892 14350
rect 8956 13870 8984 14418
rect 9048 14278 9076 14894
rect 9140 14890 9168 15914
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9126 14512 9182 14521
rect 9126 14447 9128 14456
rect 9180 14447 9182 14456
rect 9128 14418 9180 14424
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13870 9076 14214
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8956 13530 8984 13806
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8944 13184 8996 13190
rect 9048 13172 9076 13670
rect 9232 13410 9260 15914
rect 9416 15910 9444 16526
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9402 15736 9458 15745
rect 9402 15671 9458 15680
rect 9416 15162 9444 15671
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9416 14958 9444 15098
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14482 9352 14758
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9324 13841 9352 14418
rect 9416 14346 9444 14554
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9310 13832 9366 13841
rect 9310 13767 9366 13776
rect 9128 13388 9180 13394
rect 9232 13382 9352 13410
rect 9128 13330 9180 13336
rect 9140 13190 9168 13330
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8996 13144 9076 13172
rect 9128 13184 9180 13190
rect 8944 13126 8996 13132
rect 9128 13126 9180 13132
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 11898 7972 12650
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8852 12640 8904 12646
rect 8956 12628 8984 13126
rect 9140 12850 9168 13126
rect 9232 13025 9260 13262
rect 9218 13016 9274 13025
rect 9218 12951 9274 12960
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8904 12600 8984 12628
rect 8852 12582 8904 12588
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8036 11762 8064 12582
rect 8452 11996 8748 12016
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8530 11942 8532 11994
rect 8594 11942 8606 11994
rect 8668 11942 8670 11994
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8452 11920 8748 11940
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7576 10674 7604 11154
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7668 10606 7696 10950
rect 7656 10600 7708 10606
rect 7840 10600 7892 10606
rect 7656 10542 7708 10548
rect 7838 10568 7840 10577
rect 7892 10568 7894 10577
rect 7838 10503 7894 10512
rect 7932 10464 7984 10470
rect 8036 10452 8064 10950
rect 7984 10424 8064 10452
rect 7932 10406 7984 10412
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8090 7420 8774
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7484 7970 7512 8230
rect 7248 7908 7328 7936
rect 7392 7942 7512 7970
rect 7196 7890 7248 7896
rect 7208 7857 7236 7890
rect 7392 7886 7420 7942
rect 7380 7880 7432 7886
rect 7194 7848 7250 7857
rect 7576 7834 7604 9862
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7668 9042 7696 9658
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7380 7822 7432 7828
rect 7194 7783 7250 7792
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5166 7236 6258
rect 7300 6186 7328 7142
rect 7392 6934 7420 7822
rect 7484 7806 7604 7834
rect 7484 7478 7512 7806
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7484 6866 7512 7278
rect 7576 6934 7604 7686
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 7002 7696 7142
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5914 7420 6054
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7840 5840 7892 5846
rect 7378 5808 7434 5817
rect 7840 5782 7892 5788
rect 7378 5743 7434 5752
rect 7472 5772 7524 5778
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7300 4282 7328 4694
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6840 3862 6960 3890
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6748 1494 6776 2518
rect 6736 1488 6788 1494
rect 6736 1430 6788 1436
rect 6184 1420 6236 1426
rect 6184 1362 6236 1368
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 6472 800 6500 1362
rect 6840 800 6868 3674
rect 6932 2514 6960 3862
rect 7300 2514 7328 4218
rect 7392 4049 7420 5743
rect 7472 5714 7524 5720
rect 7484 5234 7512 5714
rect 7852 5302 7880 5782
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4622 7512 5170
rect 7748 5160 7800 5166
rect 7746 5128 7748 5137
rect 7800 5128 7802 5137
rect 7746 5063 7802 5072
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4826 7788 4966
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7562 4176 7618 4185
rect 7472 4140 7524 4146
rect 7562 4111 7618 4120
rect 7472 4082 7524 4088
rect 7378 4040 7434 4049
rect 7378 3975 7434 3984
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 2990 7420 3334
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7288 2508 7340 2514
rect 7484 2496 7512 4082
rect 7576 4010 7604 4111
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7576 3602 7604 3946
rect 7668 3942 7696 4626
rect 7760 4593 7788 4626
rect 7746 4584 7802 4593
rect 7746 4519 7802 4528
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4146 7880 4422
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7944 4078 7972 10066
rect 8128 9926 8156 11630
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8452 10908 8748 10928
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8530 10854 8532 10906
rect 8594 10854 8606 10906
rect 8668 10854 8670 10906
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8452 10832 8748 10852
rect 8758 10568 8814 10577
rect 8758 10503 8760 10512
rect 8812 10503 8814 10512
rect 8760 10474 8812 10480
rect 8864 10266 8892 11154
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8220 6882 8248 9930
rect 8452 9820 8748 9840
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8530 9766 8532 9818
rect 8594 9766 8606 9818
rect 8668 9766 8670 9818
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8452 9744 8748 9764
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8312 7886 8340 9522
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8588 9178 8616 9318
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8452 8732 8748 8752
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8530 8678 8532 8730
rect 8594 8678 8606 8730
rect 8668 8678 8670 8730
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8452 8656 8748 8676
rect 8482 8528 8538 8537
rect 8482 8463 8538 8472
rect 8496 8294 8524 8463
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8404 8090 8432 8230
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8666 7984 8722 7993
rect 8772 7970 8800 8230
rect 8864 8090 8892 9386
rect 8956 8809 8984 12600
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9048 11286 9076 12310
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9048 10674 9076 11222
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9140 9654 9168 11494
rect 9232 10742 9260 11698
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9324 9654 9352 13382
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 8942 8800 8998 8809
rect 8942 8735 8998 8744
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8772 7942 8892 7970
rect 8666 7919 8722 7928
rect 8680 7886 8708 7919
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8312 7342 8340 7822
rect 8452 7644 8748 7664
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8530 7590 8532 7642
rect 8594 7590 8606 7642
rect 8668 7590 8670 7642
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8452 7568 8748 7588
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 7002 8340 7278
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8220 6854 8340 6882
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8036 5370 8064 6394
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5642 8156 6190
rect 8312 5778 8340 6854
rect 8588 6730 8616 7414
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 6934 8708 7278
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8772 6730 8800 7210
rect 8864 7177 8892 7942
rect 8956 7546 8984 8570
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8942 7440 8998 7449
rect 8942 7375 8998 7384
rect 8850 7168 8906 7177
rect 8850 7103 8906 7112
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8452 6556 8748 6576
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8530 6502 8532 6554
rect 8594 6502 8606 6554
rect 8668 6502 8670 6554
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8452 6480 8748 6500
rect 8864 6254 8892 6870
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8036 4758 8064 5306
rect 8128 5302 8156 5578
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8128 4468 8156 5238
rect 8036 4440 8156 4468
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7656 2508 7708 2514
rect 7484 2468 7656 2496
rect 7288 2450 7340 2456
rect 7656 2450 7708 2456
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7300 800 7328 2246
rect 7668 2106 7696 2450
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7760 800 7788 3878
rect 8036 3602 8064 4440
rect 8220 4146 8248 5510
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8312 4078 8340 5510
rect 8452 5468 8748 5488
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8530 5414 8532 5466
rect 8594 5414 8606 5466
rect 8668 5414 8670 5466
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8452 5392 8748 5412
rect 8484 5160 8536 5166
rect 8482 5128 8484 5137
rect 8536 5128 8538 5137
rect 8482 5063 8538 5072
rect 8864 4690 8892 5646
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8956 4622 8984 7375
rect 9048 7274 9076 9522
rect 9128 9512 9180 9518
rect 9232 9489 9260 9590
rect 9128 9454 9180 9460
rect 9218 9480 9274 9489
rect 9140 9178 9168 9454
rect 9218 9415 9274 9424
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9140 9081 9168 9114
rect 9126 9072 9182 9081
rect 9126 9007 9182 9016
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9140 8498 9168 8910
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9232 8498 9260 8774
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9232 8378 9260 8434
rect 9416 8430 9444 14282
rect 9508 12102 9536 16662
rect 9600 15722 9628 19200
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9692 15978 9720 18090
rect 9968 17320 9996 19200
rect 9784 17292 10364 17320
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9600 15694 9720 15722
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9600 15366 9628 15574
rect 9588 15360 9640 15366
rect 9692 15337 9720 15694
rect 9588 15302 9640 15308
rect 9678 15328 9734 15337
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11830 9536 12038
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9508 11558 9536 11766
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9140 8350 9260 8378
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9140 7585 9168 8350
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 8090 9260 8230
rect 9508 8090 9536 10610
rect 9600 9042 9628 15302
rect 9784 15314 9812 17292
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9876 16658 9904 16934
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9876 15638 9904 16594
rect 9954 16552 10010 16561
rect 9954 16487 10010 16496
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9784 15286 9904 15314
rect 9678 15263 9734 15272
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9692 14346 9720 15098
rect 9784 15026 9812 15098
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9692 13938 9720 14282
rect 9784 14074 9812 14962
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9692 12238 9720 13398
rect 9876 13161 9904 15286
rect 9862 13152 9918 13161
rect 9862 13087 9918 13096
rect 9968 12986 9996 16487
rect 10060 16250 10088 16934
rect 10152 16794 10180 17138
rect 10336 16794 10364 17292
rect 10140 16788 10192 16794
rect 10324 16788 10376 16794
rect 10192 16748 10272 16776
rect 10140 16730 10192 16736
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10152 16114 10180 16390
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10244 15994 10272 16748
rect 10324 16730 10376 16736
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10152 15966 10272 15994
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 10060 13433 10088 15370
rect 10152 14906 10180 15966
rect 10232 15904 10284 15910
rect 10336 15892 10364 16390
rect 10428 16250 10456 19200
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10416 15904 10468 15910
rect 10336 15864 10416 15892
rect 10232 15846 10284 15852
rect 10416 15846 10468 15852
rect 10244 15638 10272 15846
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10428 15434 10456 15846
rect 10520 15706 10548 16934
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10152 14878 10272 14906
rect 10140 14816 10192 14822
rect 10138 14784 10140 14793
rect 10192 14784 10194 14793
rect 10138 14719 10194 14728
rect 10152 14006 10180 14719
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10046 13424 10102 13433
rect 10046 13359 10102 13368
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9954 12744 10010 12753
rect 9954 12679 10010 12688
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11898 9720 12038
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9876 11830 9904 12582
rect 9968 12374 9996 12679
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9864 11824 9916 11830
rect 9968 11801 9996 12174
rect 9864 11766 9916 11772
rect 9954 11792 10010 11801
rect 9954 11727 10010 11736
rect 10060 11694 10088 13359
rect 10244 13240 10272 14878
rect 10152 13212 10272 13240
rect 10152 12102 10180 13212
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10336 11880 10364 15302
rect 10612 15162 10640 17138
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15706 10732 15846
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10796 15366 10824 19200
rect 11256 17202 11284 19200
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 10950 16892 11246 16912
rect 11006 16890 11030 16892
rect 11086 16890 11110 16892
rect 11166 16890 11190 16892
rect 11028 16838 11030 16890
rect 11092 16838 11104 16890
rect 11166 16838 11168 16890
rect 11006 16836 11030 16838
rect 11086 16836 11110 16838
rect 11166 16836 11190 16838
rect 10950 16816 11246 16836
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11164 15978 11192 16662
rect 11256 16114 11284 16662
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 10950 15804 11246 15824
rect 11006 15802 11030 15804
rect 11086 15802 11110 15804
rect 11166 15802 11190 15804
rect 11028 15750 11030 15802
rect 11092 15750 11104 15802
rect 11166 15750 11168 15802
rect 11006 15748 11030 15750
rect 11086 15748 11110 15750
rect 11166 15748 11190 15750
rect 10950 15728 11246 15748
rect 11348 15706 11376 16934
rect 11440 16794 11468 17138
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11440 15502 11468 16730
rect 11624 16402 11652 19200
rect 11624 16374 12020 16402
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11532 15502 11560 16050
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10428 14482 10456 15098
rect 10612 14550 10640 15098
rect 10782 15056 10838 15065
rect 10782 14991 10838 15000
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10520 12986 10548 14486
rect 10796 13734 10824 14991
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10428 12646 10456 12922
rect 10612 12866 10640 13330
rect 10520 12850 10824 12866
rect 10508 12844 10836 12850
rect 10560 12838 10784 12844
rect 10508 12786 10560 12792
rect 10784 12786 10836 12792
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10416 12640 10468 12646
rect 10468 12600 10548 12628
rect 10416 12582 10468 12588
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10152 11852 10364 11880
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 9178 9720 11562
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9784 11150 9812 11290
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10470 9812 10950
rect 9876 10606 9904 11494
rect 10152 11234 10180 11852
rect 10428 11762 10456 12038
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 9968 11206 10180 11234
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 9586 9812 10406
rect 9876 10130 9904 10542
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9968 10010 9996 11206
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9876 9982 9996 10010
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9784 8974 9812 9522
rect 9876 9194 9904 9982
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 9518 9996 9862
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9956 9376 10008 9382
rect 9954 9344 9956 9353
rect 10008 9344 10010 9353
rect 9954 9279 10010 9288
rect 9876 9166 9996 9194
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9600 8401 9628 8570
rect 9586 8392 9642 8401
rect 9586 8327 9642 8336
rect 9588 8288 9640 8294
rect 9586 8256 9588 8265
rect 9640 8256 9642 8265
rect 9586 8191 9642 8200
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9218 7984 9274 7993
rect 9218 7919 9274 7928
rect 9496 7948 9548 7954
rect 9126 7576 9182 7585
rect 9126 7511 9182 7520
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9034 7168 9090 7177
rect 9140 7154 9168 7414
rect 9232 7290 9260 7919
rect 9496 7890 9548 7896
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9324 7410 9352 7754
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9232 7262 9352 7290
rect 9140 7126 9260 7154
rect 9034 7103 9090 7112
rect 9048 5846 9076 7103
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 9140 4826 9168 6870
rect 9232 6798 9260 7126
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6662 9260 6734
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8452 4380 8748 4400
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8530 4326 8532 4378
rect 8594 4326 8606 4378
rect 8668 4326 8670 4378
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8452 4304 8748 4324
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 2514 7972 3334
rect 8036 3058 8064 3538
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7852 1426 7880 2246
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 8128 800 8156 3946
rect 8404 3380 8432 4150
rect 8312 3352 8432 3380
rect 8312 3108 8340 3352
rect 8452 3292 8748 3312
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8530 3238 8532 3290
rect 8594 3238 8606 3290
rect 8668 3238 8670 3290
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8452 3216 8748 3236
rect 8864 3194 8892 4490
rect 9140 4434 9168 4762
rect 9232 4554 9260 6598
rect 9324 5574 9352 7262
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9140 4406 9260 4434
rect 8942 4312 8998 4321
rect 8942 4247 8998 4256
rect 8956 3398 8984 4247
rect 9126 4176 9182 4185
rect 9126 4111 9182 4120
rect 9140 4010 9168 4111
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 9232 3924 9260 4406
rect 9324 4146 9352 5510
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9416 4622 9444 5034
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9312 3936 9364 3942
rect 9232 3896 9312 3924
rect 9312 3878 9364 3884
rect 9126 3768 9182 3777
rect 9126 3703 9182 3712
rect 9140 3466 9168 3703
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8852 3188 8904 3194
rect 8772 3148 8852 3176
rect 8312 3080 8432 3108
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8312 2650 8340 2926
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2514 8432 3080
rect 8392 2508 8444 2514
rect 8772 2496 8800 3148
rect 8852 3130 8904 3136
rect 8850 3088 8906 3097
rect 9324 3074 9352 3878
rect 9416 3738 9444 4558
rect 9508 4214 9536 7890
rect 9586 7848 9642 7857
rect 9586 7783 9642 7792
rect 9600 7750 9628 7783
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 6934 9628 7686
rect 9692 7206 9720 8842
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8430 9812 8774
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9784 8090 9812 8366
rect 9876 8294 9904 9046
rect 9968 8906 9996 9166
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9692 6458 9720 6870
rect 9784 6866 9812 8026
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9876 7206 9904 7482
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9876 6662 9904 7142
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5846 9720 6054
rect 9876 5846 9904 6598
rect 9968 6458 9996 8026
rect 10060 6905 10088 11086
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10152 9178 10180 11018
rect 10244 9994 10272 11698
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 10152 7886 10180 9007
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10046 6896 10102 6905
rect 10046 6831 10102 6840
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 5370 9628 5646
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9586 5264 9642 5273
rect 9586 5199 9642 5208
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9416 3194 9444 3538
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9324 3046 9444 3074
rect 8850 3023 8906 3032
rect 8864 2650 8892 3023
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8772 2468 8984 2496
rect 8392 2450 8444 2456
rect 8452 2204 8748 2224
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8530 2150 8532 2202
rect 8594 2150 8606 2202
rect 8668 2150 8670 2202
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8452 2128 8748 2148
rect 8576 1148 8628 1154
rect 8576 1090 8628 1096
rect 8588 800 8616 1090
rect 8956 800 8984 2468
rect 9140 1154 9168 2790
rect 9416 2310 9444 3046
rect 9508 2650 9536 3878
rect 9600 3466 9628 5199
rect 9692 4078 9720 5782
rect 9876 4758 9904 5782
rect 9968 5778 9996 6394
rect 10060 6118 10088 6831
rect 10152 6458 10180 7822
rect 10244 7342 10272 9930
rect 10336 7546 10364 10066
rect 10428 8634 10456 11290
rect 10520 9466 10548 12600
rect 10612 11898 10640 12718
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 12442 10732 12582
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10598 11792 10654 11801
rect 10598 11727 10654 11736
rect 10612 9897 10640 11727
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10704 10538 10732 11086
rect 10796 11082 10824 11630
rect 10888 11286 10916 15370
rect 11072 14958 11100 15438
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10950 14716 11246 14736
rect 11006 14714 11030 14716
rect 11086 14714 11110 14716
rect 11166 14714 11190 14716
rect 11028 14662 11030 14714
rect 11092 14662 11104 14714
rect 11166 14662 11168 14714
rect 11006 14660 11030 14662
rect 11086 14660 11110 14662
rect 11166 14660 11190 14662
rect 10950 14640 11246 14660
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11256 13716 11284 14418
rect 11348 14074 11376 14962
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11532 13977 11560 14010
rect 11518 13968 11574 13977
rect 11518 13903 11574 13912
rect 11256 13688 11376 13716
rect 10950 13628 11246 13648
rect 11006 13626 11030 13628
rect 11086 13626 11110 13628
rect 11166 13626 11190 13628
rect 11028 13574 11030 13626
rect 11092 13574 11104 13626
rect 11166 13574 11168 13626
rect 11006 13572 11030 13574
rect 11086 13572 11110 13574
rect 11166 13572 11190 13574
rect 10950 13552 11246 13572
rect 11348 13462 11376 13688
rect 11624 13682 11652 16186
rect 11794 16008 11850 16017
rect 11900 15960 11928 16186
rect 11850 15952 11928 15960
rect 11794 15943 11796 15952
rect 11848 15932 11928 15952
rect 11796 15914 11848 15920
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11532 13654 11652 13682
rect 11532 13462 11560 13654
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11336 13456 11388 13462
rect 11520 13456 11572 13462
rect 11336 13398 11388 13404
rect 11518 13424 11520 13433
rect 11572 13424 11574 13433
rect 10950 12540 11246 12560
rect 11006 12538 11030 12540
rect 11086 12538 11110 12540
rect 11166 12538 11190 12540
rect 11028 12486 11030 12538
rect 11092 12486 11104 12538
rect 11166 12486 11168 12538
rect 11006 12484 11030 12486
rect 11086 12484 11110 12486
rect 11166 12484 11190 12486
rect 10950 12464 11246 12484
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10980 11762 11008 12242
rect 11348 12102 11376 13398
rect 11518 13359 11574 13368
rect 11520 13320 11572 13326
rect 11518 13288 11520 13297
rect 11572 13288 11574 13297
rect 11518 13223 11574 13232
rect 11426 13152 11482 13161
rect 11426 13087 11482 13096
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11348 11558 11376 12038
rect 11440 11898 11468 13087
rect 11532 12889 11560 13223
rect 11518 12880 11574 12889
rect 11624 12850 11652 13466
rect 11716 13190 11744 14894
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11518 12815 11574 12824
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11440 11694 11468 11834
rect 11716 11694 11744 13126
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10950 11452 11246 11472
rect 11006 11450 11030 11452
rect 11086 11450 11110 11452
rect 11166 11450 11190 11452
rect 11028 11398 11030 11450
rect 11092 11398 11104 11450
rect 11166 11398 11168 11450
rect 11006 11396 11030 11398
rect 11086 11396 11110 11398
rect 11166 11396 11190 11398
rect 10950 11376 11246 11396
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 11348 11218 11376 11494
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10704 9926 10732 10474
rect 10692 9920 10744 9926
rect 10598 9888 10654 9897
rect 10692 9862 10744 9868
rect 10598 9823 10654 9832
rect 10704 9586 10732 9862
rect 10796 9654 10824 11018
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10888 9518 10916 11086
rect 11348 10606 11376 11154
rect 11440 11150 11468 11630
rect 11518 11384 11574 11393
rect 11518 11319 11520 11328
rect 11572 11319 11574 11328
rect 11520 11290 11572 11296
rect 11518 11248 11574 11257
rect 11518 11183 11574 11192
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 10950 10364 11246 10384
rect 11006 10362 11030 10364
rect 11086 10362 11110 10364
rect 11166 10362 11190 10364
rect 11028 10310 11030 10362
rect 11092 10310 11104 10362
rect 11166 10310 11168 10362
rect 11006 10308 11030 10310
rect 11086 10308 11110 10310
rect 11166 10308 11190 10310
rect 10950 10288 11246 10308
rect 11348 10062 11376 10542
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 10876 9512 10928 9518
rect 10520 9438 10732 9466
rect 10876 9454 10928 9460
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9194 10548 9318
rect 10520 9166 10640 9194
rect 10704 9178 10732 9438
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10336 6934 10364 7346
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10428 6458 10456 7890
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7546 10548 7822
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10612 7188 10640 9166
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10888 9081 10916 9454
rect 10950 9276 11246 9296
rect 11006 9274 11030 9276
rect 11086 9274 11110 9276
rect 11166 9274 11190 9276
rect 11028 9222 11030 9274
rect 11092 9222 11104 9274
rect 11166 9222 11168 9274
rect 11006 9220 11030 9222
rect 11086 9220 11110 9222
rect 11166 9220 11190 9222
rect 10950 9200 11246 9220
rect 11152 9104 11204 9110
rect 10874 9072 10930 9081
rect 11152 9046 11204 9052
rect 10874 9007 10930 9016
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10704 8838 10732 8910
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8634 10732 8774
rect 11164 8634 11192 9046
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10704 7886 10732 8298
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 7478 10732 7822
rect 10888 7818 10916 8230
rect 10950 8188 11246 8208
rect 11006 8186 11030 8188
rect 11086 8186 11110 8188
rect 11166 8186 11190 8188
rect 11028 8134 11030 8186
rect 11092 8134 11104 8186
rect 11166 8134 11168 8186
rect 11006 8132 11030 8134
rect 11086 8132 11110 8134
rect 11166 8132 11190 8134
rect 10950 8112 11246 8132
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 11256 7546 11284 7890
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10692 7200 10744 7206
rect 10612 7160 10692 7188
rect 10692 7142 10744 7148
rect 10704 7002 10732 7142
rect 10888 7002 10916 7346
rect 10950 7100 11246 7120
rect 11006 7098 11030 7100
rect 11086 7098 11110 7100
rect 11166 7098 11190 7100
rect 11028 7046 11030 7098
rect 11092 7046 11104 7098
rect 11166 7046 11168 7098
rect 11006 7044 11030 7046
rect 11086 7044 11110 7046
rect 11166 7044 11190 7046
rect 10950 7024 11246 7044
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10152 6118 10180 6394
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4282 9812 4626
rect 10046 4584 10102 4593
rect 10046 4519 10102 4528
rect 9864 4480 9916 4486
rect 9916 4440 9996 4468
rect 9864 4422 9916 4428
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9692 3369 9720 3470
rect 9678 3360 9734 3369
rect 9678 3295 9734 3304
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9600 2446 9628 3130
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9692 2922 9720 2994
rect 9784 2990 9812 4082
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9770 2816 9826 2825
rect 9770 2751 9826 2760
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9128 1148 9180 1154
rect 9128 1090 9180 1096
rect 9416 800 9444 2246
rect 9784 800 9812 2751
rect 9876 2650 9904 3878
rect 9968 3233 9996 4440
rect 10060 4010 10088 4519
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10152 3890 10180 4150
rect 10060 3862 10180 3890
rect 9954 3224 10010 3233
rect 9954 3159 10010 3168
rect 9968 2854 9996 3159
rect 9956 2848 10008 2854
rect 10060 2825 10088 3862
rect 10244 3534 10272 4966
rect 10428 4826 10456 4966
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10520 4622 10548 5034
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10612 4457 10640 6326
rect 10888 6322 10916 6938
rect 11348 6798 11376 8502
rect 11440 7886 11468 8570
rect 11532 8514 11560 11183
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 11532 8486 11652 8514
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10704 5846 10732 6054
rect 10950 6012 11246 6032
rect 11006 6010 11030 6012
rect 11086 6010 11110 6012
rect 11166 6010 11190 6012
rect 11028 5958 11030 6010
rect 11092 5958 11104 6010
rect 11166 5958 11168 6010
rect 11006 5956 11030 5958
rect 11086 5956 11110 5958
rect 11166 5956 11190 5958
rect 10950 5936 11246 5956
rect 10692 5840 10744 5846
rect 10744 5800 10916 5828
rect 10692 5782 10744 5788
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10704 5098 10732 5170
rect 10796 5166 10824 5578
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10598 4448 10654 4457
rect 10598 4383 10654 4392
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10322 3904 10378 3913
rect 10322 3839 10378 3848
rect 10232 3528 10284 3534
rect 10138 3496 10194 3505
rect 10232 3470 10284 3476
rect 10138 3431 10194 3440
rect 10152 3194 10180 3431
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10244 3097 10272 3470
rect 10336 3398 10364 3839
rect 10428 3618 10456 4218
rect 10612 3942 10640 4383
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10520 3738 10548 3878
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10428 3590 10548 3618
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10416 3392 10468 3398
rect 10520 3369 10548 3590
rect 10416 3334 10468 3340
rect 10506 3360 10562 3369
rect 10230 3088 10286 3097
rect 10230 3023 10286 3032
rect 9956 2790 10008 2796
rect 10046 2816 10102 2825
rect 10046 2751 10102 2760
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10244 800 10272 3023
rect 10336 1562 10364 3334
rect 10428 2582 10456 3334
rect 10506 3295 10562 3304
rect 10612 2836 10640 3878
rect 10704 3534 10732 5034
rect 10796 4758 10824 5102
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10888 4690 10916 5800
rect 10950 4924 11246 4944
rect 11006 4922 11030 4924
rect 11086 4922 11110 4924
rect 11166 4922 11190 4924
rect 11028 4870 11030 4922
rect 11092 4870 11104 4922
rect 11166 4870 11168 4922
rect 11006 4868 11030 4870
rect 11086 4868 11110 4870
rect 11166 4868 11190 4870
rect 10950 4848 11246 4868
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 11152 4616 11204 4622
rect 11348 4604 11376 6598
rect 11532 5914 11560 8366
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11204 4576 11376 4604
rect 11152 4558 11204 4564
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10796 3602 10824 4218
rect 10980 4146 11008 4490
rect 11164 4214 11192 4558
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11336 4072 11388 4078
rect 10874 4040 10930 4049
rect 11336 4014 11388 4020
rect 10874 3975 10876 3984
rect 10928 3975 10930 3984
rect 10876 3946 10928 3952
rect 10950 3836 11246 3856
rect 11006 3834 11030 3836
rect 11086 3834 11110 3836
rect 11166 3834 11190 3836
rect 11028 3782 11030 3834
rect 11092 3782 11104 3834
rect 11166 3782 11168 3834
rect 11006 3780 11030 3782
rect 11086 3780 11110 3782
rect 11166 3780 11190 3782
rect 10950 3760 11246 3780
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10704 2990 10732 3470
rect 10692 2984 10744 2990
rect 10744 2944 10824 2972
rect 10692 2926 10744 2932
rect 10612 2808 10732 2836
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10324 1556 10376 1562
rect 10324 1498 10376 1504
rect 10704 800 10732 2808
rect 10796 2446 10824 2944
rect 10888 2854 10916 3470
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10950 2748 11246 2768
rect 11006 2746 11030 2748
rect 11086 2746 11110 2748
rect 11166 2746 11190 2748
rect 11028 2694 11030 2746
rect 11092 2694 11104 2746
rect 11166 2694 11168 2746
rect 11006 2692 11030 2694
rect 11086 2692 11110 2694
rect 11166 2692 11190 2694
rect 10950 2672 11246 2692
rect 11348 2650 11376 4014
rect 11440 3738 11468 5306
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11532 3618 11560 5646
rect 11624 3641 11652 8486
rect 11716 8344 11744 9415
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11808 8498 11836 8910
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11796 8356 11848 8362
rect 11716 8316 11796 8344
rect 11796 8298 11848 8304
rect 11702 7984 11758 7993
rect 11702 7919 11704 7928
rect 11756 7919 11758 7928
rect 11704 7890 11756 7896
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11716 5098 11744 5306
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11716 4622 11744 5034
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11808 4026 11836 8298
rect 11900 6118 11928 15932
rect 11992 12374 12020 16374
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 12084 11558 12112 19200
rect 12452 17241 12480 19200
rect 12912 18154 12940 19200
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 12900 18012 12952 18018
rect 12900 17954 12952 17960
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12438 17232 12494 17241
rect 12438 17167 12494 17176
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 16250 12480 17002
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12176 15638 12204 15982
rect 12544 15706 12572 17614
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12636 16794 12664 17206
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 12162 15464 12218 15473
rect 12162 15399 12164 15408
rect 12216 15399 12218 15408
rect 12164 15370 12216 15376
rect 12256 14952 12308 14958
rect 12162 14920 12218 14929
rect 12256 14894 12308 14900
rect 12162 14855 12164 14864
rect 12216 14855 12218 14864
rect 12164 14826 12216 14832
rect 12176 14550 12204 14826
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 13802 12204 13874
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11992 9722 12020 10406
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 12084 9654 12112 11222
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12084 9024 12112 9590
rect 12176 9178 12204 13738
rect 12268 13258 12296 14894
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12360 13002 12388 13670
rect 12544 13433 12572 15642
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12530 13424 12586 13433
rect 12530 13359 12586 13368
rect 12532 13320 12584 13326
rect 12530 13288 12532 13297
rect 12584 13288 12586 13297
rect 12530 13223 12586 13232
rect 12360 12974 12480 13002
rect 12452 12918 12480 12974
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12360 12442 12388 12786
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12268 11801 12296 12038
rect 12254 11792 12310 11801
rect 12360 11762 12388 12378
rect 12452 11898 12480 12718
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12254 11727 12310 11736
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12268 10810 12296 11154
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12268 9722 12296 10746
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12176 9042 12204 9114
rect 11992 8996 12112 9024
rect 12164 9036 12216 9042
rect 11992 6474 12020 8996
rect 12164 8978 12216 8984
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12084 8498 12112 8842
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12360 8430 12388 11494
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10470 12480 10950
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 8022 12296 8230
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 6662 12112 7346
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11992 6446 12388 6474
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 4146 11928 6054
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12176 4214 12204 4422
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12268 4146 12296 4694
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 11808 3998 11928 4026
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11716 3738 11744 3878
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11440 3590 11560 3618
rect 11610 3632 11666 3641
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 10968 2508 11020 2514
rect 11440 2496 11468 3590
rect 11610 3567 11666 3576
rect 11624 2990 11652 3567
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 10968 2450 11020 2456
rect 11072 2468 11468 2496
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10980 2106 11008 2450
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11072 800 11100 2468
rect 11716 2446 11744 2518
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 11532 800 11560 1498
rect 11900 800 11928 3998
rect 12268 3670 12296 4082
rect 12072 3664 12124 3670
rect 12070 3632 12072 3641
rect 12256 3664 12308 3670
rect 12124 3632 12126 3641
rect 12256 3606 12308 3612
rect 12070 3567 12126 3576
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12084 3194 12112 3470
rect 12256 3392 12308 3398
rect 12254 3360 12256 3369
rect 12308 3360 12310 3369
rect 12254 3295 12310 3304
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11978 3088 12034 3097
rect 11978 3023 11980 3032
rect 12032 3023 12034 3032
rect 11980 2994 12032 3000
rect 12256 2984 12308 2990
rect 12070 2952 12126 2961
rect 12256 2926 12308 2932
rect 12070 2887 12126 2896
rect 12084 2650 12112 2887
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12176 2496 12204 2586
rect 12084 2468 12204 2496
rect 12084 2038 12112 2468
rect 12164 2372 12216 2378
rect 12268 2360 12296 2926
rect 12216 2332 12296 2360
rect 12164 2314 12216 2320
rect 12072 2032 12124 2038
rect 12072 1974 12124 1980
rect 12360 800 12388 6446
rect 12544 3720 12572 12650
rect 12636 12646 12664 15438
rect 12728 15366 12756 15846
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12820 14906 12848 17274
rect 12912 16182 12940 17954
rect 13280 17678 13308 19200
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13648 17610 13676 19200
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12728 14878 12848 14906
rect 12728 14362 12756 14878
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12820 14618 12848 14758
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12728 14334 12848 14362
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12728 13530 12756 14214
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12714 13424 12770 13433
rect 12714 13359 12770 13368
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12636 11694 12664 12174
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10674 12664 10950
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10198 12664 10610
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 7954 12664 9998
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12728 7410 12756 13359
rect 12820 12714 12848 14334
rect 12912 13258 12940 14758
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 13004 13172 13032 17546
rect 13449 17436 13745 17456
rect 13505 17434 13529 17436
rect 13585 17434 13609 17436
rect 13665 17434 13689 17436
rect 13527 17382 13529 17434
rect 13591 17382 13603 17434
rect 13665 17382 13667 17434
rect 13505 17380 13529 17382
rect 13585 17380 13609 17382
rect 13665 17380 13689 17382
rect 13449 17360 13745 17380
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16522 13124 16934
rect 13176 16720 13228 16726
rect 13176 16662 13228 16668
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 13096 15638 13124 16458
rect 13188 16250 13216 16662
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13096 14804 13124 15574
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13188 14958 13216 15506
rect 13280 15162 13308 16594
rect 13372 16114 13400 17002
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 16726 14044 16934
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13449 16348 13745 16368
rect 13505 16346 13529 16348
rect 13585 16346 13609 16348
rect 13665 16346 13689 16348
rect 13527 16294 13529 16346
rect 13591 16294 13603 16346
rect 13665 16294 13667 16346
rect 13505 16292 13529 16294
rect 13585 16292 13609 16294
rect 13665 16292 13689 16294
rect 13449 16272 13745 16292
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13372 15026 13400 16050
rect 13740 15570 13768 16050
rect 14108 15994 14136 19200
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14016 15966 14136 15994
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13449 15260 13745 15280
rect 13505 15258 13529 15260
rect 13585 15258 13609 15260
rect 13665 15258 13689 15260
rect 13527 15206 13529 15258
rect 13591 15206 13603 15258
rect 13665 15206 13667 15258
rect 13505 15204 13529 15206
rect 13585 15204 13609 15206
rect 13665 15204 13689 15206
rect 13449 15184 13745 15204
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13096 14776 13308 14804
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 13938 13124 14282
rect 13188 14006 13216 14418
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13096 13326 13124 13874
rect 13280 13870 13308 14776
rect 13449 14172 13745 14192
rect 13505 14170 13529 14172
rect 13585 14170 13609 14172
rect 13665 14170 13689 14172
rect 13527 14118 13529 14170
rect 13591 14118 13603 14170
rect 13665 14118 13667 14170
rect 13505 14116 13529 14118
rect 13585 14116 13609 14118
rect 13665 14116 13689 14118
rect 13449 14096 13745 14116
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13372 13530 13400 13670
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13740 13326 13768 13738
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13004 13144 13124 13172
rect 12900 12776 12952 12782
rect 12898 12744 12900 12753
rect 12952 12744 12954 12753
rect 12808 12708 12860 12714
rect 12898 12679 12954 12688
rect 12808 12650 12860 12656
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 9654 12848 10474
rect 12912 10470 12940 12582
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12912 9466 12940 10406
rect 13004 9994 13032 10474
rect 13096 10266 13124 13144
rect 13449 13084 13745 13104
rect 13505 13082 13529 13084
rect 13585 13082 13609 13084
rect 13665 13082 13689 13084
rect 13527 13030 13529 13082
rect 13591 13030 13603 13082
rect 13665 13030 13667 13082
rect 13505 13028 13529 13030
rect 13585 13028 13609 13030
rect 13665 13028 13689 13030
rect 13449 13008 13745 13028
rect 14016 12986 14044 15966
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14108 15706 14136 15846
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14108 15065 14136 15438
rect 14200 15162 14228 15846
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14094 15056 14150 15065
rect 14094 14991 14150 15000
rect 14292 14822 14320 18090
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17338 14412 17478
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14476 15366 14504 19200
rect 14936 17218 14964 19200
rect 14660 17190 14964 17218
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14660 15094 14688 17190
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 15978 14780 16934
rect 14936 16454 14964 17070
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14384 14074 14412 14350
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13004 9586 13032 9930
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13084 9512 13136 9518
rect 12808 9444 12860 9450
rect 12912 9438 13032 9466
rect 13084 9454 13136 9460
rect 12808 9386 12860 9392
rect 12820 8090 12848 9386
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9178 12940 9318
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12820 7290 12848 7890
rect 13004 7698 13032 9438
rect 13096 9178 13124 9454
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13188 9058 13216 12854
rect 14016 12782 14044 12922
rect 14476 12918 14504 14826
rect 14752 13870 14780 15914
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14844 15502 14872 15642
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 15026 14872 15302
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14844 14006 14872 14962
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 10130 13308 12174
rect 13449 11996 13745 12016
rect 13505 11994 13529 11996
rect 13585 11994 13609 11996
rect 13665 11994 13689 11996
rect 13527 11942 13529 11994
rect 13591 11942 13603 11994
rect 13665 11942 13667 11994
rect 13505 11940 13529 11942
rect 13585 11940 13609 11942
rect 13665 11940 13689 11942
rect 13449 11920 13745 11940
rect 13832 11898 13860 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 13449 10908 13745 10928
rect 13505 10906 13529 10908
rect 13585 10906 13609 10908
rect 13665 10906 13689 10908
rect 13527 10854 13529 10906
rect 13591 10854 13603 10906
rect 13665 10854 13667 10906
rect 13505 10852 13529 10854
rect 13585 10852 13609 10854
rect 13665 10852 13689 10854
rect 13449 10832 13745 10852
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13372 9586 13400 9862
rect 13449 9820 13745 9840
rect 13505 9818 13529 9820
rect 13585 9818 13609 9820
rect 13665 9818 13689 9820
rect 13527 9766 13529 9818
rect 13591 9766 13603 9818
rect 13665 9766 13667 9818
rect 13505 9764 13529 9766
rect 13585 9764 13609 9766
rect 13665 9764 13689 9766
rect 13449 9744 13745 9764
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13832 9382 13860 10066
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13188 9030 13308 9058
rect 13280 9024 13308 9030
rect 13360 9036 13412 9042
rect 13280 8996 13360 9024
rect 13360 8978 13412 8984
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8634 13216 8910
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13096 7886 13124 8366
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13004 7670 13124 7698
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12728 7262 12848 7290
rect 12636 7002 12664 7210
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12728 5574 12756 7262
rect 13004 6798 13032 7346
rect 13096 7206 13124 7670
rect 13372 7528 13400 8978
rect 13832 8838 13860 9318
rect 13924 8974 13952 9930
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13449 8732 13745 8752
rect 13505 8730 13529 8732
rect 13585 8730 13609 8732
rect 13665 8730 13689 8732
rect 13527 8678 13529 8730
rect 13591 8678 13603 8730
rect 13665 8678 13667 8730
rect 13505 8676 13529 8678
rect 13585 8676 13609 8678
rect 13665 8676 13689 8678
rect 13449 8656 13745 8676
rect 13924 8634 13952 8910
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13449 7644 13745 7664
rect 13505 7642 13529 7644
rect 13585 7642 13609 7644
rect 13665 7642 13689 7644
rect 13527 7590 13529 7642
rect 13591 7590 13603 7642
rect 13665 7590 13667 7642
rect 13505 7588 13529 7590
rect 13585 7588 13609 7590
rect 13665 7588 13689 7590
rect 13449 7568 13745 7588
rect 13372 7500 13492 7528
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13096 5930 13124 7142
rect 13358 6896 13414 6905
rect 13268 6860 13320 6866
rect 13358 6831 13360 6840
rect 13268 6802 13320 6808
rect 13412 6831 13414 6840
rect 13360 6802 13412 6808
rect 13280 6322 13308 6802
rect 13464 6746 13492 7500
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13372 6718 13492 6746
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13096 5902 13216 5930
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12636 4486 12664 5034
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12452 3692 12572 3720
rect 12452 2446 12480 3692
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12636 3233 12664 3606
rect 12622 3224 12678 3233
rect 12532 3188 12584 3194
rect 12622 3159 12678 3168
rect 12532 3130 12584 3136
rect 12544 3058 12572 3130
rect 12636 3058 12664 3159
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12544 2582 12572 2994
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12728 2530 12756 5510
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12912 4690 12940 5034
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12820 2650 12848 3878
rect 12912 2990 12940 4626
rect 13188 3942 13216 5902
rect 13266 4448 13322 4457
rect 13266 4383 13322 4392
rect 13280 4282 13308 4383
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13096 3738 13124 3878
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12990 3632 13046 3641
rect 12990 3567 13046 3576
rect 13004 3398 13032 3567
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12912 2530 12940 2586
rect 12728 2502 12940 2530
rect 12440 2440 12492 2446
rect 13004 2428 13032 3334
rect 13188 3194 13216 3470
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13188 2922 13216 3130
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 13280 2802 13308 4014
rect 12440 2382 12492 2388
rect 12728 2400 13032 2428
rect 13188 2774 13308 2802
rect 12452 1426 12480 2382
rect 12440 1420 12492 1426
rect 12440 1362 12492 1368
rect 12728 800 12756 2400
rect 13188 800 13216 2774
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13280 2446 13308 2518
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13372 2020 13400 6718
rect 13449 6556 13745 6576
rect 13505 6554 13529 6556
rect 13585 6554 13609 6556
rect 13665 6554 13689 6556
rect 13527 6502 13529 6554
rect 13591 6502 13603 6554
rect 13665 6502 13667 6554
rect 13505 6500 13529 6502
rect 13585 6500 13609 6502
rect 13665 6500 13689 6502
rect 13449 6480 13745 6500
rect 13449 5468 13745 5488
rect 13505 5466 13529 5468
rect 13585 5466 13609 5468
rect 13665 5466 13689 5468
rect 13527 5414 13529 5466
rect 13591 5414 13603 5466
rect 13665 5414 13667 5466
rect 13505 5412 13529 5414
rect 13585 5412 13609 5414
rect 13665 5412 13689 5414
rect 13449 5392 13745 5412
rect 13449 4380 13745 4400
rect 13505 4378 13529 4380
rect 13585 4378 13609 4380
rect 13665 4378 13689 4380
rect 13527 4326 13529 4378
rect 13591 4326 13603 4378
rect 13665 4326 13667 4378
rect 13505 4324 13529 4326
rect 13585 4324 13609 4326
rect 13665 4324 13689 4326
rect 13449 4304 13745 4324
rect 13818 4176 13874 4185
rect 13818 4111 13874 4120
rect 13832 4078 13860 4111
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13449 3292 13745 3312
rect 13505 3290 13529 3292
rect 13585 3290 13609 3292
rect 13665 3290 13689 3292
rect 13527 3238 13529 3290
rect 13591 3238 13603 3290
rect 13665 3238 13667 3290
rect 13505 3236 13529 3238
rect 13585 3236 13609 3238
rect 13665 3236 13689 3238
rect 13449 3216 13745 3236
rect 13832 2990 13860 3334
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13924 2582 13952 7278
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14016 4282 14044 4558
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14108 4162 14136 9046
rect 14016 4134 14136 4162
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 13449 2204 13745 2224
rect 13505 2202 13529 2204
rect 13585 2202 13609 2204
rect 13665 2202 13689 2204
rect 13527 2150 13529 2202
rect 13591 2150 13603 2202
rect 13665 2150 13667 2202
rect 13505 2148 13529 2150
rect 13585 2148 13609 2150
rect 13665 2148 13689 2150
rect 13449 2128 13745 2148
rect 13372 1992 13584 2020
rect 13556 800 13584 1992
rect 14016 800 14044 4134
rect 14200 4026 14228 11494
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14384 9518 14412 9862
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14108 3998 14228 4026
rect 14108 2310 14136 3998
rect 14292 2666 14320 4966
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14384 3194 14412 4082
rect 14476 3942 14504 12854
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12306 14872 12582
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10266 14780 10406
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14660 4826 14688 5714
rect 14648 4820 14700 4826
rect 14844 4808 14872 12242
rect 14936 6066 14964 16390
rect 15304 15706 15332 19200
rect 15658 17912 15714 17921
rect 15658 17847 15714 17856
rect 15672 16114 15700 17847
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15028 15026 15056 15506
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15016 14544 15068 14550
rect 15016 14486 15068 14492
rect 15028 14074 15056 14486
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15396 13977 15424 14214
rect 15382 13968 15438 13977
rect 15382 13903 15438 13912
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 9897 15056 13806
rect 15764 11558 15792 19200
rect 16132 15638 16160 19200
rect 16592 15910 16620 19200
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 16132 11014 16160 15574
rect 16960 12850 16988 19200
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 15014 9888 15070 9897
rect 15014 9823 15070 9832
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 14936 6038 15056 6066
rect 14922 5944 14978 5953
rect 14922 5879 14978 5888
rect 14936 5846 14964 5879
rect 14924 5840 14976 5846
rect 14924 5782 14976 5788
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14648 4762 14700 4768
rect 14752 4780 14872 4808
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14660 3942 14688 4626
rect 14752 4060 14780 4780
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14844 4214 14872 4626
rect 14936 4622 14964 5034
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 14832 4208 14884 4214
rect 14832 4150 14884 4156
rect 14752 4032 14872 4060
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14476 3738 14504 3878
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14844 3194 14872 4032
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14844 2990 14872 3130
rect 14832 2984 14884 2990
rect 14752 2944 14832 2972
rect 14292 2638 14504 2666
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 2106 14136 2246
rect 14096 2100 14148 2106
rect 14096 2042 14148 2048
rect 14476 800 14504 2638
rect 14752 1834 14780 2944
rect 14832 2926 14884 2932
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 14740 1828 14792 1834
rect 14740 1770 14792 1776
rect 14844 800 14872 2790
rect 15028 2009 15056 6038
rect 15292 4616 15344 4622
rect 15198 4584 15254 4593
rect 15292 4558 15344 4564
rect 15198 4519 15254 4528
rect 15212 3942 15240 4519
rect 15304 4078 15332 4558
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15200 3936 15252 3942
rect 15252 3896 15332 3924
rect 15200 3878 15252 3884
rect 15304 3738 15332 3896
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15212 3482 15240 3674
rect 15212 3454 15332 3482
rect 15014 2000 15070 2009
rect 15014 1935 15070 1944
rect 15304 800 15332 3454
rect 15660 1420 15712 1426
rect 15660 1362 15712 1368
rect 15672 800 15700 1362
rect 16132 800 16160 9318
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16500 800 16528 3946
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16960 800 16988 2858
rect 2962 504 3018 513
rect 2962 439 3018 448
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16946 0 17002 800
<< via2 >>
rect 2778 19488 2834 19544
rect 1766 17584 1822 17640
rect 1674 16632 1730 16688
rect 3454 17434 3510 17436
rect 3534 17434 3590 17436
rect 3614 17434 3670 17436
rect 3694 17434 3750 17436
rect 3454 17382 3480 17434
rect 3480 17382 3510 17434
rect 3534 17382 3544 17434
rect 3544 17382 3590 17434
rect 3614 17382 3660 17434
rect 3660 17382 3670 17434
rect 3694 17382 3724 17434
rect 3724 17382 3750 17434
rect 3454 17380 3510 17382
rect 3534 17380 3590 17382
rect 3614 17380 3670 17382
rect 3694 17380 3750 17382
rect 4066 18536 4122 18592
rect 3454 16346 3510 16348
rect 3534 16346 3590 16348
rect 3614 16346 3670 16348
rect 3694 16346 3750 16348
rect 3454 16294 3480 16346
rect 3480 16294 3510 16346
rect 3534 16294 3544 16346
rect 3544 16294 3590 16346
rect 3614 16294 3660 16346
rect 3660 16294 3670 16346
rect 3694 16294 3724 16346
rect 3724 16294 3750 16346
rect 3454 16292 3510 16294
rect 3534 16292 3590 16294
rect 3614 16292 3670 16294
rect 3694 16292 3750 16294
rect 1766 15680 1822 15736
rect 1674 14728 1730 14784
rect 1582 13776 1638 13832
rect 1674 12824 1730 12880
rect 2594 14884 2650 14920
rect 2594 14864 2596 14884
rect 2596 14864 2648 14884
rect 2648 14864 2650 14884
rect 3146 14320 3202 14376
rect 3454 15258 3510 15260
rect 3534 15258 3590 15260
rect 3614 15258 3670 15260
rect 3694 15258 3750 15260
rect 3454 15206 3480 15258
rect 3480 15206 3510 15258
rect 3534 15206 3544 15258
rect 3544 15206 3590 15258
rect 3614 15206 3660 15258
rect 3660 15206 3670 15258
rect 3694 15206 3724 15258
rect 3724 15206 3750 15258
rect 3454 15204 3510 15206
rect 3534 15204 3590 15206
rect 3614 15204 3670 15206
rect 3694 15204 3750 15206
rect 3514 14320 3570 14376
rect 3454 14170 3510 14172
rect 3534 14170 3590 14172
rect 3614 14170 3670 14172
rect 3694 14170 3750 14172
rect 3454 14118 3480 14170
rect 3480 14118 3510 14170
rect 3534 14118 3544 14170
rect 3544 14118 3590 14170
rect 3614 14118 3660 14170
rect 3660 14118 3670 14170
rect 3694 14118 3724 14170
rect 3724 14118 3750 14170
rect 3454 14116 3510 14118
rect 3534 14116 3590 14118
rect 3614 14116 3670 14118
rect 3694 14116 3750 14118
rect 4342 14864 4398 14920
rect 3422 13912 3478 13968
rect 3790 13912 3846 13968
rect 1674 11872 1730 11928
rect 1674 10920 1730 10976
rect 1674 10004 1676 10024
rect 1676 10004 1728 10024
rect 1728 10004 1730 10024
rect 1674 9968 1730 10004
rect 3974 13404 3976 13424
rect 3976 13404 4028 13424
rect 4028 13404 4030 13424
rect 3974 13368 4030 13404
rect 3454 13082 3510 13084
rect 3534 13082 3590 13084
rect 3614 13082 3670 13084
rect 3694 13082 3750 13084
rect 3454 13030 3480 13082
rect 3480 13030 3510 13082
rect 3534 13030 3544 13082
rect 3544 13030 3590 13082
rect 3614 13030 3660 13082
rect 3660 13030 3670 13082
rect 3694 13030 3724 13082
rect 3724 13030 3750 13082
rect 3454 13028 3510 13030
rect 3534 13028 3590 13030
rect 3614 13028 3670 13030
rect 3694 13028 3750 13030
rect 3454 11994 3510 11996
rect 3534 11994 3590 11996
rect 3614 11994 3670 11996
rect 3694 11994 3750 11996
rect 3454 11942 3480 11994
rect 3480 11942 3510 11994
rect 3534 11942 3544 11994
rect 3544 11942 3590 11994
rect 3614 11942 3660 11994
rect 3660 11942 3670 11994
rect 3694 11942 3724 11994
rect 3724 11942 3750 11994
rect 3454 11940 3510 11942
rect 3534 11940 3590 11942
rect 3614 11940 3670 11942
rect 3694 11940 3750 11942
rect 2778 9016 2834 9072
rect 1766 8064 1822 8120
rect 1674 7112 1730 7168
rect 1766 6160 1822 6216
rect 2870 5752 2926 5808
rect 2318 5208 2374 5264
rect 1490 3032 1546 3088
rect 1674 4256 1730 4312
rect 2042 3732 2098 3768
rect 2042 3712 2044 3732
rect 2044 3712 2096 3732
rect 2096 3712 2098 3732
rect 1674 3304 1730 3360
rect 2042 1400 2098 1456
rect 3454 10906 3510 10908
rect 3534 10906 3590 10908
rect 3614 10906 3670 10908
rect 3694 10906 3750 10908
rect 3454 10854 3480 10906
rect 3480 10854 3510 10906
rect 3534 10854 3544 10906
rect 3544 10854 3590 10906
rect 3614 10854 3660 10906
rect 3660 10854 3670 10906
rect 3694 10854 3724 10906
rect 3724 10854 3750 10906
rect 3454 10852 3510 10854
rect 3534 10852 3590 10854
rect 3614 10852 3670 10854
rect 3694 10852 3750 10854
rect 4526 13268 4528 13288
rect 4528 13268 4580 13288
rect 4580 13268 4582 13288
rect 4526 13232 4582 13268
rect 3454 9818 3510 9820
rect 3534 9818 3590 9820
rect 3614 9818 3670 9820
rect 3694 9818 3750 9820
rect 3454 9766 3480 9818
rect 3480 9766 3510 9818
rect 3534 9766 3544 9818
rect 3544 9766 3590 9818
rect 3614 9766 3660 9818
rect 3660 9766 3670 9818
rect 3694 9766 3724 9818
rect 3724 9766 3750 9818
rect 3454 9764 3510 9766
rect 3534 9764 3590 9766
rect 3614 9764 3670 9766
rect 3694 9764 3750 9766
rect 3454 8730 3510 8732
rect 3534 8730 3590 8732
rect 3614 8730 3670 8732
rect 3694 8730 3750 8732
rect 3454 8678 3480 8730
rect 3480 8678 3510 8730
rect 3534 8678 3544 8730
rect 3544 8678 3590 8730
rect 3614 8678 3660 8730
rect 3660 8678 3670 8730
rect 3694 8678 3724 8730
rect 3724 8678 3750 8730
rect 3454 8676 3510 8678
rect 3534 8676 3590 8678
rect 3614 8676 3670 8678
rect 3694 8676 3750 8678
rect 3454 7642 3510 7644
rect 3534 7642 3590 7644
rect 3614 7642 3670 7644
rect 3694 7642 3750 7644
rect 3454 7590 3480 7642
rect 3480 7590 3510 7642
rect 3534 7590 3544 7642
rect 3544 7590 3590 7642
rect 3614 7590 3660 7642
rect 3660 7590 3670 7642
rect 3694 7590 3724 7642
rect 3724 7590 3750 7642
rect 3454 7588 3510 7590
rect 3534 7588 3590 7590
rect 3614 7588 3670 7590
rect 3694 7588 3750 7590
rect 3454 6554 3510 6556
rect 3534 6554 3590 6556
rect 3614 6554 3670 6556
rect 3694 6554 3750 6556
rect 3454 6502 3480 6554
rect 3480 6502 3510 6554
rect 3534 6502 3544 6554
rect 3544 6502 3590 6554
rect 3614 6502 3660 6554
rect 3660 6502 3670 6554
rect 3694 6502 3724 6554
rect 3724 6502 3750 6554
rect 3454 6500 3510 6502
rect 3534 6500 3590 6502
rect 3614 6500 3670 6502
rect 3694 6500 3750 6502
rect 3454 5466 3510 5468
rect 3534 5466 3590 5468
rect 3614 5466 3670 5468
rect 3694 5466 3750 5468
rect 3454 5414 3480 5466
rect 3480 5414 3510 5466
rect 3534 5414 3544 5466
rect 3544 5414 3590 5466
rect 3614 5414 3660 5466
rect 3660 5414 3670 5466
rect 3694 5414 3724 5466
rect 3724 5414 3750 5466
rect 3454 5412 3510 5414
rect 3534 5412 3590 5414
rect 3614 5412 3670 5414
rect 3694 5412 3750 5414
rect 5953 16890 6009 16892
rect 6033 16890 6089 16892
rect 6113 16890 6169 16892
rect 6193 16890 6249 16892
rect 5953 16838 5979 16890
rect 5979 16838 6009 16890
rect 6033 16838 6043 16890
rect 6043 16838 6089 16890
rect 6113 16838 6159 16890
rect 6159 16838 6169 16890
rect 6193 16838 6223 16890
rect 6223 16838 6249 16890
rect 5953 16836 6009 16838
rect 6033 16836 6089 16838
rect 6113 16836 6169 16838
rect 6193 16836 6249 16838
rect 5078 12824 5134 12880
rect 5170 10124 5226 10160
rect 5170 10104 5172 10124
rect 5172 10104 5224 10124
rect 5224 10104 5226 10124
rect 5953 15802 6009 15804
rect 6033 15802 6089 15804
rect 6113 15802 6169 15804
rect 6193 15802 6249 15804
rect 5953 15750 5979 15802
rect 5979 15750 6009 15802
rect 6033 15750 6043 15802
rect 6043 15750 6089 15802
rect 6113 15750 6159 15802
rect 6159 15750 6169 15802
rect 6193 15750 6223 15802
rect 6223 15750 6249 15802
rect 5953 15748 6009 15750
rect 6033 15748 6089 15750
rect 6113 15748 6169 15750
rect 6193 15748 6249 15750
rect 6274 15544 6330 15600
rect 5953 14714 6009 14716
rect 6033 14714 6089 14716
rect 6113 14714 6169 14716
rect 6193 14714 6249 14716
rect 5953 14662 5979 14714
rect 5979 14662 6009 14714
rect 6033 14662 6043 14714
rect 6043 14662 6089 14714
rect 6113 14662 6159 14714
rect 6159 14662 6169 14714
rect 6193 14662 6223 14714
rect 6223 14662 6249 14714
rect 5953 14660 6009 14662
rect 6033 14660 6089 14662
rect 6113 14660 6169 14662
rect 6193 14660 6249 14662
rect 5953 13626 6009 13628
rect 6033 13626 6089 13628
rect 6113 13626 6169 13628
rect 6193 13626 6249 13628
rect 5953 13574 5979 13626
rect 5979 13574 6009 13626
rect 6033 13574 6043 13626
rect 6043 13574 6089 13626
rect 6113 13574 6159 13626
rect 6159 13574 6169 13626
rect 6193 13574 6223 13626
rect 6223 13574 6249 13626
rect 5953 13572 6009 13574
rect 6033 13572 6089 13574
rect 6113 13572 6169 13574
rect 6193 13572 6249 13574
rect 5446 10124 5502 10160
rect 5446 10104 5448 10124
rect 5448 10104 5500 10124
rect 5500 10104 5502 10124
rect 6366 14184 6422 14240
rect 6274 12688 6330 12744
rect 5953 12538 6009 12540
rect 6033 12538 6089 12540
rect 6113 12538 6169 12540
rect 6193 12538 6249 12540
rect 5953 12486 5979 12538
rect 5979 12486 6009 12538
rect 6033 12486 6043 12538
rect 6043 12486 6089 12538
rect 6113 12486 6159 12538
rect 6159 12486 6169 12538
rect 6193 12486 6223 12538
rect 6223 12486 6249 12538
rect 5953 12484 6009 12486
rect 6033 12484 6089 12486
rect 6113 12484 6169 12486
rect 6193 12484 6249 12486
rect 5953 11450 6009 11452
rect 6033 11450 6089 11452
rect 6113 11450 6169 11452
rect 6193 11450 6249 11452
rect 5953 11398 5979 11450
rect 5979 11398 6009 11450
rect 6033 11398 6043 11450
rect 6043 11398 6089 11450
rect 6113 11398 6159 11450
rect 6159 11398 6169 11450
rect 6193 11398 6223 11450
rect 6223 11398 6249 11450
rect 5953 11396 6009 11398
rect 6033 11396 6089 11398
rect 6113 11396 6169 11398
rect 6193 11396 6249 11398
rect 3454 4378 3510 4380
rect 3534 4378 3590 4380
rect 3614 4378 3670 4380
rect 3694 4378 3750 4380
rect 3454 4326 3480 4378
rect 3480 4326 3510 4378
rect 3534 4326 3544 4378
rect 3544 4326 3590 4378
rect 3614 4326 3660 4378
rect 3660 4326 3670 4378
rect 3694 4326 3724 4378
rect 3724 4326 3750 4378
rect 3454 4324 3510 4326
rect 3534 4324 3590 4326
rect 3614 4324 3670 4326
rect 3694 4324 3750 4326
rect 3974 3576 4030 3632
rect 3454 3290 3510 3292
rect 3534 3290 3590 3292
rect 3614 3290 3670 3292
rect 3694 3290 3750 3292
rect 3454 3238 3480 3290
rect 3480 3238 3510 3290
rect 3534 3238 3544 3290
rect 3544 3238 3590 3290
rect 3614 3238 3660 3290
rect 3660 3238 3670 3290
rect 3694 3238 3724 3290
rect 3724 3238 3750 3290
rect 3454 3236 3510 3238
rect 3534 3236 3590 3238
rect 3614 3236 3670 3238
rect 3694 3236 3750 3238
rect 5078 8356 5134 8392
rect 5078 8336 5080 8356
rect 5080 8336 5132 8356
rect 5132 8336 5134 8356
rect 5953 10362 6009 10364
rect 6033 10362 6089 10364
rect 6113 10362 6169 10364
rect 6193 10362 6249 10364
rect 5953 10310 5979 10362
rect 5979 10310 6009 10362
rect 6033 10310 6043 10362
rect 6043 10310 6089 10362
rect 6113 10310 6159 10362
rect 6159 10310 6169 10362
rect 6193 10310 6223 10362
rect 6223 10310 6249 10362
rect 5953 10308 6009 10310
rect 6033 10308 6089 10310
rect 6113 10308 6169 10310
rect 6193 10308 6249 10310
rect 5814 9460 5816 9480
rect 5816 9460 5868 9480
rect 5868 9460 5870 9480
rect 5814 9424 5870 9460
rect 5953 9274 6009 9276
rect 6033 9274 6089 9276
rect 6113 9274 6169 9276
rect 6193 9274 6249 9276
rect 5953 9222 5979 9274
rect 5979 9222 6009 9274
rect 6033 9222 6043 9274
rect 6043 9222 6089 9274
rect 6113 9222 6159 9274
rect 6159 9222 6169 9274
rect 6193 9222 6223 9274
rect 6223 9222 6249 9274
rect 5953 9220 6009 9222
rect 6033 9220 6089 9222
rect 6113 9220 6169 9222
rect 6193 9220 6249 9222
rect 4710 4528 4766 4584
rect 6642 15952 6698 16008
rect 7378 14764 7380 14784
rect 7380 14764 7432 14784
rect 7432 14764 7434 14784
rect 7378 14728 7434 14764
rect 7746 15408 7802 15464
rect 5953 8186 6009 8188
rect 6033 8186 6089 8188
rect 6113 8186 6169 8188
rect 6193 8186 6249 8188
rect 5953 8134 5979 8186
rect 5979 8134 6009 8186
rect 6033 8134 6043 8186
rect 6043 8134 6089 8186
rect 6113 8134 6159 8186
rect 6159 8134 6169 8186
rect 6193 8134 6223 8186
rect 6223 8134 6249 8186
rect 5953 8132 6009 8134
rect 6033 8132 6089 8134
rect 6113 8132 6169 8134
rect 6193 8132 6249 8134
rect 5953 7098 6009 7100
rect 6033 7098 6089 7100
rect 6113 7098 6169 7100
rect 6193 7098 6249 7100
rect 5953 7046 5979 7098
rect 5979 7046 6009 7098
rect 6033 7046 6043 7098
rect 6043 7046 6089 7098
rect 6113 7046 6159 7098
rect 6159 7046 6169 7098
rect 6193 7046 6223 7098
rect 6223 7046 6249 7098
rect 5953 7044 6009 7046
rect 6033 7044 6089 7046
rect 6113 7044 6169 7046
rect 6193 7044 6249 7046
rect 5953 6010 6009 6012
rect 6033 6010 6089 6012
rect 6113 6010 6169 6012
rect 6193 6010 6249 6012
rect 5953 5958 5979 6010
rect 5979 5958 6009 6010
rect 6033 5958 6043 6010
rect 6043 5958 6089 6010
rect 6113 5958 6159 6010
rect 6159 5958 6169 6010
rect 6193 5958 6223 6010
rect 6223 5958 6249 6010
rect 5953 5956 6009 5958
rect 6033 5956 6089 5958
rect 6113 5956 6169 5958
rect 6193 5956 6249 5958
rect 5953 4922 6009 4924
rect 6033 4922 6089 4924
rect 6113 4922 6169 4924
rect 6193 4922 6249 4924
rect 5953 4870 5979 4922
rect 5979 4870 6009 4922
rect 6033 4870 6043 4922
rect 6043 4870 6089 4922
rect 6113 4870 6159 4922
rect 6159 4870 6169 4922
rect 6193 4870 6223 4922
rect 6223 4870 6249 4922
rect 5953 4868 6009 4870
rect 6033 4868 6089 4870
rect 6113 4868 6169 4870
rect 6193 4868 6249 4870
rect 5170 4528 5226 4584
rect 4986 3440 5042 3496
rect 5538 3712 5594 3768
rect 4802 2896 4858 2952
rect 3454 2202 3510 2204
rect 3534 2202 3590 2204
rect 3614 2202 3670 2204
rect 3694 2202 3750 2204
rect 3454 2150 3480 2202
rect 3480 2150 3510 2202
rect 3534 2150 3544 2202
rect 3544 2150 3590 2202
rect 3614 2150 3660 2202
rect 3660 2150 3670 2202
rect 3694 2150 3724 2202
rect 3724 2150 3750 2202
rect 3454 2148 3510 2150
rect 3534 2148 3590 2150
rect 3614 2148 3670 2150
rect 3694 2148 3750 2150
rect 4986 2352 5042 2408
rect 6734 5752 6790 5808
rect 5953 3834 6009 3836
rect 6033 3834 6089 3836
rect 6113 3834 6169 3836
rect 6193 3834 6249 3836
rect 5953 3782 5979 3834
rect 5979 3782 6009 3834
rect 6033 3782 6043 3834
rect 6043 3782 6089 3834
rect 6113 3782 6159 3834
rect 6159 3782 6169 3834
rect 6193 3782 6223 3834
rect 6223 3782 6249 3834
rect 5953 3780 6009 3782
rect 6033 3780 6089 3782
rect 6113 3780 6169 3782
rect 6193 3780 6249 3782
rect 6458 3712 6514 3768
rect 6366 2760 6422 2816
rect 5953 2746 6009 2748
rect 6033 2746 6089 2748
rect 6113 2746 6169 2748
rect 6193 2746 6249 2748
rect 5953 2694 5979 2746
rect 5979 2694 6009 2746
rect 6033 2694 6043 2746
rect 6043 2694 6089 2746
rect 6113 2694 6159 2746
rect 6159 2694 6169 2746
rect 6193 2694 6223 2746
rect 6223 2694 6249 2746
rect 5953 2692 6009 2694
rect 6033 2692 6089 2694
rect 6113 2692 6169 2694
rect 6193 2692 6249 2694
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8478 17434
rect 8478 17382 8508 17434
rect 8532 17382 8542 17434
rect 8542 17382 8588 17434
rect 8612 17382 8658 17434
rect 8658 17382 8668 17434
rect 8692 17382 8722 17434
rect 8722 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8758 16496 8814 16552
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8478 16346
rect 8478 16294 8508 16346
rect 8532 16294 8542 16346
rect 8542 16294 8588 16346
rect 8612 16294 8658 16346
rect 8658 16294 8668 16346
rect 8692 16294 8722 16346
rect 8722 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8206 16088 8262 16144
rect 8666 16108 8722 16144
rect 8666 16088 8668 16108
rect 8668 16088 8720 16108
rect 8720 16088 8722 16108
rect 8022 15700 8078 15736
rect 8022 15680 8024 15700
rect 8024 15680 8076 15700
rect 8076 15680 8078 15700
rect 7930 14864 7986 14920
rect 8574 15700 8630 15736
rect 8574 15680 8576 15700
rect 8576 15680 8628 15700
rect 8628 15680 8630 15700
rect 9218 16088 9274 16144
rect 9034 15680 9090 15736
rect 8758 15544 8814 15600
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8478 15258
rect 8478 15206 8508 15258
rect 8532 15206 8542 15258
rect 8542 15206 8588 15258
rect 8612 15206 8658 15258
rect 8658 15206 8668 15258
rect 8692 15206 8722 15258
rect 8722 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8758 14764 8760 14784
rect 8760 14764 8812 14784
rect 8812 14764 8814 14784
rect 8758 14728 8814 14764
rect 8758 14476 8814 14512
rect 8758 14456 8760 14476
rect 8760 14456 8812 14476
rect 8812 14456 8814 14476
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8478 14170
rect 8478 14118 8508 14170
rect 8532 14118 8542 14170
rect 8542 14118 8588 14170
rect 8612 14118 8658 14170
rect 8658 14118 8668 14170
rect 8692 14118 8722 14170
rect 8722 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8390 13812 8392 13832
rect 8392 13812 8444 13832
rect 8444 13812 8446 13832
rect 8390 13776 8446 13812
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8478 13082
rect 8478 13030 8508 13082
rect 8532 13030 8542 13082
rect 8542 13030 8588 13082
rect 8612 13030 8658 13082
rect 8658 13030 8668 13082
rect 8692 13030 8722 13082
rect 8722 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 9126 14476 9182 14512
rect 9126 14456 9128 14476
rect 9128 14456 9180 14476
rect 9180 14456 9182 14476
rect 9402 15680 9458 15736
rect 9310 13776 9366 13832
rect 9218 12960 9274 13016
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8478 11994
rect 8478 11942 8508 11994
rect 8532 11942 8542 11994
rect 8542 11942 8588 11994
rect 8612 11942 8658 11994
rect 8658 11942 8668 11994
rect 8692 11942 8722 11994
rect 8722 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 7838 10548 7840 10568
rect 7840 10548 7892 10568
rect 7892 10548 7894 10568
rect 7838 10512 7894 10548
rect 7194 7792 7250 7848
rect 7378 5752 7434 5808
rect 7746 5108 7748 5128
rect 7748 5108 7800 5128
rect 7800 5108 7802 5128
rect 7746 5072 7802 5108
rect 7562 4120 7618 4176
rect 7378 3984 7434 4040
rect 7746 4528 7802 4584
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8478 10906
rect 8478 10854 8508 10906
rect 8532 10854 8542 10906
rect 8542 10854 8588 10906
rect 8612 10854 8658 10906
rect 8658 10854 8668 10906
rect 8692 10854 8722 10906
rect 8722 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8758 10532 8814 10568
rect 8758 10512 8760 10532
rect 8760 10512 8812 10532
rect 8812 10512 8814 10532
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8478 9818
rect 8478 9766 8508 9818
rect 8532 9766 8542 9818
rect 8542 9766 8588 9818
rect 8612 9766 8658 9818
rect 8658 9766 8668 9818
rect 8692 9766 8722 9818
rect 8722 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8478 8730
rect 8478 8678 8508 8730
rect 8532 8678 8542 8730
rect 8542 8678 8588 8730
rect 8612 8678 8658 8730
rect 8658 8678 8668 8730
rect 8692 8678 8722 8730
rect 8722 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8482 8472 8538 8528
rect 8666 7928 8722 7984
rect 8942 8744 8998 8800
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8478 7642
rect 8478 7590 8508 7642
rect 8532 7590 8542 7642
rect 8542 7590 8588 7642
rect 8612 7590 8658 7642
rect 8658 7590 8668 7642
rect 8692 7590 8722 7642
rect 8722 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8942 7384 8998 7440
rect 8850 7112 8906 7168
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8478 6554
rect 8478 6502 8508 6554
rect 8532 6502 8542 6554
rect 8542 6502 8588 6554
rect 8612 6502 8658 6554
rect 8658 6502 8668 6554
rect 8692 6502 8722 6554
rect 8722 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8478 5466
rect 8478 5414 8508 5466
rect 8532 5414 8542 5466
rect 8542 5414 8588 5466
rect 8612 5414 8658 5466
rect 8658 5414 8668 5466
rect 8692 5414 8722 5466
rect 8722 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8482 5108 8484 5128
rect 8484 5108 8536 5128
rect 8536 5108 8538 5128
rect 8482 5072 8538 5108
rect 9218 9424 9274 9480
rect 9126 9016 9182 9072
rect 9678 15272 9734 15328
rect 9954 16496 10010 16552
rect 9862 13096 9918 13152
rect 10138 14764 10140 14784
rect 10140 14764 10192 14784
rect 10192 14764 10194 14784
rect 10138 14728 10194 14764
rect 10046 13368 10102 13424
rect 9954 12688 10010 12744
rect 9954 11736 10010 11792
rect 10950 16890 11006 16892
rect 11030 16890 11086 16892
rect 11110 16890 11166 16892
rect 11190 16890 11246 16892
rect 10950 16838 10976 16890
rect 10976 16838 11006 16890
rect 11030 16838 11040 16890
rect 11040 16838 11086 16890
rect 11110 16838 11156 16890
rect 11156 16838 11166 16890
rect 11190 16838 11220 16890
rect 11220 16838 11246 16890
rect 10950 16836 11006 16838
rect 11030 16836 11086 16838
rect 11110 16836 11166 16838
rect 11190 16836 11246 16838
rect 10950 15802 11006 15804
rect 11030 15802 11086 15804
rect 11110 15802 11166 15804
rect 11190 15802 11246 15804
rect 10950 15750 10976 15802
rect 10976 15750 11006 15802
rect 11030 15750 11040 15802
rect 11040 15750 11086 15802
rect 11110 15750 11156 15802
rect 11156 15750 11166 15802
rect 11190 15750 11220 15802
rect 11220 15750 11246 15802
rect 10950 15748 11006 15750
rect 11030 15748 11086 15750
rect 11110 15748 11166 15750
rect 11190 15748 11246 15750
rect 10782 15000 10838 15056
rect 9954 9324 9956 9344
rect 9956 9324 10008 9344
rect 10008 9324 10010 9344
rect 9954 9288 10010 9324
rect 9586 8336 9642 8392
rect 9586 8236 9588 8256
rect 9588 8236 9640 8256
rect 9640 8236 9642 8256
rect 9586 8200 9642 8236
rect 9218 7928 9274 7984
rect 9126 7520 9182 7576
rect 9034 7112 9090 7168
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8478 4378
rect 8478 4326 8508 4378
rect 8532 4326 8542 4378
rect 8542 4326 8588 4378
rect 8612 4326 8658 4378
rect 8658 4326 8668 4378
rect 8692 4326 8722 4378
rect 8722 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8478 3290
rect 8478 3238 8508 3290
rect 8532 3238 8542 3290
rect 8542 3238 8588 3290
rect 8612 3238 8658 3290
rect 8658 3238 8668 3290
rect 8692 3238 8722 3290
rect 8722 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8942 4256 8998 4312
rect 9126 4120 9182 4176
rect 9126 3712 9182 3768
rect 8850 3032 8906 3088
rect 9586 7792 9642 7848
rect 10138 9016 10194 9072
rect 10046 6840 10102 6896
rect 9586 5208 9642 5264
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8478 2202
rect 8478 2150 8508 2202
rect 8532 2150 8542 2202
rect 8542 2150 8588 2202
rect 8612 2150 8658 2202
rect 8658 2150 8668 2202
rect 8692 2150 8722 2202
rect 8722 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 10598 11736 10654 11792
rect 10950 14714 11006 14716
rect 11030 14714 11086 14716
rect 11110 14714 11166 14716
rect 11190 14714 11246 14716
rect 10950 14662 10976 14714
rect 10976 14662 11006 14714
rect 11030 14662 11040 14714
rect 11040 14662 11086 14714
rect 11110 14662 11156 14714
rect 11156 14662 11166 14714
rect 11190 14662 11220 14714
rect 11220 14662 11246 14714
rect 10950 14660 11006 14662
rect 11030 14660 11086 14662
rect 11110 14660 11166 14662
rect 11190 14660 11246 14662
rect 11518 13912 11574 13968
rect 10950 13626 11006 13628
rect 11030 13626 11086 13628
rect 11110 13626 11166 13628
rect 11190 13626 11246 13628
rect 10950 13574 10976 13626
rect 10976 13574 11006 13626
rect 11030 13574 11040 13626
rect 11040 13574 11086 13626
rect 11110 13574 11156 13626
rect 11156 13574 11166 13626
rect 11190 13574 11220 13626
rect 11220 13574 11246 13626
rect 10950 13572 11006 13574
rect 11030 13572 11086 13574
rect 11110 13572 11166 13574
rect 11190 13572 11246 13574
rect 11794 15972 11850 16008
rect 11794 15952 11796 15972
rect 11796 15952 11848 15972
rect 11848 15952 11850 15972
rect 11518 13404 11520 13424
rect 11520 13404 11572 13424
rect 11572 13404 11574 13424
rect 10950 12538 11006 12540
rect 11030 12538 11086 12540
rect 11110 12538 11166 12540
rect 11190 12538 11246 12540
rect 10950 12486 10976 12538
rect 10976 12486 11006 12538
rect 11030 12486 11040 12538
rect 11040 12486 11086 12538
rect 11110 12486 11156 12538
rect 11156 12486 11166 12538
rect 11190 12486 11220 12538
rect 11220 12486 11246 12538
rect 10950 12484 11006 12486
rect 11030 12484 11086 12486
rect 11110 12484 11166 12486
rect 11190 12484 11246 12486
rect 11518 13368 11574 13404
rect 11518 13268 11520 13288
rect 11520 13268 11572 13288
rect 11572 13268 11574 13288
rect 11518 13232 11574 13268
rect 11426 13096 11482 13152
rect 11518 12824 11574 12880
rect 10950 11450 11006 11452
rect 11030 11450 11086 11452
rect 11110 11450 11166 11452
rect 11190 11450 11246 11452
rect 10950 11398 10976 11450
rect 10976 11398 11006 11450
rect 11030 11398 11040 11450
rect 11040 11398 11086 11450
rect 11110 11398 11156 11450
rect 11156 11398 11166 11450
rect 11190 11398 11220 11450
rect 11220 11398 11246 11450
rect 10950 11396 11006 11398
rect 11030 11396 11086 11398
rect 11110 11396 11166 11398
rect 11190 11396 11246 11398
rect 10598 9832 10654 9888
rect 11518 11348 11574 11384
rect 11518 11328 11520 11348
rect 11520 11328 11572 11348
rect 11572 11328 11574 11348
rect 11518 11192 11574 11248
rect 10950 10362 11006 10364
rect 11030 10362 11086 10364
rect 11110 10362 11166 10364
rect 11190 10362 11246 10364
rect 10950 10310 10976 10362
rect 10976 10310 11006 10362
rect 11030 10310 11040 10362
rect 11040 10310 11086 10362
rect 11110 10310 11156 10362
rect 11156 10310 11166 10362
rect 11190 10310 11220 10362
rect 11220 10310 11246 10362
rect 10950 10308 11006 10310
rect 11030 10308 11086 10310
rect 11110 10308 11166 10310
rect 11190 10308 11246 10310
rect 10950 9274 11006 9276
rect 11030 9274 11086 9276
rect 11110 9274 11166 9276
rect 11190 9274 11246 9276
rect 10950 9222 10976 9274
rect 10976 9222 11006 9274
rect 11030 9222 11040 9274
rect 11040 9222 11086 9274
rect 11110 9222 11156 9274
rect 11156 9222 11166 9274
rect 11190 9222 11220 9274
rect 11220 9222 11246 9274
rect 10950 9220 11006 9222
rect 11030 9220 11086 9222
rect 11110 9220 11166 9222
rect 11190 9220 11246 9222
rect 10874 9016 10930 9072
rect 10950 8186 11006 8188
rect 11030 8186 11086 8188
rect 11110 8186 11166 8188
rect 11190 8186 11246 8188
rect 10950 8134 10976 8186
rect 10976 8134 11006 8186
rect 11030 8134 11040 8186
rect 11040 8134 11086 8186
rect 11110 8134 11156 8186
rect 11156 8134 11166 8186
rect 11190 8134 11220 8186
rect 11220 8134 11246 8186
rect 10950 8132 11006 8134
rect 11030 8132 11086 8134
rect 11110 8132 11166 8134
rect 11190 8132 11246 8134
rect 10950 7098 11006 7100
rect 11030 7098 11086 7100
rect 11110 7098 11166 7100
rect 11190 7098 11246 7100
rect 10950 7046 10976 7098
rect 10976 7046 11006 7098
rect 11030 7046 11040 7098
rect 11040 7046 11086 7098
rect 11110 7046 11156 7098
rect 11156 7046 11166 7098
rect 11190 7046 11220 7098
rect 11220 7046 11246 7098
rect 10950 7044 11006 7046
rect 11030 7044 11086 7046
rect 11110 7044 11166 7046
rect 11190 7044 11246 7046
rect 10046 4528 10102 4584
rect 9678 3304 9734 3360
rect 9770 2760 9826 2816
rect 9954 3168 10010 3224
rect 11702 9424 11758 9480
rect 10950 6010 11006 6012
rect 11030 6010 11086 6012
rect 11110 6010 11166 6012
rect 11190 6010 11246 6012
rect 10950 5958 10976 6010
rect 10976 5958 11006 6010
rect 11030 5958 11040 6010
rect 11040 5958 11086 6010
rect 11110 5958 11156 6010
rect 11156 5958 11166 6010
rect 11190 5958 11220 6010
rect 11220 5958 11246 6010
rect 10950 5956 11006 5958
rect 11030 5956 11086 5958
rect 11110 5956 11166 5958
rect 11190 5956 11246 5958
rect 10598 4392 10654 4448
rect 10322 3848 10378 3904
rect 10138 3440 10194 3496
rect 10230 3032 10286 3088
rect 10046 2760 10102 2816
rect 10506 3304 10562 3360
rect 10950 4922 11006 4924
rect 11030 4922 11086 4924
rect 11110 4922 11166 4924
rect 11190 4922 11246 4924
rect 10950 4870 10976 4922
rect 10976 4870 11006 4922
rect 11030 4870 11040 4922
rect 11040 4870 11086 4922
rect 11110 4870 11156 4922
rect 11156 4870 11166 4922
rect 11190 4870 11220 4922
rect 11220 4870 11246 4922
rect 10950 4868 11006 4870
rect 11030 4868 11086 4870
rect 11110 4868 11166 4870
rect 11190 4868 11246 4870
rect 10874 4004 10930 4040
rect 10874 3984 10876 4004
rect 10876 3984 10928 4004
rect 10928 3984 10930 4004
rect 10950 3834 11006 3836
rect 11030 3834 11086 3836
rect 11110 3834 11166 3836
rect 11190 3834 11246 3836
rect 10950 3782 10976 3834
rect 10976 3782 11006 3834
rect 11030 3782 11040 3834
rect 11040 3782 11086 3834
rect 11110 3782 11156 3834
rect 11156 3782 11166 3834
rect 11190 3782 11220 3834
rect 11220 3782 11246 3834
rect 10950 3780 11006 3782
rect 11030 3780 11086 3782
rect 11110 3780 11166 3782
rect 11190 3780 11246 3782
rect 10950 2746 11006 2748
rect 11030 2746 11086 2748
rect 11110 2746 11166 2748
rect 11190 2746 11246 2748
rect 10950 2694 10976 2746
rect 10976 2694 11006 2746
rect 11030 2694 11040 2746
rect 11040 2694 11086 2746
rect 11110 2694 11156 2746
rect 11156 2694 11166 2746
rect 11190 2694 11220 2746
rect 11220 2694 11246 2746
rect 10950 2692 11006 2694
rect 11030 2692 11086 2694
rect 11110 2692 11166 2694
rect 11190 2692 11246 2694
rect 11702 7948 11758 7984
rect 11702 7928 11704 7948
rect 11704 7928 11756 7948
rect 11756 7928 11758 7948
rect 12438 17176 12494 17232
rect 12162 15428 12218 15464
rect 12162 15408 12164 15428
rect 12164 15408 12216 15428
rect 12216 15408 12218 15428
rect 12162 14884 12218 14920
rect 12162 14864 12164 14884
rect 12164 14864 12216 14884
rect 12216 14864 12218 14884
rect 12530 13368 12586 13424
rect 12530 13268 12532 13288
rect 12532 13268 12584 13288
rect 12584 13268 12586 13288
rect 12530 13232 12586 13268
rect 12254 11736 12310 11792
rect 11610 3576 11666 3632
rect 12070 3612 12072 3632
rect 12072 3612 12124 3632
rect 12124 3612 12126 3632
rect 12070 3576 12126 3612
rect 12254 3340 12256 3360
rect 12256 3340 12308 3360
rect 12308 3340 12310 3360
rect 12254 3304 12310 3340
rect 11978 3052 12034 3088
rect 11978 3032 11980 3052
rect 11980 3032 12032 3052
rect 12032 3032 12034 3052
rect 12070 2896 12126 2952
rect 12714 13368 12770 13424
rect 13449 17434 13505 17436
rect 13529 17434 13585 17436
rect 13609 17434 13665 17436
rect 13689 17434 13745 17436
rect 13449 17382 13475 17434
rect 13475 17382 13505 17434
rect 13529 17382 13539 17434
rect 13539 17382 13585 17434
rect 13609 17382 13655 17434
rect 13655 17382 13665 17434
rect 13689 17382 13719 17434
rect 13719 17382 13745 17434
rect 13449 17380 13505 17382
rect 13529 17380 13585 17382
rect 13609 17380 13665 17382
rect 13689 17380 13745 17382
rect 13449 16346 13505 16348
rect 13529 16346 13585 16348
rect 13609 16346 13665 16348
rect 13689 16346 13745 16348
rect 13449 16294 13475 16346
rect 13475 16294 13505 16346
rect 13529 16294 13539 16346
rect 13539 16294 13585 16346
rect 13609 16294 13655 16346
rect 13655 16294 13665 16346
rect 13689 16294 13719 16346
rect 13719 16294 13745 16346
rect 13449 16292 13505 16294
rect 13529 16292 13585 16294
rect 13609 16292 13665 16294
rect 13689 16292 13745 16294
rect 13449 15258 13505 15260
rect 13529 15258 13585 15260
rect 13609 15258 13665 15260
rect 13689 15258 13745 15260
rect 13449 15206 13475 15258
rect 13475 15206 13505 15258
rect 13529 15206 13539 15258
rect 13539 15206 13585 15258
rect 13609 15206 13655 15258
rect 13655 15206 13665 15258
rect 13689 15206 13719 15258
rect 13719 15206 13745 15258
rect 13449 15204 13505 15206
rect 13529 15204 13585 15206
rect 13609 15204 13665 15206
rect 13689 15204 13745 15206
rect 13449 14170 13505 14172
rect 13529 14170 13585 14172
rect 13609 14170 13665 14172
rect 13689 14170 13745 14172
rect 13449 14118 13475 14170
rect 13475 14118 13505 14170
rect 13529 14118 13539 14170
rect 13539 14118 13585 14170
rect 13609 14118 13655 14170
rect 13655 14118 13665 14170
rect 13689 14118 13719 14170
rect 13719 14118 13745 14170
rect 13449 14116 13505 14118
rect 13529 14116 13585 14118
rect 13609 14116 13665 14118
rect 13689 14116 13745 14118
rect 12898 12724 12900 12744
rect 12900 12724 12952 12744
rect 12952 12724 12954 12744
rect 12898 12688 12954 12724
rect 13449 13082 13505 13084
rect 13529 13082 13585 13084
rect 13609 13082 13665 13084
rect 13689 13082 13745 13084
rect 13449 13030 13475 13082
rect 13475 13030 13505 13082
rect 13529 13030 13539 13082
rect 13539 13030 13585 13082
rect 13609 13030 13655 13082
rect 13655 13030 13665 13082
rect 13689 13030 13719 13082
rect 13719 13030 13745 13082
rect 13449 13028 13505 13030
rect 13529 13028 13585 13030
rect 13609 13028 13665 13030
rect 13689 13028 13745 13030
rect 14094 15000 14150 15056
rect 13449 11994 13505 11996
rect 13529 11994 13585 11996
rect 13609 11994 13665 11996
rect 13689 11994 13745 11996
rect 13449 11942 13475 11994
rect 13475 11942 13505 11994
rect 13529 11942 13539 11994
rect 13539 11942 13585 11994
rect 13609 11942 13655 11994
rect 13655 11942 13665 11994
rect 13689 11942 13719 11994
rect 13719 11942 13745 11994
rect 13449 11940 13505 11942
rect 13529 11940 13585 11942
rect 13609 11940 13665 11942
rect 13689 11940 13745 11942
rect 13449 10906 13505 10908
rect 13529 10906 13585 10908
rect 13609 10906 13665 10908
rect 13689 10906 13745 10908
rect 13449 10854 13475 10906
rect 13475 10854 13505 10906
rect 13529 10854 13539 10906
rect 13539 10854 13585 10906
rect 13609 10854 13655 10906
rect 13655 10854 13665 10906
rect 13689 10854 13719 10906
rect 13719 10854 13745 10906
rect 13449 10852 13505 10854
rect 13529 10852 13585 10854
rect 13609 10852 13665 10854
rect 13689 10852 13745 10854
rect 13449 9818 13505 9820
rect 13529 9818 13585 9820
rect 13609 9818 13665 9820
rect 13689 9818 13745 9820
rect 13449 9766 13475 9818
rect 13475 9766 13505 9818
rect 13529 9766 13539 9818
rect 13539 9766 13585 9818
rect 13609 9766 13655 9818
rect 13655 9766 13665 9818
rect 13689 9766 13719 9818
rect 13719 9766 13745 9818
rect 13449 9764 13505 9766
rect 13529 9764 13585 9766
rect 13609 9764 13665 9766
rect 13689 9764 13745 9766
rect 13449 8730 13505 8732
rect 13529 8730 13585 8732
rect 13609 8730 13665 8732
rect 13689 8730 13745 8732
rect 13449 8678 13475 8730
rect 13475 8678 13505 8730
rect 13529 8678 13539 8730
rect 13539 8678 13585 8730
rect 13609 8678 13655 8730
rect 13655 8678 13665 8730
rect 13689 8678 13719 8730
rect 13719 8678 13745 8730
rect 13449 8676 13505 8678
rect 13529 8676 13585 8678
rect 13609 8676 13665 8678
rect 13689 8676 13745 8678
rect 13449 7642 13505 7644
rect 13529 7642 13585 7644
rect 13609 7642 13665 7644
rect 13689 7642 13745 7644
rect 13449 7590 13475 7642
rect 13475 7590 13505 7642
rect 13529 7590 13539 7642
rect 13539 7590 13585 7642
rect 13609 7590 13655 7642
rect 13655 7590 13665 7642
rect 13689 7590 13719 7642
rect 13719 7590 13745 7642
rect 13449 7588 13505 7590
rect 13529 7588 13585 7590
rect 13609 7588 13665 7590
rect 13689 7588 13745 7590
rect 13358 6860 13414 6896
rect 13358 6840 13360 6860
rect 13360 6840 13412 6860
rect 13412 6840 13414 6860
rect 12622 3168 12678 3224
rect 13266 4392 13322 4448
rect 12990 3576 13046 3632
rect 13449 6554 13505 6556
rect 13529 6554 13585 6556
rect 13609 6554 13665 6556
rect 13689 6554 13745 6556
rect 13449 6502 13475 6554
rect 13475 6502 13505 6554
rect 13529 6502 13539 6554
rect 13539 6502 13585 6554
rect 13609 6502 13655 6554
rect 13655 6502 13665 6554
rect 13689 6502 13719 6554
rect 13719 6502 13745 6554
rect 13449 6500 13505 6502
rect 13529 6500 13585 6502
rect 13609 6500 13665 6502
rect 13689 6500 13745 6502
rect 13449 5466 13505 5468
rect 13529 5466 13585 5468
rect 13609 5466 13665 5468
rect 13689 5466 13745 5468
rect 13449 5414 13475 5466
rect 13475 5414 13505 5466
rect 13529 5414 13539 5466
rect 13539 5414 13585 5466
rect 13609 5414 13655 5466
rect 13655 5414 13665 5466
rect 13689 5414 13719 5466
rect 13719 5414 13745 5466
rect 13449 5412 13505 5414
rect 13529 5412 13585 5414
rect 13609 5412 13665 5414
rect 13689 5412 13745 5414
rect 13449 4378 13505 4380
rect 13529 4378 13585 4380
rect 13609 4378 13665 4380
rect 13689 4378 13745 4380
rect 13449 4326 13475 4378
rect 13475 4326 13505 4378
rect 13529 4326 13539 4378
rect 13539 4326 13585 4378
rect 13609 4326 13655 4378
rect 13655 4326 13665 4378
rect 13689 4326 13719 4378
rect 13719 4326 13745 4378
rect 13449 4324 13505 4326
rect 13529 4324 13585 4326
rect 13609 4324 13665 4326
rect 13689 4324 13745 4326
rect 13818 4120 13874 4176
rect 13449 3290 13505 3292
rect 13529 3290 13585 3292
rect 13609 3290 13665 3292
rect 13689 3290 13745 3292
rect 13449 3238 13475 3290
rect 13475 3238 13505 3290
rect 13529 3238 13539 3290
rect 13539 3238 13585 3290
rect 13609 3238 13655 3290
rect 13655 3238 13665 3290
rect 13689 3238 13719 3290
rect 13719 3238 13745 3290
rect 13449 3236 13505 3238
rect 13529 3236 13585 3238
rect 13609 3236 13665 3238
rect 13689 3236 13745 3238
rect 13449 2202 13505 2204
rect 13529 2202 13585 2204
rect 13609 2202 13665 2204
rect 13689 2202 13745 2204
rect 13449 2150 13475 2202
rect 13475 2150 13505 2202
rect 13529 2150 13539 2202
rect 13539 2150 13585 2202
rect 13609 2150 13655 2202
rect 13655 2150 13665 2202
rect 13689 2150 13719 2202
rect 13719 2150 13745 2202
rect 13449 2148 13505 2150
rect 13529 2148 13585 2150
rect 13609 2148 13665 2150
rect 13689 2148 13745 2150
rect 15658 17856 15714 17912
rect 15382 13912 15438 13968
rect 15014 9832 15070 9888
rect 14922 5888 14978 5944
rect 15198 4528 15254 4584
rect 15014 1944 15070 2000
rect 2962 448 3018 504
<< metal3 >>
rect 0 19546 800 19576
rect 2773 19546 2839 19549
rect 0 19544 2839 19546
rect 0 19488 2778 19544
rect 2834 19488 2839 19544
rect 0 19486 2839 19488
rect 0 19456 800 19486
rect 2773 19483 2839 19486
rect 0 18594 800 18624
rect 4061 18594 4127 18597
rect 0 18592 4127 18594
rect 0 18536 4066 18592
rect 4122 18536 4127 18592
rect 0 18534 4127 18536
rect 0 18504 800 18534
rect 4061 18531 4127 18534
rect 15653 17914 15719 17917
rect 16400 17914 17200 17944
rect 15653 17912 17200 17914
rect 15653 17856 15658 17912
rect 15714 17856 17200 17912
rect 15653 17854 17200 17856
rect 15653 17851 15719 17854
rect 16400 17824 17200 17854
rect 0 17642 800 17672
rect 1761 17642 1827 17645
rect 0 17640 1827 17642
rect 0 17584 1766 17640
rect 1822 17584 1827 17640
rect 0 17582 1827 17584
rect 0 17552 800 17582
rect 1761 17579 1827 17582
rect 3442 17440 3762 17441
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3762 17440
rect 3442 17375 3762 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 13437 17440 13757 17441
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 17375 13757 17376
rect 11646 17172 11652 17236
rect 11716 17234 11722 17236
rect 12433 17234 12499 17237
rect 11716 17232 12499 17234
rect 11716 17176 12438 17232
rect 12494 17176 12499 17232
rect 11716 17174 12499 17176
rect 11716 17172 11722 17174
rect 12433 17171 12499 17174
rect 5941 16896 6261 16897
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 16831 6261 16832
rect 10938 16896 11258 16897
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11258 16896
rect 10938 16831 11258 16832
rect 0 16690 800 16720
rect 1669 16690 1735 16693
rect 0 16688 1735 16690
rect 0 16632 1674 16688
rect 1730 16632 1735 16688
rect 0 16630 1735 16632
rect 0 16600 800 16630
rect 1669 16627 1735 16630
rect 8753 16554 8819 16557
rect 9949 16554 10015 16557
rect 8753 16552 10015 16554
rect 8753 16496 8758 16552
rect 8814 16496 9954 16552
rect 10010 16496 10015 16552
rect 8753 16494 10015 16496
rect 8753 16491 8819 16494
rect 9949 16491 10015 16494
rect 3442 16352 3762 16353
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3762 16352
rect 3442 16287 3762 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 13437 16352 13757 16353
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 16287 13757 16288
rect 8201 16146 8267 16149
rect 8661 16146 8727 16149
rect 9213 16146 9279 16149
rect 8201 16144 9279 16146
rect 8201 16088 8206 16144
rect 8262 16088 8666 16144
rect 8722 16088 9218 16144
rect 9274 16088 9279 16144
rect 8201 16086 9279 16088
rect 8201 16083 8267 16086
rect 8661 16083 8727 16086
rect 9213 16083 9279 16086
rect 6637 16010 6703 16013
rect 11789 16010 11855 16013
rect 6637 16008 11855 16010
rect 6637 15952 6642 16008
rect 6698 15952 11794 16008
rect 11850 15952 11855 16008
rect 6637 15950 11855 15952
rect 6637 15947 6703 15950
rect 11789 15947 11855 15950
rect 5941 15808 6261 15809
rect 0 15738 800 15768
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 15743 6261 15744
rect 10938 15808 11258 15809
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11258 15808
rect 10938 15743 11258 15744
rect 1761 15738 1827 15741
rect 0 15736 1827 15738
rect 0 15680 1766 15736
rect 1822 15680 1827 15736
rect 0 15678 1827 15680
rect 0 15648 800 15678
rect 1761 15675 1827 15678
rect 8017 15738 8083 15741
rect 8569 15738 8635 15741
rect 8017 15736 8635 15738
rect 8017 15680 8022 15736
rect 8078 15680 8574 15736
rect 8630 15680 8635 15736
rect 8017 15678 8635 15680
rect 8017 15675 8083 15678
rect 8569 15675 8635 15678
rect 9029 15738 9095 15741
rect 9397 15738 9463 15741
rect 9029 15736 9463 15738
rect 9029 15680 9034 15736
rect 9090 15680 9402 15736
rect 9458 15680 9463 15736
rect 9029 15678 9463 15680
rect 9029 15675 9095 15678
rect 9397 15675 9463 15678
rect 6269 15602 6335 15605
rect 8753 15602 8819 15605
rect 6269 15600 8819 15602
rect 6269 15544 6274 15600
rect 6330 15544 8758 15600
rect 8814 15544 8819 15600
rect 6269 15542 8819 15544
rect 6269 15539 6335 15542
rect 8753 15539 8819 15542
rect 7741 15466 7807 15469
rect 12157 15466 12223 15469
rect 7741 15464 12223 15466
rect 7741 15408 7746 15464
rect 7802 15408 12162 15464
rect 12218 15408 12223 15464
rect 7741 15406 12223 15408
rect 7741 15403 7807 15406
rect 12157 15403 12223 15406
rect 9673 15330 9739 15333
rect 9630 15328 9739 15330
rect 9630 15272 9678 15328
rect 9734 15272 9739 15328
rect 9630 15267 9739 15272
rect 3442 15264 3762 15265
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3762 15264
rect 3442 15199 3762 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 2589 14922 2655 14925
rect 4337 14922 4403 14925
rect 7925 14922 7991 14925
rect 8886 14922 8892 14924
rect 2589 14920 7436 14922
rect 2589 14864 2594 14920
rect 2650 14864 4342 14920
rect 4398 14864 7436 14920
rect 2589 14862 7436 14864
rect 2589 14859 2655 14862
rect 4337 14859 4403 14862
rect 0 14786 800 14816
rect 7376 14789 7436 14862
rect 7925 14920 8892 14922
rect 7925 14864 7930 14920
rect 7986 14864 8892 14920
rect 7925 14862 8892 14864
rect 7925 14859 7991 14862
rect 8886 14860 8892 14862
rect 8956 14922 8962 14924
rect 9630 14922 9690 15267
rect 13437 15264 13757 15265
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 15199 13757 15200
rect 10777 15058 10843 15061
rect 14089 15058 14155 15061
rect 10777 15056 14155 15058
rect 10777 15000 10782 15056
rect 10838 15000 14094 15056
rect 14150 15000 14155 15056
rect 10777 14998 14155 15000
rect 10777 14995 10843 14998
rect 14089 14995 14155 14998
rect 12157 14922 12223 14925
rect 8956 14920 12223 14922
rect 8956 14864 12162 14920
rect 12218 14864 12223 14920
rect 8956 14862 12223 14864
rect 8956 14860 8962 14862
rect 12157 14859 12223 14862
rect 1669 14786 1735 14789
rect 0 14784 1735 14786
rect 0 14728 1674 14784
rect 1730 14728 1735 14784
rect 0 14726 1735 14728
rect 0 14696 800 14726
rect 1669 14723 1735 14726
rect 7373 14786 7439 14789
rect 8753 14786 8819 14789
rect 10133 14786 10199 14789
rect 7373 14784 10199 14786
rect 7373 14728 7378 14784
rect 7434 14728 8758 14784
rect 8814 14728 10138 14784
rect 10194 14728 10199 14784
rect 7373 14726 10199 14728
rect 7373 14723 7439 14726
rect 8753 14723 8819 14726
rect 10133 14723 10199 14726
rect 5941 14720 6261 14721
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 14655 6261 14656
rect 10938 14720 11258 14721
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11258 14720
rect 10938 14655 11258 14656
rect 8753 14514 8819 14517
rect 9121 14514 9187 14517
rect 8753 14512 9187 14514
rect 8753 14456 8758 14512
rect 8814 14456 9126 14512
rect 9182 14456 9187 14512
rect 8753 14454 9187 14456
rect 8753 14451 8819 14454
rect 9121 14451 9187 14454
rect 3141 14378 3207 14381
rect 3509 14378 3575 14381
rect 3141 14376 3575 14378
rect 3141 14320 3146 14376
rect 3202 14320 3514 14376
rect 3570 14320 3575 14376
rect 3141 14318 3575 14320
rect 3141 14315 3207 14318
rect 3509 14315 3575 14318
rect 5574 14180 5580 14244
rect 5644 14242 5650 14244
rect 6361 14242 6427 14245
rect 5644 14240 6427 14242
rect 5644 14184 6366 14240
rect 6422 14184 6427 14240
rect 5644 14182 6427 14184
rect 5644 14180 5650 14182
rect 6361 14179 6427 14182
rect 3442 14176 3762 14177
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3762 14176
rect 3442 14111 3762 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 13437 14176 13757 14177
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 14111 13757 14112
rect 3417 13970 3483 13973
rect 3785 13970 3851 13973
rect 11513 13970 11579 13973
rect 3417 13968 11579 13970
rect 3417 13912 3422 13968
rect 3478 13912 3790 13968
rect 3846 13912 11518 13968
rect 11574 13912 11579 13968
rect 3417 13910 11579 13912
rect 3417 13907 3483 13910
rect 3785 13907 3851 13910
rect 11513 13907 11579 13910
rect 15377 13970 15443 13973
rect 16400 13970 17200 14000
rect 15377 13968 17200 13970
rect 15377 13912 15382 13968
rect 15438 13912 17200 13968
rect 15377 13910 17200 13912
rect 15377 13907 15443 13910
rect 16400 13880 17200 13910
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 8385 13834 8451 13837
rect 9305 13834 9371 13837
rect 8385 13832 9371 13834
rect 8385 13776 8390 13832
rect 8446 13776 9310 13832
rect 9366 13776 9371 13832
rect 8385 13774 9371 13776
rect 8385 13771 8451 13774
rect 9305 13771 9371 13774
rect 5941 13632 6261 13633
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 13567 6261 13568
rect 10938 13632 11258 13633
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11258 13632
rect 10938 13567 11258 13568
rect 3969 13426 4035 13429
rect 10041 13426 10107 13429
rect 11513 13428 11579 13429
rect 11462 13426 11468 13428
rect 3969 13424 10107 13426
rect 3969 13368 3974 13424
rect 4030 13368 10046 13424
rect 10102 13368 10107 13424
rect 3969 13366 10107 13368
rect 11422 13366 11468 13426
rect 11532 13424 11579 13428
rect 11574 13368 11579 13424
rect 3969 13363 4035 13366
rect 10041 13363 10107 13366
rect 11462 13364 11468 13366
rect 11532 13364 11579 13368
rect 11513 13363 11579 13364
rect 12525 13426 12591 13429
rect 12709 13426 12775 13429
rect 12525 13424 12775 13426
rect 12525 13368 12530 13424
rect 12586 13368 12714 13424
rect 12770 13368 12775 13424
rect 12525 13366 12775 13368
rect 12525 13363 12591 13366
rect 12709 13363 12775 13366
rect 4521 13290 4587 13293
rect 11513 13290 11579 13293
rect 12525 13290 12591 13293
rect 4521 13288 8954 13290
rect 4521 13232 4526 13288
rect 4582 13232 8954 13288
rect 4521 13230 8954 13232
rect 4521 13227 4587 13230
rect 8894 13154 8954 13230
rect 11513 13288 12591 13290
rect 11513 13232 11518 13288
rect 11574 13232 12530 13288
rect 12586 13232 12591 13288
rect 11513 13230 12591 13232
rect 11513 13227 11579 13230
rect 12525 13227 12591 13230
rect 9857 13154 9923 13157
rect 11421 13154 11487 13157
rect 8894 13152 11487 13154
rect 8894 13096 9862 13152
rect 9918 13096 11426 13152
rect 11482 13096 11487 13152
rect 8894 13094 11487 13096
rect 9857 13091 9923 13094
rect 11421 13091 11487 13094
rect 3442 13088 3762 13089
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3762 13088
rect 3442 13023 3762 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 13437 13088 13757 13089
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 13023 13757 13024
rect 8886 12956 8892 13020
rect 8956 13018 8962 13020
rect 9213 13018 9279 13021
rect 8956 13016 9279 13018
rect 8956 12960 9218 13016
rect 9274 12960 9279 13016
rect 8956 12958 9279 12960
rect 8956 12956 8962 12958
rect 9213 12955 9279 12958
rect 0 12882 800 12912
rect 1669 12882 1735 12885
rect 0 12880 1735 12882
rect 0 12824 1674 12880
rect 1730 12824 1735 12880
rect 0 12822 1735 12824
rect 0 12792 800 12822
rect 1669 12819 1735 12822
rect 5073 12882 5139 12885
rect 11513 12882 11579 12885
rect 5073 12880 11579 12882
rect 5073 12824 5078 12880
rect 5134 12824 11518 12880
rect 11574 12824 11579 12880
rect 5073 12822 11579 12824
rect 5073 12819 5139 12822
rect 11513 12819 11579 12822
rect 5206 12684 5212 12748
rect 5276 12746 5282 12748
rect 6269 12746 6335 12749
rect 5276 12744 6335 12746
rect 5276 12688 6274 12744
rect 6330 12688 6335 12744
rect 5276 12686 6335 12688
rect 5276 12684 5282 12686
rect 6269 12683 6335 12686
rect 9949 12746 10015 12749
rect 12893 12746 12959 12749
rect 9949 12744 12959 12746
rect 9949 12688 9954 12744
rect 10010 12688 12898 12744
rect 12954 12688 12959 12744
rect 9949 12686 12959 12688
rect 9949 12683 10015 12686
rect 12893 12683 12959 12686
rect 5941 12544 6261 12545
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 12479 6261 12480
rect 10938 12544 11258 12545
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11258 12544
rect 10938 12479 11258 12480
rect 3442 12000 3762 12001
rect 0 11930 800 11960
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3762 12000
rect 3442 11935 3762 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 13437 12000 13757 12001
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 11935 13757 11936
rect 1669 11930 1735 11933
rect 0 11928 1735 11930
rect 0 11872 1674 11928
rect 1730 11872 1735 11928
rect 0 11870 1735 11872
rect 0 11840 800 11870
rect 1669 11867 1735 11870
rect 9949 11794 10015 11797
rect 10593 11794 10659 11797
rect 12249 11794 12315 11797
rect 9949 11792 12315 11794
rect 9949 11736 9954 11792
rect 10010 11736 10598 11792
rect 10654 11736 12254 11792
rect 12310 11736 12315 11792
rect 9949 11734 12315 11736
rect 9949 11731 10015 11734
rect 10593 11731 10659 11734
rect 12249 11731 12315 11734
rect 5941 11456 6261 11457
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 11391 6261 11392
rect 10938 11456 11258 11457
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11258 11456
rect 10938 11391 11258 11392
rect 11513 11386 11579 11389
rect 11646 11386 11652 11388
rect 11513 11384 11652 11386
rect 11513 11328 11518 11384
rect 11574 11328 11652 11384
rect 11513 11326 11652 11328
rect 11513 11323 11579 11326
rect 11646 11324 11652 11326
rect 11716 11324 11722 11388
rect 11513 11252 11579 11253
rect 11462 11188 11468 11252
rect 11532 11250 11579 11252
rect 11532 11248 11624 11250
rect 11574 11192 11624 11248
rect 11532 11190 11624 11192
rect 11532 11188 11579 11190
rect 11513 11187 11579 11188
rect 0 10978 800 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 800 10918
rect 1669 10915 1735 10918
rect 3442 10912 3762 10913
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3762 10912
rect 3442 10847 3762 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 13437 10912 13757 10913
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 10847 13757 10848
rect 7833 10570 7899 10573
rect 8753 10570 8819 10573
rect 7833 10568 8819 10570
rect 7833 10512 7838 10568
rect 7894 10512 8758 10568
rect 8814 10512 8819 10568
rect 7833 10510 8819 10512
rect 7833 10507 7899 10510
rect 8753 10507 8819 10510
rect 5941 10368 6261 10369
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 10303 6261 10304
rect 10938 10368 11258 10369
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11258 10368
rect 10938 10303 11258 10304
rect 5165 10164 5231 10165
rect 5165 10162 5212 10164
rect 5120 10160 5212 10162
rect 5120 10104 5170 10160
rect 5120 10102 5212 10104
rect 5165 10100 5212 10102
rect 5276 10100 5282 10164
rect 5441 10162 5507 10165
rect 5574 10162 5580 10164
rect 5441 10160 5580 10162
rect 5441 10104 5446 10160
rect 5502 10104 5580 10160
rect 5441 10102 5580 10104
rect 5165 10099 5231 10100
rect 5441 10099 5507 10102
rect 5574 10100 5580 10102
rect 5644 10100 5650 10164
rect 0 10026 800 10056
rect 1669 10026 1735 10029
rect 0 10024 1735 10026
rect 0 9968 1674 10024
rect 1730 9968 1735 10024
rect 0 9966 1735 9968
rect 0 9936 800 9966
rect 1669 9963 1735 9966
rect 10593 9888 10659 9893
rect 10593 9832 10598 9888
rect 10654 9832 10659 9888
rect 10593 9827 10659 9832
rect 15009 9890 15075 9893
rect 16400 9890 17200 9920
rect 15009 9888 17200 9890
rect 15009 9832 15014 9888
rect 15070 9832 17200 9888
rect 15009 9830 17200 9832
rect 15009 9827 15075 9830
rect 3442 9824 3762 9825
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3762 9824
rect 3442 9759 3762 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 10596 9618 10656 9827
rect 13437 9824 13757 9825
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 16400 9800 17200 9830
rect 13437 9759 13757 9760
rect 10726 9618 10732 9620
rect 10596 9558 10732 9618
rect 10726 9556 10732 9558
rect 10796 9556 10802 9620
rect 5809 9482 5875 9485
rect 9213 9482 9279 9485
rect 11697 9482 11763 9485
rect 5809 9480 9279 9482
rect 5809 9424 5814 9480
rect 5870 9424 9218 9480
rect 9274 9424 9279 9480
rect 5809 9422 9279 9424
rect 5809 9419 5875 9422
rect 9213 9419 9279 9422
rect 9998 9480 11763 9482
rect 9998 9424 11702 9480
rect 11758 9424 11763 9480
rect 9998 9422 11763 9424
rect 9998 9349 10058 9422
rect 11697 9419 11763 9422
rect 9949 9344 10058 9349
rect 9949 9288 9954 9344
rect 10010 9288 10058 9344
rect 9949 9286 10058 9288
rect 9949 9283 10015 9286
rect 5941 9280 6261 9281
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 9215 6261 9216
rect 10938 9280 11258 9281
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11258 9280
rect 10938 9215 11258 9216
rect 0 9074 800 9104
rect 2773 9074 2839 9077
rect 0 9072 2839 9074
rect 0 9016 2778 9072
rect 2834 9016 2839 9072
rect 0 9014 2839 9016
rect 0 8984 800 9014
rect 2773 9011 2839 9014
rect 9121 9074 9187 9077
rect 9254 9074 9260 9076
rect 9121 9072 9260 9074
rect 9121 9016 9126 9072
rect 9182 9016 9260 9072
rect 9121 9014 9260 9016
rect 9121 9011 9187 9014
rect 9254 9012 9260 9014
rect 9324 9012 9330 9076
rect 10133 9074 10199 9077
rect 10869 9074 10935 9077
rect 10133 9072 10935 9074
rect 10133 9016 10138 9072
rect 10194 9016 10874 9072
rect 10930 9016 10935 9072
rect 10133 9014 10935 9016
rect 10133 9011 10199 9014
rect 10869 9011 10935 9014
rect 8937 8802 9003 8805
rect 9070 8802 9076 8804
rect 8937 8800 9076 8802
rect 8937 8744 8942 8800
rect 8998 8744 9076 8800
rect 8937 8742 9076 8744
rect 8937 8739 9003 8742
rect 9070 8740 9076 8742
rect 9140 8740 9146 8804
rect 3442 8736 3762 8737
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3762 8736
rect 3442 8671 3762 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 13437 8736 13757 8737
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 8671 13757 8672
rect 8477 8530 8543 8533
rect 8886 8530 8892 8532
rect 8477 8528 8892 8530
rect 8477 8472 8482 8528
rect 8538 8472 8892 8528
rect 8477 8470 8892 8472
rect 8477 8467 8543 8470
rect 8886 8468 8892 8470
rect 8956 8468 8962 8532
rect 5073 8394 5139 8397
rect 9581 8394 9647 8397
rect 5073 8392 9647 8394
rect 5073 8336 5078 8392
rect 5134 8336 9586 8392
rect 9642 8336 9647 8392
rect 5073 8334 9647 8336
rect 5073 8331 5139 8334
rect 9581 8331 9647 8334
rect 9438 8196 9444 8260
rect 9508 8258 9514 8260
rect 9581 8258 9647 8261
rect 9508 8256 9647 8258
rect 9508 8200 9586 8256
rect 9642 8200 9647 8256
rect 9508 8198 9647 8200
rect 9508 8196 9514 8198
rect 9581 8195 9647 8198
rect 5941 8192 6261 8193
rect 0 8122 800 8152
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 8127 6261 8128
rect 10938 8192 11258 8193
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11258 8192
rect 10938 8127 11258 8128
rect 1761 8122 1827 8125
rect 0 8120 1827 8122
rect 0 8064 1766 8120
rect 1822 8064 1827 8120
rect 0 8062 1827 8064
rect 0 8032 800 8062
rect 1761 8059 1827 8062
rect 8661 7986 8727 7989
rect 9213 7986 9279 7989
rect 11697 7986 11763 7989
rect 8661 7984 11763 7986
rect 8661 7928 8666 7984
rect 8722 7928 9218 7984
rect 9274 7928 11702 7984
rect 11758 7928 11763 7984
rect 8661 7926 11763 7928
rect 8661 7923 8727 7926
rect 9213 7923 9279 7926
rect 11697 7923 11763 7926
rect 7189 7850 7255 7853
rect 9581 7850 9647 7853
rect 7189 7848 9647 7850
rect 7189 7792 7194 7848
rect 7250 7792 9586 7848
rect 9642 7792 9647 7848
rect 7189 7790 9647 7792
rect 7189 7787 7255 7790
rect 9581 7787 9647 7790
rect 3442 7648 3762 7649
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3762 7648
rect 3442 7583 3762 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 13437 7648 13757 7649
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 7583 13757 7584
rect 9121 7578 9187 7581
rect 8940 7576 9187 7578
rect 8940 7520 9126 7576
rect 9182 7520 9187 7576
rect 8940 7518 9187 7520
rect 8940 7445 9000 7518
rect 9121 7515 9187 7518
rect 8937 7440 9003 7445
rect 8937 7384 8942 7440
rect 8998 7384 9003 7440
rect 8937 7379 9003 7384
rect 0 7170 800 7200
rect 1669 7170 1735 7173
rect 0 7168 1735 7170
rect 0 7112 1674 7168
rect 1730 7112 1735 7168
rect 0 7110 1735 7112
rect 0 7080 800 7110
rect 1669 7107 1735 7110
rect 8845 7170 8911 7173
rect 9029 7170 9095 7173
rect 8845 7168 9095 7170
rect 8845 7112 8850 7168
rect 8906 7112 9034 7168
rect 9090 7112 9095 7168
rect 8845 7110 9095 7112
rect 8845 7107 8911 7110
rect 9029 7107 9095 7110
rect 5941 7104 6261 7105
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 7039 6261 7040
rect 10938 7104 11258 7105
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11258 7104
rect 10938 7039 11258 7040
rect 10041 6898 10107 6901
rect 13353 6898 13419 6901
rect 10041 6896 13419 6898
rect 10041 6840 10046 6896
rect 10102 6840 13358 6896
rect 13414 6840 13419 6896
rect 10041 6838 13419 6840
rect 10041 6835 10107 6838
rect 13353 6835 13419 6838
rect 3442 6560 3762 6561
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3762 6560
rect 3442 6495 3762 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 13437 6560 13757 6561
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 6495 13757 6496
rect 0 6218 800 6248
rect 1761 6218 1827 6221
rect 0 6216 1827 6218
rect 0 6160 1766 6216
rect 1822 6160 1827 6216
rect 0 6158 1827 6160
rect 0 6128 800 6158
rect 1761 6155 1827 6158
rect 5941 6016 6261 6017
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 5951 6261 5952
rect 10938 6016 11258 6017
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11258 6016
rect 10938 5951 11258 5952
rect 14917 5946 14983 5949
rect 16400 5946 17200 5976
rect 14917 5944 17200 5946
rect 14917 5888 14922 5944
rect 14978 5888 17200 5944
rect 14917 5886 17200 5888
rect 14917 5883 14983 5886
rect 16400 5856 17200 5886
rect 2865 5810 2931 5813
rect 6729 5810 6795 5813
rect 7373 5810 7439 5813
rect 2865 5808 7439 5810
rect 2865 5752 2870 5808
rect 2926 5752 6734 5808
rect 6790 5752 7378 5808
rect 7434 5752 7439 5808
rect 2865 5750 7439 5752
rect 2865 5747 2931 5750
rect 6729 5747 6795 5750
rect 7373 5747 7439 5750
rect 3442 5472 3762 5473
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3762 5472
rect 3442 5407 3762 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 13437 5472 13757 5473
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 5407 13757 5408
rect 0 5266 800 5296
rect 2313 5266 2379 5269
rect 0 5264 2379 5266
rect 0 5208 2318 5264
rect 2374 5208 2379 5264
rect 0 5206 2379 5208
rect 0 5176 800 5206
rect 2313 5203 2379 5206
rect 9438 5204 9444 5268
rect 9508 5266 9514 5268
rect 9581 5266 9647 5269
rect 9508 5264 9647 5266
rect 9508 5208 9586 5264
rect 9642 5208 9647 5264
rect 9508 5206 9647 5208
rect 9508 5204 9514 5206
rect 9581 5203 9647 5206
rect 7741 5130 7807 5133
rect 8477 5130 8543 5133
rect 7741 5128 8543 5130
rect 7741 5072 7746 5128
rect 7802 5072 8482 5128
rect 8538 5072 8543 5128
rect 7741 5070 8543 5072
rect 7741 5067 7807 5070
rect 8477 5067 8543 5070
rect 5941 4928 6261 4929
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 4863 6261 4864
rect 10938 4928 11258 4929
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11258 4928
rect 10938 4863 11258 4864
rect 4705 4586 4771 4589
rect 5165 4586 5231 4589
rect 7741 4586 7807 4589
rect 4705 4584 7807 4586
rect 4705 4528 4710 4584
rect 4766 4528 5170 4584
rect 5226 4528 7746 4584
rect 7802 4528 7807 4584
rect 4705 4526 7807 4528
rect 4705 4523 4771 4526
rect 5165 4523 5231 4526
rect 7741 4523 7807 4526
rect 10041 4586 10107 4589
rect 15193 4586 15259 4589
rect 10041 4584 15259 4586
rect 10041 4528 10046 4584
rect 10102 4528 15198 4584
rect 15254 4528 15259 4584
rect 10041 4526 15259 4528
rect 10041 4523 10107 4526
rect 15193 4523 15259 4526
rect 10593 4450 10659 4453
rect 13261 4450 13327 4453
rect 10593 4448 13327 4450
rect 10593 4392 10598 4448
rect 10654 4392 13266 4448
rect 13322 4392 13327 4448
rect 10593 4390 13327 4392
rect 10593 4387 10659 4390
rect 13261 4387 13327 4390
rect 3442 4384 3762 4385
rect 0 4314 800 4344
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3762 4384
rect 3442 4319 3762 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 13437 4384 13757 4385
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 4319 13757 4320
rect 1669 4314 1735 4317
rect 0 4312 1735 4314
rect 0 4256 1674 4312
rect 1730 4256 1735 4312
rect 0 4254 1735 4256
rect 0 4224 800 4254
rect 1669 4251 1735 4254
rect 8937 4314 9003 4317
rect 9254 4314 9260 4316
rect 8937 4312 9260 4314
rect 8937 4256 8942 4312
rect 8998 4256 9260 4312
rect 8937 4254 9260 4256
rect 8937 4251 9003 4254
rect 9254 4252 9260 4254
rect 9324 4314 9330 4316
rect 9324 4254 12634 4314
rect 9324 4252 9330 4254
rect 7557 4178 7623 4181
rect 9121 4180 9187 4181
rect 9070 4178 9076 4180
rect 7557 4176 9076 4178
rect 9140 4178 9187 4180
rect 12574 4178 12634 4254
rect 13813 4178 13879 4181
rect 9140 4176 9232 4178
rect 7557 4120 7562 4176
rect 7618 4120 9076 4176
rect 9182 4120 9232 4176
rect 7557 4118 9076 4120
rect 7557 4115 7623 4118
rect 9070 4116 9076 4118
rect 9140 4118 9232 4120
rect 12574 4176 13879 4178
rect 12574 4120 13818 4176
rect 13874 4120 13879 4176
rect 12574 4118 13879 4120
rect 9140 4116 9187 4118
rect 9121 4115 9187 4116
rect 13813 4115 13879 4118
rect 7373 4042 7439 4045
rect 10869 4042 10935 4045
rect 7373 4040 10935 4042
rect 7373 3984 7378 4040
rect 7434 3984 10874 4040
rect 10930 3984 10935 4040
rect 7373 3982 10935 3984
rect 7373 3979 7439 3982
rect 10869 3979 10935 3982
rect 10317 3906 10383 3909
rect 10726 3906 10732 3908
rect 10317 3904 10732 3906
rect 10317 3848 10322 3904
rect 10378 3848 10732 3904
rect 10317 3846 10732 3848
rect 10317 3843 10383 3846
rect 10726 3844 10732 3846
rect 10796 3844 10802 3908
rect 5941 3840 6261 3841
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 3775 6261 3776
rect 10938 3840 11258 3841
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11258 3840
rect 10938 3775 11258 3776
rect 2037 3770 2103 3773
rect 5533 3770 5599 3773
rect 2037 3768 5599 3770
rect 2037 3712 2042 3768
rect 2098 3712 5538 3768
rect 5594 3712 5599 3768
rect 2037 3710 5599 3712
rect 2037 3707 2103 3710
rect 5533 3707 5599 3710
rect 6453 3770 6519 3773
rect 9121 3770 9187 3773
rect 6453 3768 9187 3770
rect 6453 3712 6458 3768
rect 6514 3712 9126 3768
rect 9182 3712 9187 3768
rect 6453 3710 9187 3712
rect 6453 3707 6519 3710
rect 9121 3707 9187 3710
rect 3969 3634 4035 3637
rect 11605 3634 11671 3637
rect 3969 3632 11671 3634
rect 3969 3576 3974 3632
rect 4030 3576 11610 3632
rect 11666 3576 11671 3632
rect 3969 3574 11671 3576
rect 3969 3571 4035 3574
rect 11605 3571 11671 3574
rect 12065 3634 12131 3637
rect 12985 3634 13051 3637
rect 12065 3632 13051 3634
rect 12065 3576 12070 3632
rect 12126 3576 12990 3632
rect 13046 3576 13051 3632
rect 12065 3574 13051 3576
rect 12065 3571 12131 3574
rect 12985 3571 13051 3574
rect 4981 3498 5047 3501
rect 10133 3498 10199 3501
rect 4981 3496 10199 3498
rect 4981 3440 4986 3496
rect 5042 3440 10138 3496
rect 10194 3440 10199 3496
rect 4981 3438 10199 3440
rect 4981 3435 5047 3438
rect 10133 3435 10199 3438
rect 0 3362 800 3392
rect 1669 3362 1735 3365
rect 0 3360 1735 3362
rect 0 3304 1674 3360
rect 1730 3304 1735 3360
rect 0 3302 1735 3304
rect 0 3272 800 3302
rect 1669 3299 1735 3302
rect 9673 3362 9739 3365
rect 10501 3362 10567 3365
rect 12249 3362 12315 3365
rect 9673 3360 12315 3362
rect 9673 3304 9678 3360
rect 9734 3304 10506 3360
rect 10562 3304 12254 3360
rect 12310 3304 12315 3360
rect 9673 3302 12315 3304
rect 9673 3299 9739 3302
rect 10501 3299 10567 3302
rect 12249 3299 12315 3302
rect 3442 3296 3762 3297
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3762 3296
rect 3442 3231 3762 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 13437 3296 13757 3297
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 13437 3231 13757 3232
rect 9949 3226 10015 3229
rect 12617 3226 12683 3229
rect 9949 3224 12683 3226
rect 9949 3168 9954 3224
rect 10010 3168 12622 3224
rect 12678 3168 12683 3224
rect 9949 3166 12683 3168
rect 9949 3163 10015 3166
rect 12617 3163 12683 3166
rect 1485 3090 1551 3093
rect 8845 3090 8911 3093
rect 1485 3088 8911 3090
rect 1485 3032 1490 3088
rect 1546 3032 8850 3088
rect 8906 3032 8911 3088
rect 1485 3030 8911 3032
rect 1485 3027 1551 3030
rect 8845 3027 8911 3030
rect 10225 3090 10291 3093
rect 11973 3090 12039 3093
rect 10225 3088 12039 3090
rect 10225 3032 10230 3088
rect 10286 3032 11978 3088
rect 12034 3032 12039 3088
rect 10225 3030 12039 3032
rect 10225 3027 10291 3030
rect 11973 3027 12039 3030
rect 4797 2954 4863 2957
rect 12065 2954 12131 2957
rect 4797 2952 12131 2954
rect 4797 2896 4802 2952
rect 4858 2896 12070 2952
rect 12126 2896 12131 2952
rect 4797 2894 12131 2896
rect 4797 2891 4863 2894
rect 12065 2891 12131 2894
rect 6361 2818 6427 2821
rect 9765 2818 9831 2821
rect 10041 2818 10107 2821
rect 6361 2816 10107 2818
rect 6361 2760 6366 2816
rect 6422 2760 9770 2816
rect 9826 2760 10046 2816
rect 10102 2760 10107 2816
rect 6361 2758 10107 2760
rect 6361 2755 6427 2758
rect 9765 2755 9831 2758
rect 10041 2755 10107 2758
rect 5941 2752 6261 2753
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2687 6261 2688
rect 10938 2752 11258 2753
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11258 2752
rect 10938 2687 11258 2688
rect 0 2410 800 2440
rect 4981 2410 5047 2413
rect 0 2408 5047 2410
rect 0 2352 4986 2408
rect 5042 2352 5047 2408
rect 0 2350 5047 2352
rect 0 2320 800 2350
rect 4981 2347 5047 2350
rect 3442 2208 3762 2209
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3762 2208
rect 3442 2143 3762 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 13437 2208 13757 2209
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2143 13757 2144
rect 15009 2002 15075 2005
rect 16400 2002 17200 2032
rect 15009 2000 17200 2002
rect 15009 1944 15014 2000
rect 15070 1944 17200 2000
rect 15009 1942 17200 1944
rect 15009 1939 15075 1942
rect 16400 1912 17200 1942
rect 0 1458 800 1488
rect 2037 1458 2103 1461
rect 0 1456 2103 1458
rect 0 1400 2042 1456
rect 2098 1400 2103 1456
rect 0 1398 2103 1400
rect 0 1368 800 1398
rect 2037 1395 2103 1398
rect 0 506 800 536
rect 2957 506 3023 509
rect 0 504 3023 506
rect 0 448 2962 504
rect 3018 448 3023 504
rect 0 446 3023 448
rect 0 416 800 446
rect 2957 443 3023 446
<< via3 >>
rect 3450 17436 3514 17440
rect 3450 17380 3454 17436
rect 3454 17380 3510 17436
rect 3510 17380 3514 17436
rect 3450 17376 3514 17380
rect 3530 17436 3594 17440
rect 3530 17380 3534 17436
rect 3534 17380 3590 17436
rect 3590 17380 3594 17436
rect 3530 17376 3594 17380
rect 3610 17436 3674 17440
rect 3610 17380 3614 17436
rect 3614 17380 3670 17436
rect 3670 17380 3674 17436
rect 3610 17376 3674 17380
rect 3690 17436 3754 17440
rect 3690 17380 3694 17436
rect 3694 17380 3750 17436
rect 3750 17380 3754 17436
rect 3690 17376 3754 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 13445 17436 13509 17440
rect 13445 17380 13449 17436
rect 13449 17380 13505 17436
rect 13505 17380 13509 17436
rect 13445 17376 13509 17380
rect 13525 17436 13589 17440
rect 13525 17380 13529 17436
rect 13529 17380 13585 17436
rect 13585 17380 13589 17436
rect 13525 17376 13589 17380
rect 13605 17436 13669 17440
rect 13605 17380 13609 17436
rect 13609 17380 13665 17436
rect 13665 17380 13669 17436
rect 13605 17376 13669 17380
rect 13685 17436 13749 17440
rect 13685 17380 13689 17436
rect 13689 17380 13745 17436
rect 13745 17380 13749 17436
rect 13685 17376 13749 17380
rect 11652 17172 11716 17236
rect 5949 16892 6013 16896
rect 5949 16836 5953 16892
rect 5953 16836 6009 16892
rect 6009 16836 6013 16892
rect 5949 16832 6013 16836
rect 6029 16892 6093 16896
rect 6029 16836 6033 16892
rect 6033 16836 6089 16892
rect 6089 16836 6093 16892
rect 6029 16832 6093 16836
rect 6109 16892 6173 16896
rect 6109 16836 6113 16892
rect 6113 16836 6169 16892
rect 6169 16836 6173 16892
rect 6109 16832 6173 16836
rect 6189 16892 6253 16896
rect 6189 16836 6193 16892
rect 6193 16836 6249 16892
rect 6249 16836 6253 16892
rect 6189 16832 6253 16836
rect 10946 16892 11010 16896
rect 10946 16836 10950 16892
rect 10950 16836 11006 16892
rect 11006 16836 11010 16892
rect 10946 16832 11010 16836
rect 11026 16892 11090 16896
rect 11026 16836 11030 16892
rect 11030 16836 11086 16892
rect 11086 16836 11090 16892
rect 11026 16832 11090 16836
rect 11106 16892 11170 16896
rect 11106 16836 11110 16892
rect 11110 16836 11166 16892
rect 11166 16836 11170 16892
rect 11106 16832 11170 16836
rect 11186 16892 11250 16896
rect 11186 16836 11190 16892
rect 11190 16836 11246 16892
rect 11246 16836 11250 16892
rect 11186 16832 11250 16836
rect 3450 16348 3514 16352
rect 3450 16292 3454 16348
rect 3454 16292 3510 16348
rect 3510 16292 3514 16348
rect 3450 16288 3514 16292
rect 3530 16348 3594 16352
rect 3530 16292 3534 16348
rect 3534 16292 3590 16348
rect 3590 16292 3594 16348
rect 3530 16288 3594 16292
rect 3610 16348 3674 16352
rect 3610 16292 3614 16348
rect 3614 16292 3670 16348
rect 3670 16292 3674 16348
rect 3610 16288 3674 16292
rect 3690 16348 3754 16352
rect 3690 16292 3694 16348
rect 3694 16292 3750 16348
rect 3750 16292 3754 16348
rect 3690 16288 3754 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 13445 16348 13509 16352
rect 13445 16292 13449 16348
rect 13449 16292 13505 16348
rect 13505 16292 13509 16348
rect 13445 16288 13509 16292
rect 13525 16348 13589 16352
rect 13525 16292 13529 16348
rect 13529 16292 13585 16348
rect 13585 16292 13589 16348
rect 13525 16288 13589 16292
rect 13605 16348 13669 16352
rect 13605 16292 13609 16348
rect 13609 16292 13665 16348
rect 13665 16292 13669 16348
rect 13605 16288 13669 16292
rect 13685 16348 13749 16352
rect 13685 16292 13689 16348
rect 13689 16292 13745 16348
rect 13745 16292 13749 16348
rect 13685 16288 13749 16292
rect 5949 15804 6013 15808
rect 5949 15748 5953 15804
rect 5953 15748 6009 15804
rect 6009 15748 6013 15804
rect 5949 15744 6013 15748
rect 6029 15804 6093 15808
rect 6029 15748 6033 15804
rect 6033 15748 6089 15804
rect 6089 15748 6093 15804
rect 6029 15744 6093 15748
rect 6109 15804 6173 15808
rect 6109 15748 6113 15804
rect 6113 15748 6169 15804
rect 6169 15748 6173 15804
rect 6109 15744 6173 15748
rect 6189 15804 6253 15808
rect 6189 15748 6193 15804
rect 6193 15748 6249 15804
rect 6249 15748 6253 15804
rect 6189 15744 6253 15748
rect 10946 15804 11010 15808
rect 10946 15748 10950 15804
rect 10950 15748 11006 15804
rect 11006 15748 11010 15804
rect 10946 15744 11010 15748
rect 11026 15804 11090 15808
rect 11026 15748 11030 15804
rect 11030 15748 11086 15804
rect 11086 15748 11090 15804
rect 11026 15744 11090 15748
rect 11106 15804 11170 15808
rect 11106 15748 11110 15804
rect 11110 15748 11166 15804
rect 11166 15748 11170 15804
rect 11106 15744 11170 15748
rect 11186 15804 11250 15808
rect 11186 15748 11190 15804
rect 11190 15748 11246 15804
rect 11246 15748 11250 15804
rect 11186 15744 11250 15748
rect 3450 15260 3514 15264
rect 3450 15204 3454 15260
rect 3454 15204 3510 15260
rect 3510 15204 3514 15260
rect 3450 15200 3514 15204
rect 3530 15260 3594 15264
rect 3530 15204 3534 15260
rect 3534 15204 3590 15260
rect 3590 15204 3594 15260
rect 3530 15200 3594 15204
rect 3610 15260 3674 15264
rect 3610 15204 3614 15260
rect 3614 15204 3670 15260
rect 3670 15204 3674 15260
rect 3610 15200 3674 15204
rect 3690 15260 3754 15264
rect 3690 15204 3694 15260
rect 3694 15204 3750 15260
rect 3750 15204 3754 15260
rect 3690 15200 3754 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 8892 14860 8956 14924
rect 13445 15260 13509 15264
rect 13445 15204 13449 15260
rect 13449 15204 13505 15260
rect 13505 15204 13509 15260
rect 13445 15200 13509 15204
rect 13525 15260 13589 15264
rect 13525 15204 13529 15260
rect 13529 15204 13585 15260
rect 13585 15204 13589 15260
rect 13525 15200 13589 15204
rect 13605 15260 13669 15264
rect 13605 15204 13609 15260
rect 13609 15204 13665 15260
rect 13665 15204 13669 15260
rect 13605 15200 13669 15204
rect 13685 15260 13749 15264
rect 13685 15204 13689 15260
rect 13689 15204 13745 15260
rect 13745 15204 13749 15260
rect 13685 15200 13749 15204
rect 5949 14716 6013 14720
rect 5949 14660 5953 14716
rect 5953 14660 6009 14716
rect 6009 14660 6013 14716
rect 5949 14656 6013 14660
rect 6029 14716 6093 14720
rect 6029 14660 6033 14716
rect 6033 14660 6089 14716
rect 6089 14660 6093 14716
rect 6029 14656 6093 14660
rect 6109 14716 6173 14720
rect 6109 14660 6113 14716
rect 6113 14660 6169 14716
rect 6169 14660 6173 14716
rect 6109 14656 6173 14660
rect 6189 14716 6253 14720
rect 6189 14660 6193 14716
rect 6193 14660 6249 14716
rect 6249 14660 6253 14716
rect 6189 14656 6253 14660
rect 10946 14716 11010 14720
rect 10946 14660 10950 14716
rect 10950 14660 11006 14716
rect 11006 14660 11010 14716
rect 10946 14656 11010 14660
rect 11026 14716 11090 14720
rect 11026 14660 11030 14716
rect 11030 14660 11086 14716
rect 11086 14660 11090 14716
rect 11026 14656 11090 14660
rect 11106 14716 11170 14720
rect 11106 14660 11110 14716
rect 11110 14660 11166 14716
rect 11166 14660 11170 14716
rect 11106 14656 11170 14660
rect 11186 14716 11250 14720
rect 11186 14660 11190 14716
rect 11190 14660 11246 14716
rect 11246 14660 11250 14716
rect 11186 14656 11250 14660
rect 5580 14180 5644 14244
rect 3450 14172 3514 14176
rect 3450 14116 3454 14172
rect 3454 14116 3510 14172
rect 3510 14116 3514 14172
rect 3450 14112 3514 14116
rect 3530 14172 3594 14176
rect 3530 14116 3534 14172
rect 3534 14116 3590 14172
rect 3590 14116 3594 14172
rect 3530 14112 3594 14116
rect 3610 14172 3674 14176
rect 3610 14116 3614 14172
rect 3614 14116 3670 14172
rect 3670 14116 3674 14172
rect 3610 14112 3674 14116
rect 3690 14172 3754 14176
rect 3690 14116 3694 14172
rect 3694 14116 3750 14172
rect 3750 14116 3754 14172
rect 3690 14112 3754 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 13445 14172 13509 14176
rect 13445 14116 13449 14172
rect 13449 14116 13505 14172
rect 13505 14116 13509 14172
rect 13445 14112 13509 14116
rect 13525 14172 13589 14176
rect 13525 14116 13529 14172
rect 13529 14116 13585 14172
rect 13585 14116 13589 14172
rect 13525 14112 13589 14116
rect 13605 14172 13669 14176
rect 13605 14116 13609 14172
rect 13609 14116 13665 14172
rect 13665 14116 13669 14172
rect 13605 14112 13669 14116
rect 13685 14172 13749 14176
rect 13685 14116 13689 14172
rect 13689 14116 13745 14172
rect 13745 14116 13749 14172
rect 13685 14112 13749 14116
rect 5949 13628 6013 13632
rect 5949 13572 5953 13628
rect 5953 13572 6009 13628
rect 6009 13572 6013 13628
rect 5949 13568 6013 13572
rect 6029 13628 6093 13632
rect 6029 13572 6033 13628
rect 6033 13572 6089 13628
rect 6089 13572 6093 13628
rect 6029 13568 6093 13572
rect 6109 13628 6173 13632
rect 6109 13572 6113 13628
rect 6113 13572 6169 13628
rect 6169 13572 6173 13628
rect 6109 13568 6173 13572
rect 6189 13628 6253 13632
rect 6189 13572 6193 13628
rect 6193 13572 6249 13628
rect 6249 13572 6253 13628
rect 6189 13568 6253 13572
rect 10946 13628 11010 13632
rect 10946 13572 10950 13628
rect 10950 13572 11006 13628
rect 11006 13572 11010 13628
rect 10946 13568 11010 13572
rect 11026 13628 11090 13632
rect 11026 13572 11030 13628
rect 11030 13572 11086 13628
rect 11086 13572 11090 13628
rect 11026 13568 11090 13572
rect 11106 13628 11170 13632
rect 11106 13572 11110 13628
rect 11110 13572 11166 13628
rect 11166 13572 11170 13628
rect 11106 13568 11170 13572
rect 11186 13628 11250 13632
rect 11186 13572 11190 13628
rect 11190 13572 11246 13628
rect 11246 13572 11250 13628
rect 11186 13568 11250 13572
rect 11468 13424 11532 13428
rect 11468 13368 11518 13424
rect 11518 13368 11532 13424
rect 11468 13364 11532 13368
rect 3450 13084 3514 13088
rect 3450 13028 3454 13084
rect 3454 13028 3510 13084
rect 3510 13028 3514 13084
rect 3450 13024 3514 13028
rect 3530 13084 3594 13088
rect 3530 13028 3534 13084
rect 3534 13028 3590 13084
rect 3590 13028 3594 13084
rect 3530 13024 3594 13028
rect 3610 13084 3674 13088
rect 3610 13028 3614 13084
rect 3614 13028 3670 13084
rect 3670 13028 3674 13084
rect 3610 13024 3674 13028
rect 3690 13084 3754 13088
rect 3690 13028 3694 13084
rect 3694 13028 3750 13084
rect 3750 13028 3754 13084
rect 3690 13024 3754 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 13445 13084 13509 13088
rect 13445 13028 13449 13084
rect 13449 13028 13505 13084
rect 13505 13028 13509 13084
rect 13445 13024 13509 13028
rect 13525 13084 13589 13088
rect 13525 13028 13529 13084
rect 13529 13028 13585 13084
rect 13585 13028 13589 13084
rect 13525 13024 13589 13028
rect 13605 13084 13669 13088
rect 13605 13028 13609 13084
rect 13609 13028 13665 13084
rect 13665 13028 13669 13084
rect 13605 13024 13669 13028
rect 13685 13084 13749 13088
rect 13685 13028 13689 13084
rect 13689 13028 13745 13084
rect 13745 13028 13749 13084
rect 13685 13024 13749 13028
rect 8892 12956 8956 13020
rect 5212 12684 5276 12748
rect 5949 12540 6013 12544
rect 5949 12484 5953 12540
rect 5953 12484 6009 12540
rect 6009 12484 6013 12540
rect 5949 12480 6013 12484
rect 6029 12540 6093 12544
rect 6029 12484 6033 12540
rect 6033 12484 6089 12540
rect 6089 12484 6093 12540
rect 6029 12480 6093 12484
rect 6109 12540 6173 12544
rect 6109 12484 6113 12540
rect 6113 12484 6169 12540
rect 6169 12484 6173 12540
rect 6109 12480 6173 12484
rect 6189 12540 6253 12544
rect 6189 12484 6193 12540
rect 6193 12484 6249 12540
rect 6249 12484 6253 12540
rect 6189 12480 6253 12484
rect 10946 12540 11010 12544
rect 10946 12484 10950 12540
rect 10950 12484 11006 12540
rect 11006 12484 11010 12540
rect 10946 12480 11010 12484
rect 11026 12540 11090 12544
rect 11026 12484 11030 12540
rect 11030 12484 11086 12540
rect 11086 12484 11090 12540
rect 11026 12480 11090 12484
rect 11106 12540 11170 12544
rect 11106 12484 11110 12540
rect 11110 12484 11166 12540
rect 11166 12484 11170 12540
rect 11106 12480 11170 12484
rect 11186 12540 11250 12544
rect 11186 12484 11190 12540
rect 11190 12484 11246 12540
rect 11246 12484 11250 12540
rect 11186 12480 11250 12484
rect 3450 11996 3514 12000
rect 3450 11940 3454 11996
rect 3454 11940 3510 11996
rect 3510 11940 3514 11996
rect 3450 11936 3514 11940
rect 3530 11996 3594 12000
rect 3530 11940 3534 11996
rect 3534 11940 3590 11996
rect 3590 11940 3594 11996
rect 3530 11936 3594 11940
rect 3610 11996 3674 12000
rect 3610 11940 3614 11996
rect 3614 11940 3670 11996
rect 3670 11940 3674 11996
rect 3610 11936 3674 11940
rect 3690 11996 3754 12000
rect 3690 11940 3694 11996
rect 3694 11940 3750 11996
rect 3750 11940 3754 11996
rect 3690 11936 3754 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 13445 11996 13509 12000
rect 13445 11940 13449 11996
rect 13449 11940 13505 11996
rect 13505 11940 13509 11996
rect 13445 11936 13509 11940
rect 13525 11996 13589 12000
rect 13525 11940 13529 11996
rect 13529 11940 13585 11996
rect 13585 11940 13589 11996
rect 13525 11936 13589 11940
rect 13605 11996 13669 12000
rect 13605 11940 13609 11996
rect 13609 11940 13665 11996
rect 13665 11940 13669 11996
rect 13605 11936 13669 11940
rect 13685 11996 13749 12000
rect 13685 11940 13689 11996
rect 13689 11940 13745 11996
rect 13745 11940 13749 11996
rect 13685 11936 13749 11940
rect 5949 11452 6013 11456
rect 5949 11396 5953 11452
rect 5953 11396 6009 11452
rect 6009 11396 6013 11452
rect 5949 11392 6013 11396
rect 6029 11452 6093 11456
rect 6029 11396 6033 11452
rect 6033 11396 6089 11452
rect 6089 11396 6093 11452
rect 6029 11392 6093 11396
rect 6109 11452 6173 11456
rect 6109 11396 6113 11452
rect 6113 11396 6169 11452
rect 6169 11396 6173 11452
rect 6109 11392 6173 11396
rect 6189 11452 6253 11456
rect 6189 11396 6193 11452
rect 6193 11396 6249 11452
rect 6249 11396 6253 11452
rect 6189 11392 6253 11396
rect 10946 11452 11010 11456
rect 10946 11396 10950 11452
rect 10950 11396 11006 11452
rect 11006 11396 11010 11452
rect 10946 11392 11010 11396
rect 11026 11452 11090 11456
rect 11026 11396 11030 11452
rect 11030 11396 11086 11452
rect 11086 11396 11090 11452
rect 11026 11392 11090 11396
rect 11106 11452 11170 11456
rect 11106 11396 11110 11452
rect 11110 11396 11166 11452
rect 11166 11396 11170 11452
rect 11106 11392 11170 11396
rect 11186 11452 11250 11456
rect 11186 11396 11190 11452
rect 11190 11396 11246 11452
rect 11246 11396 11250 11452
rect 11186 11392 11250 11396
rect 11652 11324 11716 11388
rect 11468 11248 11532 11252
rect 11468 11192 11518 11248
rect 11518 11192 11532 11248
rect 11468 11188 11532 11192
rect 3450 10908 3514 10912
rect 3450 10852 3454 10908
rect 3454 10852 3510 10908
rect 3510 10852 3514 10908
rect 3450 10848 3514 10852
rect 3530 10908 3594 10912
rect 3530 10852 3534 10908
rect 3534 10852 3590 10908
rect 3590 10852 3594 10908
rect 3530 10848 3594 10852
rect 3610 10908 3674 10912
rect 3610 10852 3614 10908
rect 3614 10852 3670 10908
rect 3670 10852 3674 10908
rect 3610 10848 3674 10852
rect 3690 10908 3754 10912
rect 3690 10852 3694 10908
rect 3694 10852 3750 10908
rect 3750 10852 3754 10908
rect 3690 10848 3754 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 13445 10908 13509 10912
rect 13445 10852 13449 10908
rect 13449 10852 13505 10908
rect 13505 10852 13509 10908
rect 13445 10848 13509 10852
rect 13525 10908 13589 10912
rect 13525 10852 13529 10908
rect 13529 10852 13585 10908
rect 13585 10852 13589 10908
rect 13525 10848 13589 10852
rect 13605 10908 13669 10912
rect 13605 10852 13609 10908
rect 13609 10852 13665 10908
rect 13665 10852 13669 10908
rect 13605 10848 13669 10852
rect 13685 10908 13749 10912
rect 13685 10852 13689 10908
rect 13689 10852 13745 10908
rect 13745 10852 13749 10908
rect 13685 10848 13749 10852
rect 5949 10364 6013 10368
rect 5949 10308 5953 10364
rect 5953 10308 6009 10364
rect 6009 10308 6013 10364
rect 5949 10304 6013 10308
rect 6029 10364 6093 10368
rect 6029 10308 6033 10364
rect 6033 10308 6089 10364
rect 6089 10308 6093 10364
rect 6029 10304 6093 10308
rect 6109 10364 6173 10368
rect 6109 10308 6113 10364
rect 6113 10308 6169 10364
rect 6169 10308 6173 10364
rect 6109 10304 6173 10308
rect 6189 10364 6253 10368
rect 6189 10308 6193 10364
rect 6193 10308 6249 10364
rect 6249 10308 6253 10364
rect 6189 10304 6253 10308
rect 10946 10364 11010 10368
rect 10946 10308 10950 10364
rect 10950 10308 11006 10364
rect 11006 10308 11010 10364
rect 10946 10304 11010 10308
rect 11026 10364 11090 10368
rect 11026 10308 11030 10364
rect 11030 10308 11086 10364
rect 11086 10308 11090 10364
rect 11026 10304 11090 10308
rect 11106 10364 11170 10368
rect 11106 10308 11110 10364
rect 11110 10308 11166 10364
rect 11166 10308 11170 10364
rect 11106 10304 11170 10308
rect 11186 10364 11250 10368
rect 11186 10308 11190 10364
rect 11190 10308 11246 10364
rect 11246 10308 11250 10364
rect 11186 10304 11250 10308
rect 5212 10160 5276 10164
rect 5212 10104 5226 10160
rect 5226 10104 5276 10160
rect 5212 10100 5276 10104
rect 5580 10100 5644 10164
rect 3450 9820 3514 9824
rect 3450 9764 3454 9820
rect 3454 9764 3510 9820
rect 3510 9764 3514 9820
rect 3450 9760 3514 9764
rect 3530 9820 3594 9824
rect 3530 9764 3534 9820
rect 3534 9764 3590 9820
rect 3590 9764 3594 9820
rect 3530 9760 3594 9764
rect 3610 9820 3674 9824
rect 3610 9764 3614 9820
rect 3614 9764 3670 9820
rect 3670 9764 3674 9820
rect 3610 9760 3674 9764
rect 3690 9820 3754 9824
rect 3690 9764 3694 9820
rect 3694 9764 3750 9820
rect 3750 9764 3754 9820
rect 3690 9760 3754 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 13445 9820 13509 9824
rect 13445 9764 13449 9820
rect 13449 9764 13505 9820
rect 13505 9764 13509 9820
rect 13445 9760 13509 9764
rect 13525 9820 13589 9824
rect 13525 9764 13529 9820
rect 13529 9764 13585 9820
rect 13585 9764 13589 9820
rect 13525 9760 13589 9764
rect 13605 9820 13669 9824
rect 13605 9764 13609 9820
rect 13609 9764 13665 9820
rect 13665 9764 13669 9820
rect 13605 9760 13669 9764
rect 13685 9820 13749 9824
rect 13685 9764 13689 9820
rect 13689 9764 13745 9820
rect 13745 9764 13749 9820
rect 13685 9760 13749 9764
rect 10732 9556 10796 9620
rect 5949 9276 6013 9280
rect 5949 9220 5953 9276
rect 5953 9220 6009 9276
rect 6009 9220 6013 9276
rect 5949 9216 6013 9220
rect 6029 9276 6093 9280
rect 6029 9220 6033 9276
rect 6033 9220 6089 9276
rect 6089 9220 6093 9276
rect 6029 9216 6093 9220
rect 6109 9276 6173 9280
rect 6109 9220 6113 9276
rect 6113 9220 6169 9276
rect 6169 9220 6173 9276
rect 6109 9216 6173 9220
rect 6189 9276 6253 9280
rect 6189 9220 6193 9276
rect 6193 9220 6249 9276
rect 6249 9220 6253 9276
rect 6189 9216 6253 9220
rect 10946 9276 11010 9280
rect 10946 9220 10950 9276
rect 10950 9220 11006 9276
rect 11006 9220 11010 9276
rect 10946 9216 11010 9220
rect 11026 9276 11090 9280
rect 11026 9220 11030 9276
rect 11030 9220 11086 9276
rect 11086 9220 11090 9276
rect 11026 9216 11090 9220
rect 11106 9276 11170 9280
rect 11106 9220 11110 9276
rect 11110 9220 11166 9276
rect 11166 9220 11170 9276
rect 11106 9216 11170 9220
rect 11186 9276 11250 9280
rect 11186 9220 11190 9276
rect 11190 9220 11246 9276
rect 11246 9220 11250 9276
rect 11186 9216 11250 9220
rect 9260 9012 9324 9076
rect 9076 8740 9140 8804
rect 3450 8732 3514 8736
rect 3450 8676 3454 8732
rect 3454 8676 3510 8732
rect 3510 8676 3514 8732
rect 3450 8672 3514 8676
rect 3530 8732 3594 8736
rect 3530 8676 3534 8732
rect 3534 8676 3590 8732
rect 3590 8676 3594 8732
rect 3530 8672 3594 8676
rect 3610 8732 3674 8736
rect 3610 8676 3614 8732
rect 3614 8676 3670 8732
rect 3670 8676 3674 8732
rect 3610 8672 3674 8676
rect 3690 8732 3754 8736
rect 3690 8676 3694 8732
rect 3694 8676 3750 8732
rect 3750 8676 3754 8732
rect 3690 8672 3754 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 13445 8732 13509 8736
rect 13445 8676 13449 8732
rect 13449 8676 13505 8732
rect 13505 8676 13509 8732
rect 13445 8672 13509 8676
rect 13525 8732 13589 8736
rect 13525 8676 13529 8732
rect 13529 8676 13585 8732
rect 13585 8676 13589 8732
rect 13525 8672 13589 8676
rect 13605 8732 13669 8736
rect 13605 8676 13609 8732
rect 13609 8676 13665 8732
rect 13665 8676 13669 8732
rect 13605 8672 13669 8676
rect 13685 8732 13749 8736
rect 13685 8676 13689 8732
rect 13689 8676 13745 8732
rect 13745 8676 13749 8732
rect 13685 8672 13749 8676
rect 8892 8468 8956 8532
rect 9444 8196 9508 8260
rect 5949 8188 6013 8192
rect 5949 8132 5953 8188
rect 5953 8132 6009 8188
rect 6009 8132 6013 8188
rect 5949 8128 6013 8132
rect 6029 8188 6093 8192
rect 6029 8132 6033 8188
rect 6033 8132 6089 8188
rect 6089 8132 6093 8188
rect 6029 8128 6093 8132
rect 6109 8188 6173 8192
rect 6109 8132 6113 8188
rect 6113 8132 6169 8188
rect 6169 8132 6173 8188
rect 6109 8128 6173 8132
rect 6189 8188 6253 8192
rect 6189 8132 6193 8188
rect 6193 8132 6249 8188
rect 6249 8132 6253 8188
rect 6189 8128 6253 8132
rect 10946 8188 11010 8192
rect 10946 8132 10950 8188
rect 10950 8132 11006 8188
rect 11006 8132 11010 8188
rect 10946 8128 11010 8132
rect 11026 8188 11090 8192
rect 11026 8132 11030 8188
rect 11030 8132 11086 8188
rect 11086 8132 11090 8188
rect 11026 8128 11090 8132
rect 11106 8188 11170 8192
rect 11106 8132 11110 8188
rect 11110 8132 11166 8188
rect 11166 8132 11170 8188
rect 11106 8128 11170 8132
rect 11186 8188 11250 8192
rect 11186 8132 11190 8188
rect 11190 8132 11246 8188
rect 11246 8132 11250 8188
rect 11186 8128 11250 8132
rect 3450 7644 3514 7648
rect 3450 7588 3454 7644
rect 3454 7588 3510 7644
rect 3510 7588 3514 7644
rect 3450 7584 3514 7588
rect 3530 7644 3594 7648
rect 3530 7588 3534 7644
rect 3534 7588 3590 7644
rect 3590 7588 3594 7644
rect 3530 7584 3594 7588
rect 3610 7644 3674 7648
rect 3610 7588 3614 7644
rect 3614 7588 3670 7644
rect 3670 7588 3674 7644
rect 3610 7584 3674 7588
rect 3690 7644 3754 7648
rect 3690 7588 3694 7644
rect 3694 7588 3750 7644
rect 3750 7588 3754 7644
rect 3690 7584 3754 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 13445 7644 13509 7648
rect 13445 7588 13449 7644
rect 13449 7588 13505 7644
rect 13505 7588 13509 7644
rect 13445 7584 13509 7588
rect 13525 7644 13589 7648
rect 13525 7588 13529 7644
rect 13529 7588 13585 7644
rect 13585 7588 13589 7644
rect 13525 7584 13589 7588
rect 13605 7644 13669 7648
rect 13605 7588 13609 7644
rect 13609 7588 13665 7644
rect 13665 7588 13669 7644
rect 13605 7584 13669 7588
rect 13685 7644 13749 7648
rect 13685 7588 13689 7644
rect 13689 7588 13745 7644
rect 13745 7588 13749 7644
rect 13685 7584 13749 7588
rect 5949 7100 6013 7104
rect 5949 7044 5953 7100
rect 5953 7044 6009 7100
rect 6009 7044 6013 7100
rect 5949 7040 6013 7044
rect 6029 7100 6093 7104
rect 6029 7044 6033 7100
rect 6033 7044 6089 7100
rect 6089 7044 6093 7100
rect 6029 7040 6093 7044
rect 6109 7100 6173 7104
rect 6109 7044 6113 7100
rect 6113 7044 6169 7100
rect 6169 7044 6173 7100
rect 6109 7040 6173 7044
rect 6189 7100 6253 7104
rect 6189 7044 6193 7100
rect 6193 7044 6249 7100
rect 6249 7044 6253 7100
rect 6189 7040 6253 7044
rect 10946 7100 11010 7104
rect 10946 7044 10950 7100
rect 10950 7044 11006 7100
rect 11006 7044 11010 7100
rect 10946 7040 11010 7044
rect 11026 7100 11090 7104
rect 11026 7044 11030 7100
rect 11030 7044 11086 7100
rect 11086 7044 11090 7100
rect 11026 7040 11090 7044
rect 11106 7100 11170 7104
rect 11106 7044 11110 7100
rect 11110 7044 11166 7100
rect 11166 7044 11170 7100
rect 11106 7040 11170 7044
rect 11186 7100 11250 7104
rect 11186 7044 11190 7100
rect 11190 7044 11246 7100
rect 11246 7044 11250 7100
rect 11186 7040 11250 7044
rect 3450 6556 3514 6560
rect 3450 6500 3454 6556
rect 3454 6500 3510 6556
rect 3510 6500 3514 6556
rect 3450 6496 3514 6500
rect 3530 6556 3594 6560
rect 3530 6500 3534 6556
rect 3534 6500 3590 6556
rect 3590 6500 3594 6556
rect 3530 6496 3594 6500
rect 3610 6556 3674 6560
rect 3610 6500 3614 6556
rect 3614 6500 3670 6556
rect 3670 6500 3674 6556
rect 3610 6496 3674 6500
rect 3690 6556 3754 6560
rect 3690 6500 3694 6556
rect 3694 6500 3750 6556
rect 3750 6500 3754 6556
rect 3690 6496 3754 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 13445 6556 13509 6560
rect 13445 6500 13449 6556
rect 13449 6500 13505 6556
rect 13505 6500 13509 6556
rect 13445 6496 13509 6500
rect 13525 6556 13589 6560
rect 13525 6500 13529 6556
rect 13529 6500 13585 6556
rect 13585 6500 13589 6556
rect 13525 6496 13589 6500
rect 13605 6556 13669 6560
rect 13605 6500 13609 6556
rect 13609 6500 13665 6556
rect 13665 6500 13669 6556
rect 13605 6496 13669 6500
rect 13685 6556 13749 6560
rect 13685 6500 13689 6556
rect 13689 6500 13745 6556
rect 13745 6500 13749 6556
rect 13685 6496 13749 6500
rect 5949 6012 6013 6016
rect 5949 5956 5953 6012
rect 5953 5956 6009 6012
rect 6009 5956 6013 6012
rect 5949 5952 6013 5956
rect 6029 6012 6093 6016
rect 6029 5956 6033 6012
rect 6033 5956 6089 6012
rect 6089 5956 6093 6012
rect 6029 5952 6093 5956
rect 6109 6012 6173 6016
rect 6109 5956 6113 6012
rect 6113 5956 6169 6012
rect 6169 5956 6173 6012
rect 6109 5952 6173 5956
rect 6189 6012 6253 6016
rect 6189 5956 6193 6012
rect 6193 5956 6249 6012
rect 6249 5956 6253 6012
rect 6189 5952 6253 5956
rect 10946 6012 11010 6016
rect 10946 5956 10950 6012
rect 10950 5956 11006 6012
rect 11006 5956 11010 6012
rect 10946 5952 11010 5956
rect 11026 6012 11090 6016
rect 11026 5956 11030 6012
rect 11030 5956 11086 6012
rect 11086 5956 11090 6012
rect 11026 5952 11090 5956
rect 11106 6012 11170 6016
rect 11106 5956 11110 6012
rect 11110 5956 11166 6012
rect 11166 5956 11170 6012
rect 11106 5952 11170 5956
rect 11186 6012 11250 6016
rect 11186 5956 11190 6012
rect 11190 5956 11246 6012
rect 11246 5956 11250 6012
rect 11186 5952 11250 5956
rect 3450 5468 3514 5472
rect 3450 5412 3454 5468
rect 3454 5412 3510 5468
rect 3510 5412 3514 5468
rect 3450 5408 3514 5412
rect 3530 5468 3594 5472
rect 3530 5412 3534 5468
rect 3534 5412 3590 5468
rect 3590 5412 3594 5468
rect 3530 5408 3594 5412
rect 3610 5468 3674 5472
rect 3610 5412 3614 5468
rect 3614 5412 3670 5468
rect 3670 5412 3674 5468
rect 3610 5408 3674 5412
rect 3690 5468 3754 5472
rect 3690 5412 3694 5468
rect 3694 5412 3750 5468
rect 3750 5412 3754 5468
rect 3690 5408 3754 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 13445 5468 13509 5472
rect 13445 5412 13449 5468
rect 13449 5412 13505 5468
rect 13505 5412 13509 5468
rect 13445 5408 13509 5412
rect 13525 5468 13589 5472
rect 13525 5412 13529 5468
rect 13529 5412 13585 5468
rect 13585 5412 13589 5468
rect 13525 5408 13589 5412
rect 13605 5468 13669 5472
rect 13605 5412 13609 5468
rect 13609 5412 13665 5468
rect 13665 5412 13669 5468
rect 13605 5408 13669 5412
rect 13685 5468 13749 5472
rect 13685 5412 13689 5468
rect 13689 5412 13745 5468
rect 13745 5412 13749 5468
rect 13685 5408 13749 5412
rect 9444 5204 9508 5268
rect 5949 4924 6013 4928
rect 5949 4868 5953 4924
rect 5953 4868 6009 4924
rect 6009 4868 6013 4924
rect 5949 4864 6013 4868
rect 6029 4924 6093 4928
rect 6029 4868 6033 4924
rect 6033 4868 6089 4924
rect 6089 4868 6093 4924
rect 6029 4864 6093 4868
rect 6109 4924 6173 4928
rect 6109 4868 6113 4924
rect 6113 4868 6169 4924
rect 6169 4868 6173 4924
rect 6109 4864 6173 4868
rect 6189 4924 6253 4928
rect 6189 4868 6193 4924
rect 6193 4868 6249 4924
rect 6249 4868 6253 4924
rect 6189 4864 6253 4868
rect 10946 4924 11010 4928
rect 10946 4868 10950 4924
rect 10950 4868 11006 4924
rect 11006 4868 11010 4924
rect 10946 4864 11010 4868
rect 11026 4924 11090 4928
rect 11026 4868 11030 4924
rect 11030 4868 11086 4924
rect 11086 4868 11090 4924
rect 11026 4864 11090 4868
rect 11106 4924 11170 4928
rect 11106 4868 11110 4924
rect 11110 4868 11166 4924
rect 11166 4868 11170 4924
rect 11106 4864 11170 4868
rect 11186 4924 11250 4928
rect 11186 4868 11190 4924
rect 11190 4868 11246 4924
rect 11246 4868 11250 4924
rect 11186 4864 11250 4868
rect 3450 4380 3514 4384
rect 3450 4324 3454 4380
rect 3454 4324 3510 4380
rect 3510 4324 3514 4380
rect 3450 4320 3514 4324
rect 3530 4380 3594 4384
rect 3530 4324 3534 4380
rect 3534 4324 3590 4380
rect 3590 4324 3594 4380
rect 3530 4320 3594 4324
rect 3610 4380 3674 4384
rect 3610 4324 3614 4380
rect 3614 4324 3670 4380
rect 3670 4324 3674 4380
rect 3610 4320 3674 4324
rect 3690 4380 3754 4384
rect 3690 4324 3694 4380
rect 3694 4324 3750 4380
rect 3750 4324 3754 4380
rect 3690 4320 3754 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 13445 4380 13509 4384
rect 13445 4324 13449 4380
rect 13449 4324 13505 4380
rect 13505 4324 13509 4380
rect 13445 4320 13509 4324
rect 13525 4380 13589 4384
rect 13525 4324 13529 4380
rect 13529 4324 13585 4380
rect 13585 4324 13589 4380
rect 13525 4320 13589 4324
rect 13605 4380 13669 4384
rect 13605 4324 13609 4380
rect 13609 4324 13665 4380
rect 13665 4324 13669 4380
rect 13605 4320 13669 4324
rect 13685 4380 13749 4384
rect 13685 4324 13689 4380
rect 13689 4324 13745 4380
rect 13745 4324 13749 4380
rect 13685 4320 13749 4324
rect 9260 4252 9324 4316
rect 9076 4176 9140 4180
rect 9076 4120 9126 4176
rect 9126 4120 9140 4176
rect 9076 4116 9140 4120
rect 10732 3844 10796 3908
rect 5949 3836 6013 3840
rect 5949 3780 5953 3836
rect 5953 3780 6009 3836
rect 6009 3780 6013 3836
rect 5949 3776 6013 3780
rect 6029 3836 6093 3840
rect 6029 3780 6033 3836
rect 6033 3780 6089 3836
rect 6089 3780 6093 3836
rect 6029 3776 6093 3780
rect 6109 3836 6173 3840
rect 6109 3780 6113 3836
rect 6113 3780 6169 3836
rect 6169 3780 6173 3836
rect 6109 3776 6173 3780
rect 6189 3836 6253 3840
rect 6189 3780 6193 3836
rect 6193 3780 6249 3836
rect 6249 3780 6253 3836
rect 6189 3776 6253 3780
rect 10946 3836 11010 3840
rect 10946 3780 10950 3836
rect 10950 3780 11006 3836
rect 11006 3780 11010 3836
rect 10946 3776 11010 3780
rect 11026 3836 11090 3840
rect 11026 3780 11030 3836
rect 11030 3780 11086 3836
rect 11086 3780 11090 3836
rect 11026 3776 11090 3780
rect 11106 3836 11170 3840
rect 11106 3780 11110 3836
rect 11110 3780 11166 3836
rect 11166 3780 11170 3836
rect 11106 3776 11170 3780
rect 11186 3836 11250 3840
rect 11186 3780 11190 3836
rect 11190 3780 11246 3836
rect 11246 3780 11250 3836
rect 11186 3776 11250 3780
rect 3450 3292 3514 3296
rect 3450 3236 3454 3292
rect 3454 3236 3510 3292
rect 3510 3236 3514 3292
rect 3450 3232 3514 3236
rect 3530 3292 3594 3296
rect 3530 3236 3534 3292
rect 3534 3236 3590 3292
rect 3590 3236 3594 3292
rect 3530 3232 3594 3236
rect 3610 3292 3674 3296
rect 3610 3236 3614 3292
rect 3614 3236 3670 3292
rect 3670 3236 3674 3292
rect 3610 3232 3674 3236
rect 3690 3292 3754 3296
rect 3690 3236 3694 3292
rect 3694 3236 3750 3292
rect 3750 3236 3754 3292
rect 3690 3232 3754 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 13445 3292 13509 3296
rect 13445 3236 13449 3292
rect 13449 3236 13505 3292
rect 13505 3236 13509 3292
rect 13445 3232 13509 3236
rect 13525 3292 13589 3296
rect 13525 3236 13529 3292
rect 13529 3236 13585 3292
rect 13585 3236 13589 3292
rect 13525 3232 13589 3236
rect 13605 3292 13669 3296
rect 13605 3236 13609 3292
rect 13609 3236 13665 3292
rect 13665 3236 13669 3292
rect 13605 3232 13669 3236
rect 13685 3292 13749 3296
rect 13685 3236 13689 3292
rect 13689 3236 13745 3292
rect 13745 3236 13749 3292
rect 13685 3232 13749 3236
rect 5949 2748 6013 2752
rect 5949 2692 5953 2748
rect 5953 2692 6009 2748
rect 6009 2692 6013 2748
rect 5949 2688 6013 2692
rect 6029 2748 6093 2752
rect 6029 2692 6033 2748
rect 6033 2692 6089 2748
rect 6089 2692 6093 2748
rect 6029 2688 6093 2692
rect 6109 2748 6173 2752
rect 6109 2692 6113 2748
rect 6113 2692 6169 2748
rect 6169 2692 6173 2748
rect 6109 2688 6173 2692
rect 6189 2748 6253 2752
rect 6189 2692 6193 2748
rect 6193 2692 6249 2748
rect 6249 2692 6253 2748
rect 6189 2688 6253 2692
rect 10946 2748 11010 2752
rect 10946 2692 10950 2748
rect 10950 2692 11006 2748
rect 11006 2692 11010 2748
rect 10946 2688 11010 2692
rect 11026 2748 11090 2752
rect 11026 2692 11030 2748
rect 11030 2692 11086 2748
rect 11086 2692 11090 2748
rect 11026 2688 11090 2692
rect 11106 2748 11170 2752
rect 11106 2692 11110 2748
rect 11110 2692 11166 2748
rect 11166 2692 11170 2748
rect 11106 2688 11170 2692
rect 11186 2748 11250 2752
rect 11186 2692 11190 2748
rect 11190 2692 11246 2748
rect 11246 2692 11250 2748
rect 11186 2688 11250 2692
rect 3450 2204 3514 2208
rect 3450 2148 3454 2204
rect 3454 2148 3510 2204
rect 3510 2148 3514 2204
rect 3450 2144 3514 2148
rect 3530 2204 3594 2208
rect 3530 2148 3534 2204
rect 3534 2148 3590 2204
rect 3590 2148 3594 2204
rect 3530 2144 3594 2148
rect 3610 2204 3674 2208
rect 3610 2148 3614 2204
rect 3614 2148 3670 2204
rect 3670 2148 3674 2204
rect 3610 2144 3674 2148
rect 3690 2204 3754 2208
rect 3690 2148 3694 2204
rect 3694 2148 3750 2204
rect 3750 2148 3754 2204
rect 3690 2144 3754 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 13445 2204 13509 2208
rect 13445 2148 13449 2204
rect 13449 2148 13505 2204
rect 13505 2148 13509 2204
rect 13445 2144 13509 2148
rect 13525 2204 13589 2208
rect 13525 2148 13529 2204
rect 13529 2148 13585 2204
rect 13585 2148 13589 2204
rect 13525 2144 13589 2148
rect 13605 2204 13669 2208
rect 13605 2148 13609 2204
rect 13609 2148 13665 2204
rect 13665 2148 13669 2204
rect 13605 2144 13669 2148
rect 13685 2204 13749 2208
rect 13685 2148 13689 2204
rect 13689 2148 13745 2204
rect 13745 2148 13749 2204
rect 13685 2144 13749 2148
<< metal4 >>
rect 3442 17440 3763 17456
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3763 17440
rect 3442 16352 3763 17376
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3763 16352
rect 3442 15264 3763 16288
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3763 15264
rect 3442 14176 3763 15200
rect 5941 16896 6261 17456
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 15808 6261 16832
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 14720 6261 15744
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5579 14244 5645 14245
rect 5579 14180 5580 14244
rect 5644 14180 5645 14244
rect 5579 14179 5645 14180
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3763 14176
rect 3442 13088 3763 14112
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3763 13088
rect 3442 12000 3763 13024
rect 5211 12748 5277 12749
rect 5211 12684 5212 12748
rect 5276 12684 5277 12748
rect 5211 12683 5277 12684
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3763 12000
rect 3442 10912 3763 11936
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3763 10912
rect 3442 9824 3763 10848
rect 5214 10165 5274 12683
rect 5582 10165 5642 14179
rect 5941 13632 6261 14656
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 12544 6261 13568
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 11456 6261 12480
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 10368 6261 11392
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5211 10164 5277 10165
rect 5211 10100 5212 10164
rect 5276 10100 5277 10164
rect 5211 10099 5277 10100
rect 5579 10164 5645 10165
rect 5579 10100 5580 10164
rect 5644 10100 5645 10164
rect 5579 10099 5645 10100
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3763 9824
rect 3442 8736 3763 9760
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3763 8736
rect 3442 7648 3763 8672
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3763 7648
rect 3442 6560 3763 7584
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3763 6560
rect 3442 5472 3763 6496
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3763 5472
rect 3442 4384 3763 5408
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3763 4384
rect 3442 3296 3763 4320
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3763 3296
rect 3442 2208 3763 3232
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3763 2208
rect 3442 2128 3763 2144
rect 5941 9280 6261 10304
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 8192 6261 9216
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 7104 6261 8128
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 6016 6261 7040
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 4928 6261 5952
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 3840 6261 4864
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 2752 6261 3776
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2128 6261 2688
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 10938 16896 11259 17456
rect 13437 17440 13757 17456
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 11651 17236 11717 17237
rect 11651 17172 11652 17236
rect 11716 17172 11717 17236
rect 11651 17171 11717 17172
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11259 16896
rect 10938 15808 11259 16832
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11259 15808
rect 8891 14924 8957 14925
rect 8891 14860 8892 14924
rect 8956 14860 8957 14924
rect 8891 14859 8957 14860
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8894 13021 8954 14859
rect 10938 14720 11259 15744
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11259 14720
rect 10938 13632 11259 14656
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11259 13632
rect 8891 13020 8957 13021
rect 8891 12956 8892 13020
rect 8956 12956 8957 13020
rect 8891 12955 8957 12956
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8894 8533 8954 12955
rect 10938 12544 11259 13568
rect 11467 13428 11533 13429
rect 11467 13364 11468 13428
rect 11532 13364 11533 13428
rect 11467 13363 11533 13364
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11259 12544
rect 10938 11456 11259 12480
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11259 11456
rect 10938 10368 11259 11392
rect 11470 11253 11530 13363
rect 11654 11389 11714 17171
rect 13437 16352 13757 17376
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 15264 13757 16288
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 14176 13757 15200
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 13088 13757 14112
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 12000 13757 13024
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 11651 11388 11717 11389
rect 11651 11324 11652 11388
rect 11716 11324 11717 11388
rect 11651 11323 11717 11324
rect 11467 11252 11533 11253
rect 11467 11188 11468 11252
rect 11532 11188 11533 11252
rect 11467 11187 11533 11188
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11259 10368
rect 10731 9620 10797 9621
rect 10731 9556 10732 9620
rect 10796 9556 10797 9620
rect 10731 9555 10797 9556
rect 9259 9076 9325 9077
rect 9259 9012 9260 9076
rect 9324 9012 9325 9076
rect 9259 9011 9325 9012
rect 9075 8804 9141 8805
rect 9075 8740 9076 8804
rect 9140 8740 9141 8804
rect 9075 8739 9141 8740
rect 8891 8532 8957 8533
rect 8891 8468 8892 8532
rect 8956 8468 8957 8532
rect 8891 8467 8957 8468
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 9078 4181 9138 8739
rect 9262 4317 9322 9011
rect 9443 8260 9509 8261
rect 9443 8196 9444 8260
rect 9508 8196 9509 8260
rect 9443 8195 9509 8196
rect 9446 5269 9506 8195
rect 9443 5268 9509 5269
rect 9443 5204 9444 5268
rect 9508 5204 9509 5268
rect 9443 5203 9509 5204
rect 9259 4316 9325 4317
rect 9259 4252 9260 4316
rect 9324 4252 9325 4316
rect 9259 4251 9325 4252
rect 9075 4180 9141 4181
rect 9075 4116 9076 4180
rect 9140 4116 9141 4180
rect 9075 4115 9141 4116
rect 10734 3909 10794 9555
rect 10938 9280 11259 10304
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11259 9280
rect 10938 8192 11259 9216
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11259 8192
rect 10938 7104 11259 8128
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11259 7104
rect 10938 6016 11259 7040
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11259 6016
rect 10938 4928 11259 5952
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11259 4928
rect 10731 3908 10797 3909
rect 10731 3844 10732 3908
rect 10796 3844 10797 3908
rect 10731 3843 10797 3844
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10938 3840 11259 4864
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11259 3840
rect 10938 2752 11259 3776
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11259 2752
rect 10938 2128 11259 2688
rect 13437 10912 13757 11936
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 9824 13757 10848
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 8736 13757 9760
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 7648 13757 8672
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 6560 13757 7584
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 5472 13757 6496
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 4384 13757 5408
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 3296 13757 4320
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 13437 2208 13757 3232
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2128 13757 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9
timestamp 1608910539
transform 1 0 1932 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1472 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _35_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608910539
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608910539
transform 1 0 2760 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608910539
transform 1 0 2392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2208 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1608910539
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1608910539
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608910539
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608910539
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4140 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4048 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5060 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5612 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608910539
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608910539
transform 1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _31_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1608910539
transform 1 0 8740 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 8464 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608910539
transform 1 0 7636 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608910539
transform 1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608910539
transform 1 0 8372 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98
timestamp 1608910539
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8832 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10212 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9936 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_112
timestamp 1608910539
transform 1 0 11408 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 11040 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11500 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1608910539
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 12236 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608910539
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_128
timestamp 1608910539
transform 1 0 12880 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1608910539
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1608910539
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12972 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_157 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1608910539
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1608910539
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1608910539
transform 1 0 14996 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_16
timestamp 1608910539
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_11
timestamp 1608910539
transform 1 0 2116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1608910539
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1608910539
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1608910539
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1608910539
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608910539
transform 1 0 1564 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4140 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5980 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608910539
transform 1 0 5612 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1608910539
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8004 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608910539
transform 1 0 7452 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1608910539
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10028 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10856 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11684 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12512 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_139
timestamp 1608910539
transform 1 0 13892 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608910539
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp 1608910539
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1472 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_38
timestamp 1608910539
transform 1 0 4600 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1608910539
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608910539
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1608910539
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 6440 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1608910539
transform 1 0 6900 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1608910539
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1608910539
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1608910539
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7636 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608910539
transform 1 0 8464 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_90
timestamp 1608910539
transform 1 0 9384 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9476 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10304 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608910539
transform 1 0 8832 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1608910539
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_158
timestamp 1608910539
transform 1 0 15640 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14812 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_16
timestamp 1608910539
transform 1 0 2576 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2668 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1608910539
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1608910539
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 3680 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 3496 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4508 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_49
timestamp 1608910539
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 1608910539
transform 1 0 4968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1608910539
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1608910539
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1608910539
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6992 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7820 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8648 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_95
timestamp 1608910539
transform 1 0 9844 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1608910539
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10120 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp 1608910539
transform 1 0 11776 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11868 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1608910539
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 14352 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 13524 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_157
timestamp 1608910539
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 16008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2576 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4232 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1608910539
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp 1608910539
transform 1 0 5060 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5152 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6900 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8372 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608910539
transform 1 0 7728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1608910539
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608910539
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10764 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13892 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_155
timestamp 1608910539
transform 1 0 15364 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1608910539
transform 1 0 2852 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 2024 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2852 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1608910539
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 3680 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3220 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1608910539
transform 1 0 5060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_52
timestamp 1608910539
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_48
timestamp 1608910539
transform 1 0 5520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608910539
transform 1 0 5612 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1608910539
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 5980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5980 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6808 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1608910539
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7360 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8280 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8280 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608910539
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1608910539
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_97
timestamp 1608910539
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1608910539
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 10120 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10396 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_118
timestamp 1608910539
transform 1 0 11960 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_112
timestamp 1608910539
transform 1 0 11408 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1608910539
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1608910539
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608910539
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1608910539
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_141
timestamp 1608910539
transform 1 0 14076 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1608910539
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1608910539
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1608910539
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14628 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2208 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1608910539
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_21
timestamp 1608910539
transform 1 0 3036 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_62
timestamp 1608910539
transform 1 0 6808 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5980 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_79
timestamp 1608910539
transform 1 0 8372 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6900 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_87
timestamp 1608910539
transform 1 0 9108 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1608910539
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11408 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_139
timestamp 1608910539
transform 1 0 13892 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1608910539
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1608910539
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1932 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_41
timestamp 1608910539
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3404 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1608910539
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1608910539
transform 1 0 5244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5612 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 7452 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9752 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8924 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1608910539
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1608910539
transform 1 0 11408 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_136
timestamp 1608910539
transform 1 0 13616 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_156
timestamp 1608910539
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_148
timestamp 1608910539
transform 1 0 14720 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_10
timestamp 1608910539
transform 1 0 2024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2300 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1608910539
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 4508 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4784 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5612 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1608910539
transform 1 0 7636 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10028 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_117
timestamp 1608910539
transform 1 0 11868 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12512 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1608910539
transform 1 0 10856 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1608910539
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_133
timestamp 1608910539
transform 1 0 13340 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1608910539
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_16
timestamp 1608910539
transform 1 0 2576 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_22
timestamp 1608910539
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3220 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4876 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_78
timestamp 1608910539
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1608910539
transform 1 0 9660 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9752 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608910539
transform 1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_112
timestamp 1608910539
transform 1 0 11408 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11500 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_145
timestamp 1608910539
transform 1 0 14444 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_127
timestamp 1608910539
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12972 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1608910539
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608910539
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608910539
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4416 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5888 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10672 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1608910539
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1608910539
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608910539
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_10
timestamp 1608910539
transform 1 0 2024 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1608910539
transform 1 0 2852 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1608910539
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2576 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2944 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_38
timestamp 1608910539
transform 1 0 4600 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1608910539
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_36
timestamp 1608910539
transform 1 0 4416 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_42
timestamp 1608910539
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_49
timestamp 1608910539
transform 1 0 5612 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_45
timestamp 1608910539
transform 1 0 5244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608910539
transform 1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1608910539
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_56
timestamp 1608910539
transform 1 0 6256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5888 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 1608910539
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7636 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8096 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1608910539
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1608910539
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9752 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8924 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10028 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9936 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1608910539
transform 1 0 11316 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_105
timestamp 1608910539
transform 1 0 10764 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_110
timestamp 1608910539
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11408 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1608910539
transform 1 0 13432 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_128
timestamp 1608910539
transform 1 0 12880 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_141
timestamp 1608910539
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1608910539
transform 1 0 13248 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13524 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1608910539
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_158
timestamp 1608910539
transform 1 0 15640 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_146
timestamp 1608910539
transform 1 0 14536 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_10
timestamp 1608910539
transform 1 0 2024 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3404 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4232 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1608910539
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6992 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7820 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_94
timestamp 1608910539
transform 1 0 9752 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_91
timestamp 1608910539
transform 1 0 9476 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10028 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_145
timestamp 1608910539
transform 1 0 14444 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12696 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1608910539
transform 1 0 14168 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1608910539
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_19
timestamp 1608910539
transform 1 0 2852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1608910539
transform 1 0 1932 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_52
timestamp 1608910539
transform 1 0 5888 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_48
timestamp 1608910539
transform 1 0 5520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5980 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608910539
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_71
timestamp 1608910539
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 8740 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1608910539
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10120 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_113
timestamp 1608910539
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 11684 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_143
timestamp 1608910539
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_131
timestamp 1608910539
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1608910539
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1608910539
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_19
timestamp 1608910539
transform 1 0 2852 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4140 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1608910539
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5796 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_81
timestamp 1608910539
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1608910539
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8648 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608910539
transform 1 0 7636 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_91
timestamp 1608910539
transform 1 0 9476 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10580 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9752 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608910539
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1608910539
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_136
timestamp 1608910539
transform 1 0 13616 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_156
timestamp 1608910539
transform 1 0 15456 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_148
timestamp 1608910539
transform 1 0 14720 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_10
timestamp 1608910539
transform 1 0 2024 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2116 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_39
timestamp 1608910539
transform 1 0 4692 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4784 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6256 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7728 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1608910539
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1608910539
transform 1 0 9844 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10672 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608910539
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_140
timestamp 1608910539
transform 1 0 13984 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_127
timestamp 1608910539
transform 1 0 12788 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 12880 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1608910539
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1608910539
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_18
timestamp 1608910539
transform 1 0 2760 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_10
timestamp 1608910539
transform 1 0 2024 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_10
timestamp 1608910539
transform 1 0 2024 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2852 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2392 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_36
timestamp 1608910539
transform 1 0 4416 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1608910539
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_39
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3220 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1608910539
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_45
timestamp 1608910539
transform 1 0 5244 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5152 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5336 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_59
timestamp 1608910539
transform 1 0 6532 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1608910539
transform 1 0 5980 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1608910539
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_62
timestamp 1608910539
transform 1 0 6808 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_80
timestamp 1608910539
transform 1 0 8464 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7636 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 7544 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_96
timestamp 1608910539
transform 1 0 9936 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608910539
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10212 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9384 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10028 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_113
timestamp 1608910539
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1608910539
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1608910539
transform 1 0 11040 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_137
timestamp 1608910539
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_136
timestamp 1608910539
transform 1 0 13616 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1608910539
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_148
timestamp 1608910539
transform 1 0 14720 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1608910539
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1608910539
transform 1 0 14996 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1608910539
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1608910539
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 16008 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_10
timestamp 1608910539
transform 1 0 2024 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2300 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4784 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1608910539
transform 1 0 3956 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1608910539
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5612 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_78
timestamp 1608910539
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8372 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_95
timestamp 1608910539
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_115
timestamp 1608910539
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_107
timestamp 1608910539
transform 1 0 10948 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12512 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13340 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_21_153
timestamp 1608910539
transform 1 0 15180 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_149
timestamp 1608910539
transform 1 0 14812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14904 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1656 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4140 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6440 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5612 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_78
timestamp 1608910539
transform 1 0 8280 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7452 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8372 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1608910539
transform 1 0 12604 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11132 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1608910539
transform 1 0 13892 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12696 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13984 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_22_156
timestamp 1608910539
transform 1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1608910539
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1608910539
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 2668 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608910539
transform 1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608910539
transform 1 0 1564 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4140 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608910539
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_52
timestamp 1608910539
transform 1 0 5888 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 5244 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608910539
transform 1 0 4968 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_69
timestamp 1608910539
transform 1 0 7452 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_64
timestamp 1608910539
transform 1 0 6992 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7544 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9200 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10212 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1608910539
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 11684 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_141
timestamp 1608910539
transform 1 0 14076 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13248 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1608910539
transform 1 0 14168 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_158
timestamp 1608910539
transform 1 0 15640 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608910539
transform 1 0 14996 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_10
timestamp 1608910539
transform 1 0 2024 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1608910539
transform 1 0 6716 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_44
timestamp 1608910539
transform 1 0 5152 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5244 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_65
timestamp 1608910539
transform 1 0 7084 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7176 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1608910539
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608910539
transform 1 0 8832 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1608910539
transform 1 0 12512 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 12144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1608910539
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14352 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12880 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_156
timestamp 1608910539
transform 1 0 15456 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_20
timestamp 1608910539
transform 1 0 2944 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1608910539
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 1608910539
transform 1 0 2024 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1608910539
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1608910539
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_38
timestamp 1608910539
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1608910539
transform 1 0 4048 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_29
timestamp 1608910539
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1608910539
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1608910539
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1608910539
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1608910539
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608910539
transform 1 0 3220 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_51
timestamp 1608910539
transform 1 0 5796 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1608910539
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1608910539
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1608910539
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1608910539
transform 1 0 5244 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_78
timestamp 1608910539
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8740 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10212 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608910539
transform 1 0 11868 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_134
timestamp 1608910539
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1608910539
transform 1 0 13708 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1608910539
transform 1 0 14536 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608910539
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_11
timestamp 1608910539
transform 1 0 2116 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1608910539
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608910539
transform 1 0 2392 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608910539
transform 1 0 2024 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_19
timestamp 1608910539
transform 1 0 2852 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608910539
transform 1 0 2760 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_28
timestamp 1608910539
transform 1 0 3680 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1608910539
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1608910539
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1608910539
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1608910539
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608910539
transform 1 0 3496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608910539
transform 1 0 3128 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_36
timestamp 1608910539
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608910539
transform 1 0 4876 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608910539
transform 1 0 4508 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1608910539
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_44
timestamp 1608910539
transform 1 0 5152 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608910539
transform 1 0 5612 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_55
timestamp 1608910539
transform 1 0 6164 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_52
timestamp 1608910539
transform 1 0 5888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1608910539
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 6348 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 5980 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 6716 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_67
timestamp 1608910539
transform 1 0 7268 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1608910539
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1608910539
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1608910539
transform 1 0 6900 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1608910539
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 7084 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_80
timestamp 1608910539
transform 1 0 8464 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp 1608910539
transform 1 0 7820 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1608910539
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608910539
transform 1 0 7912 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7360 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_90
timestamp 1608910539
transform 1 0 9384 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1608910539
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608910539
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608910539
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_96
timestamp 1608910539
transform 1 0 9936 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1608910539
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1608910539
transform 1 0 10028 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_115
timestamp 1608910539
transform 1 0 11684 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_124
timestamp 1608910539
transform 1 0 12512 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1608910539
transform 1 0 10856 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12604 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11040 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_27_141
timestamp 1608910539
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12788 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13616 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_27_156
timestamp 1608910539
transform 1 0 15456 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1608910539
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1608910539
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14536 0 1 16864
box -38 -48 866 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 16400 1912 17200 2032 6 ccff_tail
port 2 nsew signal tristate
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_in[10]
port 4 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_in[11]
port 5 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_in[12]
port 6 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_in[13]
port 7 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 chany_bottom_in[14]
port 8 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_in[15]
port 9 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 chany_bottom_in[16]
port 10 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_in[17]
port 11 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_in[18]
port 12 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_in[19]
port 13 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[1]
port 14 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[2]
port 15 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[3]
port 16 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[4]
port 17 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[5]
port 18 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[6]
port 19 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 chany_bottom_in[7]
port 20 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[8]
port 21 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[9]
port 22 nsew signal input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 23 nsew signal tristate
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_out[10]
port 24 nsew signal tristate
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_out[11]
port 25 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_out[12]
port 26 nsew signal tristate
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_out[13]
port 27 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_out[14]
port 28 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_out[15]
port 29 nsew signal tristate
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_out[16]
port 30 nsew signal tristate
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_out[17]
port 31 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_out[18]
port 32 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_out[19]
port 33 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 34 nsew signal tristate
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 35 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[3]
port 36 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 37 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 chany_bottom_out[5]
port 38 nsew signal tristate
rlabel metal2 s 2686 0 2742 800 6 chany_bottom_out[6]
port 39 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_out[7]
port 40 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[8]
port 41 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_out[9]
port 42 nsew signal tristate
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_in[0]
port 43 nsew signal input
rlabel metal2 s 12898 19200 12954 20000 6 chany_top_in[10]
port 44 nsew signal input
rlabel metal2 s 13266 19200 13322 20000 6 chany_top_in[11]
port 45 nsew signal input
rlabel metal2 s 13634 19200 13690 20000 6 chany_top_in[12]
port 46 nsew signal input
rlabel metal2 s 14094 19200 14150 20000 6 chany_top_in[13]
port 47 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[14]
port 48 nsew signal input
rlabel metal2 s 14922 19200 14978 20000 6 chany_top_in[15]
port 49 nsew signal input
rlabel metal2 s 15290 19200 15346 20000 6 chany_top_in[16]
port 50 nsew signal input
rlabel metal2 s 15750 19200 15806 20000 6 chany_top_in[17]
port 51 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[18]
port 52 nsew signal input
rlabel metal2 s 16578 19200 16634 20000 6 chany_top_in[19]
port 53 nsew signal input
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_in[1]
port 54 nsew signal input
rlabel metal2 s 9586 19200 9642 20000 6 chany_top_in[2]
port 55 nsew signal input
rlabel metal2 s 9954 19200 10010 20000 6 chany_top_in[3]
port 56 nsew signal input
rlabel metal2 s 10414 19200 10470 20000 6 chany_top_in[4]
port 57 nsew signal input
rlabel metal2 s 10782 19200 10838 20000 6 chany_top_in[5]
port 58 nsew signal input
rlabel metal2 s 11242 19200 11298 20000 6 chany_top_in[6]
port 59 nsew signal input
rlabel metal2 s 11610 19200 11666 20000 6 chany_top_in[7]
port 60 nsew signal input
rlabel metal2 s 12070 19200 12126 20000 6 chany_top_in[8]
port 61 nsew signal input
rlabel metal2 s 12438 19200 12494 20000 6 chany_top_in[9]
port 62 nsew signal input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 63 nsew signal tristate
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_out[10]
port 64 nsew signal tristate
rlabel metal2 s 5078 19200 5134 20000 6 chany_top_out[11]
port 65 nsew signal tristate
rlabel metal2 s 5446 19200 5502 20000 6 chany_top_out[12]
port 66 nsew signal tristate
rlabel metal2 s 5906 19200 5962 20000 6 chany_top_out[13]
port 67 nsew signal tristate
rlabel metal2 s 6274 19200 6330 20000 6 chany_top_out[14]
port 68 nsew signal tristate
rlabel metal2 s 6734 19200 6790 20000 6 chany_top_out[15]
port 69 nsew signal tristate
rlabel metal2 s 7102 19200 7158 20000 6 chany_top_out[16]
port 70 nsew signal tristate
rlabel metal2 s 7562 19200 7618 20000 6 chany_top_out[17]
port 71 nsew signal tristate
rlabel metal2 s 7930 19200 7986 20000 6 chany_top_out[18]
port 72 nsew signal tristate
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[19]
port 73 nsew signal tristate
rlabel metal2 s 938 19200 994 20000 6 chany_top_out[1]
port 74 nsew signal tristate
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 75 nsew signal tristate
rlabel metal2 s 1766 19200 1822 20000 6 chany_top_out[3]
port 76 nsew signal tristate
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 77 nsew signal tristate
rlabel metal2 s 2594 19200 2650 20000 6 chany_top_out[5]
port 78 nsew signal tristate
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 79 nsew signal tristate
rlabel metal2 s 3422 19200 3478 20000 6 chany_top_out[7]
port 80 nsew signal tristate
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_out[8]
port 81 nsew signal tristate
rlabel metal2 s 4250 19200 4306 20000 6 chany_top_out[9]
port 82 nsew signal tristate
rlabel metal3 s 16400 9800 17200 9920 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew signal tristate
rlabel metal3 s 16400 13880 17200 14000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew signal input
rlabel metal3 s 16400 17824 17200 17944 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew signal tristate
rlabel metal3 s 0 3272 800 3392 6 left_grid_pin_16_
port 86 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 left_grid_pin_17_
port 87 nsew signal tristate
rlabel metal3 s 0 5176 800 5296 6 left_grid_pin_18_
port 88 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 left_grid_pin_19_
port 89 nsew signal tristate
rlabel metal3 s 0 7080 800 7200 6 left_grid_pin_20_
port 90 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 left_grid_pin_21_
port 91 nsew signal tristate
rlabel metal3 s 0 8984 800 9104 6 left_grid_pin_22_
port 92 nsew signal tristate
rlabel metal3 s 0 9936 800 10056 6 left_grid_pin_23_
port 93 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 left_grid_pin_24_
port 94 nsew signal tristate
rlabel metal3 s 0 11840 800 11960 6 left_grid_pin_25_
port 95 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 left_grid_pin_26_
port 96 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 left_grid_pin_27_
port 97 nsew signal tristate
rlabel metal3 s 0 14696 800 14816 6 left_grid_pin_28_
port 98 nsew signal tristate
rlabel metal3 s 0 15648 800 15768 6 left_grid_pin_29_
port 99 nsew signal tristate
rlabel metal3 s 0 16600 800 16720 6 left_grid_pin_30_
port 100 nsew signal tristate
rlabel metal3 s 0 17552 800 17672 6 left_grid_pin_31_
port 101 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 left_width_0_height_0__pin_0_
port 102 nsew signal input
rlabel metal3 s 0 416 800 536 6 left_width_0_height_0__pin_1_lower
port 103 nsew signal tristate
rlabel metal3 s 0 19456 800 19576 6 left_width_0_height_0__pin_1_upper
port 104 nsew signal tristate
rlabel metal2 s 16946 19200 17002 20000 6 prog_clk_0_N_out
port 105 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 prog_clk_0_S_out
port 106 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 prog_clk_0_W_in
port 107 nsew signal input
rlabel metal3 s 16400 5856 17200 5976 6 right_grid_pin_0_
port 108 nsew signal tristate
rlabel metal4 s 13437 2128 13757 17456 6 VPWR
port 109 nsew power bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VPWR
port 110 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 17456 6 VPWR
port 111 nsew power bidirectional
rlabel metal4 s 10939 2128 11259 17456 6 VGND
port 112 nsew ground bidirectional
rlabel metal4 s 5941 2128 6261 17456 6 VGND
port 113 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
