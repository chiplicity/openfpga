magic
tech EFS8A
magscale 1 2
timestamp 1602873085
<< locali >>
rect 2789 12631 2823 12733
rect 6653 11679 6687 11781
rect 6135 11169 6170 11203
rect 7147 11169 7182 11203
rect 18371 11169 18498 11203
rect 19475 11169 19510 11203
rect 5675 10557 5802 10591
rect 18003 10557 18130 10591
rect 21097 10523 21131 10625
rect 19383 10081 19418 10115
rect 25455 10081 25490 10115
rect 33701 9503 33735 9537
rect 33701 9469 33862 9503
rect 15663 9129 15669 9163
rect 15663 9061 15697 9129
rect 22787 8993 22822 9027
rect 30423 8993 30458 9027
rect 34069 8347 34103 8585
rect 15571 8279 15605 8347
rect 15571 8245 15577 8279
rect 15663 8041 15669 8075
rect 18975 8041 18981 8075
rect 26887 8041 26893 8075
rect 15663 7973 15697 8041
rect 18975 7973 19009 8041
rect 26887 7973 26921 8041
rect 5089 7327 5123 7429
rect 2520 7225 2592 7259
rect 22655 6953 22661 6987
rect 34155 6953 34161 6987
rect 22655 6885 22689 6953
rect 24328 6885 24396 6919
rect 34155 6885 34189 6953
rect 24961 6103 24995 6409
rect 28917 6239 28951 6409
rect 25599 6103 25633 6171
rect 25599 6069 25605 6103
rect 8027 5865 8033 5899
rect 24403 5865 24409 5899
rect 34247 5865 34253 5899
rect 8027 5797 8061 5865
rect 5089 5559 5123 5797
rect 22201 5763 22235 5865
rect 24403 5797 24437 5865
rect 34247 5797 34281 5865
rect 11621 5083 11655 5253
rect 12081 5015 12115 5117
rect 23305 5083 23339 5321
rect 8211 4777 8217 4811
rect 8211 4709 8245 4777
rect 35483 4709 35528 4743
rect 1535 4029 1662 4063
rect 22747 3689 22753 3723
rect 14105 3587 14139 3689
rect 22747 3621 22781 3689
rect 17049 3451 17083 3553
rect 24501 2907 24535 3077
rect 35725 2907 35759 3077
rect 9315 2839 9349 2907
rect 9315 2805 9321 2839
rect 13829 2295 13863 2397
rect 31953 2295 31987 2397
<< viali >>
rect 1593 12937 1627 12971
rect 35633 12937 35667 12971
rect 1409 12733 1443 12767
rect 2580 12733 2614 12767
rect 2789 12733 2823 12767
rect 4972 12733 5006 12767
rect 13001 12733 13035 12767
rect 13461 12733 13495 12767
rect 35449 12733 35483 12767
rect 36001 12733 36035 12767
rect 2053 12665 2087 12699
rect 2651 12597 2685 12631
rect 2789 12597 2823 12631
rect 3065 12597 3099 12631
rect 5043 12597 5077 12631
rect 5457 12597 5491 12631
rect 13185 12597 13219 12631
rect 1593 12393 1627 12427
rect 1409 12257 1443 12291
rect 2513 12257 2547 12291
rect 4123 12257 4157 12291
rect 5984 12257 6018 12291
rect 10241 12257 10275 12291
rect 11320 12257 11354 12291
rect 13093 12257 13127 12291
rect 2697 12121 2731 12155
rect 2053 12053 2087 12087
rect 2329 12053 2363 12087
rect 4215 12053 4249 12087
rect 6055 12053 6089 12087
rect 10425 12053 10459 12087
rect 11391 12053 11425 12087
rect 13277 12053 13311 12087
rect 14289 12053 14323 12087
rect 2973 11849 3007 11883
rect 14105 11849 14139 11883
rect 3617 11781 3651 11815
rect 6653 11781 6687 11815
rect 10425 11781 10459 11815
rect 1685 11713 1719 11747
rect 2145 11645 2179 11679
rect 2329 11645 2363 11679
rect 3341 11645 3375 11679
rect 3433 11645 3467 11679
rect 4956 11645 4990 11679
rect 5365 11645 5399 11679
rect 6653 11645 6687 11679
rect 6888 11645 6922 11679
rect 10241 11645 10275 11679
rect 11069 11645 11103 11679
rect 11320 11645 11354 11679
rect 14289 11645 14323 11679
rect 14749 11645 14783 11679
rect 18496 11645 18530 11679
rect 19752 11645 19786 11679
rect 20177 11645 20211 11679
rect 5043 11577 5077 11611
rect 6975 11577 7009 11611
rect 12173 11577 12207 11611
rect 15025 11577 15059 11611
rect 19855 11577 19889 11611
rect 2145 11509 2179 11543
rect 4169 11509 4203 11543
rect 6009 11509 6043 11543
rect 7389 11509 7423 11543
rect 10701 11509 10735 11543
rect 11391 11509 11425 11543
rect 11805 11509 11839 11543
rect 12449 11509 12483 11543
rect 13185 11509 13219 11543
rect 18567 11509 18601 11543
rect 18981 11509 19015 11543
rect 17003 11305 17037 11339
rect 35633 11305 35667 11339
rect 1869 11169 1903 11203
rect 2329 11169 2363 11203
rect 4112 11169 4146 11203
rect 4629 11169 4663 11203
rect 5156 11169 5190 11203
rect 6101 11169 6135 11203
rect 7113 11169 7147 11203
rect 8192 11169 8226 11203
rect 9689 11169 9723 11203
rect 10768 11169 10802 11203
rect 11805 11169 11839 11203
rect 13553 11169 13587 11203
rect 13645 11169 13679 11203
rect 14105 11169 14139 11203
rect 16900 11169 16934 11203
rect 18337 11169 18371 11203
rect 19441 11169 19475 11203
rect 22084 11169 22118 11203
rect 26684 11169 26718 11203
rect 34412 11169 34446 11203
rect 35449 11169 35483 11203
rect 2421 11101 2455 11135
rect 12449 11101 12483 11135
rect 14381 11101 14415 11135
rect 15669 11101 15703 11135
rect 5227 11033 5261 11067
rect 8263 11033 8297 11067
rect 9873 11033 9907 11067
rect 1777 10965 1811 10999
rect 4215 10965 4249 10999
rect 6239 10965 6273 10999
rect 7251 10965 7285 10999
rect 10839 10965 10873 10999
rect 18567 10965 18601 10999
rect 19579 10965 19613 10999
rect 22155 10965 22189 10999
rect 26755 10965 26789 10999
rect 34483 10965 34517 10999
rect 1593 10761 1627 10795
rect 4537 10761 4571 10795
rect 5181 10761 5215 10795
rect 5871 10761 5905 10795
rect 15301 10761 15335 10795
rect 18521 10761 18555 10795
rect 22661 10761 22695 10795
rect 26249 10761 26283 10795
rect 35357 10761 35391 10795
rect 13737 10693 13771 10727
rect 35633 10693 35667 10727
rect 2697 10625 2731 10659
rect 7573 10625 7607 10659
rect 8585 10625 8619 10659
rect 11805 10625 11839 10659
rect 18889 10625 18923 10659
rect 21097 10625 21131 10659
rect 1409 10557 1443 10591
rect 2789 10557 2823 10591
rect 3341 10557 3375 10591
rect 4353 10557 4387 10591
rect 5641 10557 5675 10591
rect 6561 10557 6595 10591
rect 8033 10557 8067 10591
rect 10368 10557 10402 10591
rect 10793 10557 10827 10591
rect 11380 10557 11414 10591
rect 11483 10557 11517 10591
rect 12541 10557 12575 10591
rect 14197 10557 14231 10591
rect 14565 10557 14599 10591
rect 15853 10557 15887 10591
rect 16405 10557 16439 10591
rect 17969 10557 18003 10591
rect 19108 10557 19142 10591
rect 19901 10557 19935 10591
rect 20872 10557 20906 10591
rect 21868 10557 21902 10591
rect 22293 10557 22327 10591
rect 25764 10557 25798 10591
rect 26744 10557 26778 10591
rect 27169 10557 27203 10591
rect 27788 10557 27822 10591
rect 28181 10557 28215 10591
rect 33308 10557 33342 10591
rect 35449 10557 35483 10591
rect 36001 10557 36035 10591
rect 2053 10489 2087 10523
rect 10471 10489 10505 10523
rect 14841 10489 14875 10523
rect 15761 10489 15795 10523
rect 16589 10489 16623 10523
rect 19211 10489 19245 10523
rect 21097 10489 21131 10523
rect 21373 10489 21407 10523
rect 26847 10489 26881 10523
rect 2881 10421 2915 10455
rect 4077 10421 4111 10455
rect 6193 10421 6227 10455
rect 7021 10421 7055 10455
rect 8217 10421 8251 10455
rect 8861 10421 8895 10455
rect 9321 10421 9355 10455
rect 9873 10421 9907 10455
rect 11253 10421 11287 10455
rect 12173 10421 12207 10455
rect 12725 10421 12759 10455
rect 16865 10421 16899 10455
rect 18199 10421 18233 10455
rect 19533 10421 19567 10455
rect 20959 10421 20993 10455
rect 21971 10421 22005 10455
rect 25835 10421 25869 10455
rect 26617 10421 26651 10455
rect 27859 10421 27893 10455
rect 33379 10421 33413 10455
rect 33701 10421 33735 10455
rect 34437 10421 34471 10455
rect 3525 10217 3559 10251
rect 4169 10217 4203 10251
rect 6745 10217 6779 10251
rect 13461 10217 13495 10251
rect 14105 10217 14139 10251
rect 27169 10217 27203 10251
rect 35633 10217 35667 10251
rect 27445 10149 27479 10183
rect 1685 10081 1719 10115
rect 1869 10081 1903 10115
rect 3008 10081 3042 10115
rect 4353 10081 4387 10115
rect 4537 10081 4571 10115
rect 5708 10081 5742 10115
rect 6929 10081 6963 10115
rect 7113 10081 7147 10115
rect 8652 10081 8686 10115
rect 10517 10081 10551 10115
rect 10977 10081 11011 10115
rect 12817 10081 12851 10115
rect 16129 10081 16163 10115
rect 16451 10081 16485 10115
rect 17785 10081 17819 10115
rect 18245 10081 18279 10115
rect 19349 10081 19383 10115
rect 20948 10081 20982 10115
rect 21992 10081 22026 10115
rect 22937 10081 22971 10115
rect 24409 10081 24443 10115
rect 25421 10081 25455 10115
rect 28860 10081 28894 10115
rect 33492 10081 33526 10115
rect 34488 10081 34522 10115
rect 35449 10081 35483 10115
rect 36588 10081 36622 10115
rect 1961 10013 1995 10047
rect 2513 10013 2547 10047
rect 11069 10013 11103 10047
rect 13185 10013 13219 10047
rect 16313 10013 16347 10047
rect 18521 10013 18555 10047
rect 21465 10013 21499 10047
rect 27353 10013 27387 10047
rect 27997 10013 28031 10047
rect 34575 10013 34609 10047
rect 8723 9945 8757 9979
rect 12982 9945 13016 9979
rect 28963 9945 28997 9979
rect 33563 9945 33597 9979
rect 2789 9877 2823 9911
rect 3111 9877 3145 9911
rect 5779 9877 5813 9911
rect 11713 9877 11747 9911
rect 12541 9877 12575 9911
rect 13093 9877 13127 9911
rect 14565 9877 14599 9911
rect 19487 9877 19521 9911
rect 19901 9877 19935 9911
rect 21051 9877 21085 9911
rect 21741 9877 21775 9911
rect 22063 9877 22097 9911
rect 23121 9877 23155 9911
rect 24133 9877 24167 9911
rect 24593 9877 24627 9911
rect 25559 9877 25593 9911
rect 36691 9877 36725 9911
rect 4077 9673 4111 9707
rect 6561 9673 6595 9707
rect 8217 9673 8251 9707
rect 10241 9673 10275 9707
rect 11529 9673 11563 9707
rect 11805 9673 11839 9707
rect 15485 9673 15519 9707
rect 15853 9673 15887 9707
rect 17509 9673 17543 9707
rect 19349 9673 19383 9707
rect 20913 9673 20947 9707
rect 22385 9673 22419 9707
rect 32229 9673 32263 9707
rect 33517 9673 33551 9707
rect 35541 9673 35575 9707
rect 35909 9673 35943 9707
rect 36645 9673 36679 9707
rect 6285 9605 6319 9639
rect 13461 9605 13495 9639
rect 25513 9605 25547 9639
rect 29423 9605 29457 9639
rect 3065 9537 3099 9571
rect 7205 9537 7239 9571
rect 9965 9537 9999 9571
rect 12541 9537 12575 9571
rect 16037 9537 16071 9571
rect 16957 9537 16991 9571
rect 21741 9537 21775 9571
rect 23949 9537 23983 9571
rect 27445 9537 27479 9571
rect 33701 9537 33735 9571
rect 34345 9537 34379 9571
rect 1593 9469 1627 9503
rect 1961 9469 1995 9503
rect 2513 9469 2547 9503
rect 4445 9469 4479 9503
rect 5089 9469 5123 9503
rect 5273 9469 5307 9503
rect 8585 9469 8619 9503
rect 8861 9469 8895 9503
rect 10609 9469 10643 9503
rect 10977 9469 11011 9503
rect 13185 9469 13219 9503
rect 15025 9469 15059 9503
rect 18337 9469 18371 9503
rect 18613 9469 18647 9503
rect 19901 9469 19935 9503
rect 20177 9469 20211 9503
rect 24133 9469 24167 9503
rect 24593 9469 24627 9503
rect 26408 9469 26442 9503
rect 29352 9469 29386 9503
rect 29837 9469 29871 9503
rect 30297 9469 30331 9503
rect 30757 9469 30791 9503
rect 31820 9469 31854 9503
rect 32816 9469 32850 9503
rect 35357 9469 35391 9503
rect 36461 9469 36495 9503
rect 37013 9469 37047 9503
rect 2145 9401 2179 9435
rect 3157 9401 3191 9435
rect 3709 9401 3743 9435
rect 6929 9401 6963 9435
rect 7021 9401 7055 9435
rect 12633 9401 12667 9435
rect 13829 9401 13863 9435
rect 14289 9401 14323 9435
rect 16129 9401 16163 9435
rect 16681 9401 16715 9435
rect 21465 9401 21499 9435
rect 21557 9401 21591 9435
rect 24869 9401 24903 9435
rect 27261 9401 27295 9435
rect 27537 9401 27571 9435
rect 28089 9401 28123 9435
rect 31907 9401 31941 9435
rect 35173 9401 35207 9435
rect 2789 9333 2823 9367
rect 5733 9333 5767 9367
rect 7849 9333 7883 9367
rect 8493 9333 8527 9367
rect 9413 9333 9447 9367
rect 10517 9333 10551 9367
rect 12265 9333 12299 9367
rect 14657 9333 14691 9367
rect 17877 9333 17911 9367
rect 18153 9333 18187 9367
rect 19901 9333 19935 9367
rect 22937 9333 22971 9367
rect 26479 9333 26513 9367
rect 26893 9333 26927 9367
rect 28365 9333 28399 9367
rect 28825 9333 28859 9367
rect 30481 9333 30515 9367
rect 32597 9333 32631 9367
rect 32919 9333 32953 9367
rect 33931 9333 33965 9367
rect 34713 9333 34747 9367
rect 37473 9333 37507 9367
rect 1961 9129 1995 9163
rect 3433 9129 3467 9163
rect 11069 9129 11103 9163
rect 11529 9129 11563 9163
rect 15669 9129 15703 9163
rect 16221 9129 16255 9163
rect 16497 9129 16531 9163
rect 18153 9129 18187 9163
rect 18705 9129 18739 9163
rect 20085 9129 20119 9163
rect 23903 9129 23937 9163
rect 24409 9129 24443 9163
rect 28273 9129 28307 9163
rect 28641 9129 28675 9163
rect 2329 9061 2363 9095
rect 2605 9061 2639 9095
rect 3157 9061 3191 9095
rect 4261 9061 4295 9095
rect 7389 9061 7423 9095
rect 11805 9061 11839 9095
rect 13369 9061 13403 9095
rect 17233 9061 17267 9095
rect 18521 9061 18555 9095
rect 21281 9061 21315 9095
rect 21373 9061 21407 9095
rect 27353 9061 27387 9095
rect 27445 9061 27479 9095
rect 29009 9061 29043 9095
rect 34069 9061 34103 9095
rect 35633 9061 35667 9095
rect 1476 8993 1510 9027
rect 5641 8993 5675 9027
rect 5917 8993 5951 9027
rect 10057 8993 10091 9027
rect 10517 8993 10551 9027
rect 15301 8993 15335 9027
rect 18613 8993 18647 9027
rect 19165 8993 19199 9027
rect 22753 8993 22787 9027
rect 23832 8993 23866 9027
rect 24869 8993 24903 9027
rect 25421 8993 25455 9027
rect 30389 8993 30423 9027
rect 32321 8993 32355 9027
rect 32689 8993 32723 9027
rect 2513 8925 2547 8959
rect 4169 8925 4203 8959
rect 6101 8925 6135 8959
rect 7297 8925 7331 8959
rect 7573 8925 7607 8959
rect 10609 8925 10643 8959
rect 11713 8925 11747 8959
rect 11989 8925 12023 8959
rect 13277 8925 13311 8959
rect 13553 8925 13587 8959
rect 17141 8925 17175 8959
rect 17417 8925 17451 8959
rect 21925 8925 21959 8959
rect 25605 8925 25639 8959
rect 27997 8925 28031 8959
rect 28917 8925 28951 8959
rect 29193 8925 29227 8959
rect 32873 8925 32907 8959
rect 33977 8925 34011 8959
rect 34253 8925 34287 8959
rect 35541 8925 35575 8959
rect 4721 8857 4755 8891
rect 5733 8857 5767 8891
rect 8493 8857 8527 8891
rect 16865 8857 16899 8891
rect 19717 8857 19751 8891
rect 30527 8857 30561 8891
rect 36093 8857 36127 8891
rect 1547 8789 1581 8823
rect 3893 8789 3927 8823
rect 5273 8789 5307 8823
rect 6929 8789 6963 8823
rect 8861 8789 8895 8823
rect 12817 8789 12851 8823
rect 22293 8789 22327 8823
rect 22891 8789 22925 8823
rect 27169 8789 27203 8823
rect 31309 8789 31343 8823
rect 33241 8789 33275 8823
rect 33609 8789 33643 8823
rect 34989 8789 35023 8823
rect 2421 8585 2455 8619
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 8033 8585 8067 8619
rect 8677 8585 8711 8619
rect 10149 8585 10183 8619
rect 13461 8585 13495 8619
rect 17095 8585 17129 8619
rect 22385 8585 22419 8619
rect 22753 8585 22787 8619
rect 23949 8585 23983 8619
rect 25329 8585 25363 8619
rect 26801 8585 26835 8619
rect 28733 8585 28767 8619
rect 32781 8585 32815 8619
rect 34069 8585 34103 8619
rect 36001 8585 36035 8619
rect 36277 8585 36311 8619
rect 36645 8585 36679 8619
rect 3617 8517 3651 8551
rect 8309 8517 8343 8551
rect 10425 8517 10459 8551
rect 13829 8517 13863 8551
rect 18889 8517 18923 8551
rect 19257 8517 19291 8551
rect 1501 8449 1535 8483
rect 2145 8449 2179 8483
rect 5273 8449 5307 8483
rect 5641 8449 5675 8483
rect 10885 8449 10919 8483
rect 11529 8449 11563 8483
rect 12817 8449 12851 8483
rect 17877 8449 17911 8483
rect 18337 8449 18371 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 21465 8449 21499 8483
rect 27721 8449 27755 8483
rect 29653 8449 29687 8483
rect 33333 8449 33367 8483
rect 33977 8449 34011 8483
rect 7113 8381 7147 8415
rect 8861 8381 8895 8415
rect 9321 8381 9355 8415
rect 14048 8381 14082 8415
rect 15209 8381 15243 8415
rect 16773 8381 16807 8415
rect 16992 8381 17026 8415
rect 21189 8381 21223 8415
rect 24317 8381 24351 8415
rect 24777 8381 24811 8415
rect 25053 8381 25087 8415
rect 25881 8381 25915 8415
rect 31217 8381 31251 8415
rect 32137 8381 32171 8415
rect 35541 8517 35575 8551
rect 34989 8449 35023 8483
rect 37703 8449 37737 8483
rect 36461 8381 36495 8415
rect 37616 8381 37650 8415
rect 38025 8381 38059 8415
rect 1593 8313 1627 8347
rect 3065 8313 3099 8347
rect 3157 8313 3191 8347
rect 5365 8313 5399 8347
rect 7434 8313 7468 8347
rect 10977 8313 11011 8347
rect 12541 8313 12575 8347
rect 12633 8313 12667 8347
rect 14151 8313 14185 8347
rect 18429 8313 18463 8347
rect 19993 8313 20027 8347
rect 21557 8313 21591 8347
rect 22109 8313 22143 8347
rect 23489 8313 23523 8347
rect 26243 8313 26277 8347
rect 27813 8313 27847 8347
rect 28365 8313 28399 8347
rect 29377 8313 29411 8347
rect 29469 8313 29503 8347
rect 31125 8313 31159 8347
rect 31538 8313 31572 8347
rect 33425 8313 33459 8347
rect 34069 8313 34103 8347
rect 34713 8313 34747 8347
rect 35081 8313 35115 8347
rect 2881 8245 2915 8279
rect 4997 8245 5031 8279
rect 6193 8245 6227 8279
rect 6653 8245 6687 8279
rect 8953 8245 8987 8279
rect 11897 8245 11931 8279
rect 12265 8245 12299 8279
rect 14565 8245 14599 8279
rect 15117 8245 15151 8279
rect 15577 8245 15611 8279
rect 16129 8245 16163 8279
rect 16497 8245 16531 8279
rect 17417 8245 17451 8279
rect 19625 8245 19659 8279
rect 20821 8245 20855 8279
rect 25789 8245 25823 8279
rect 27261 8245 27295 8279
rect 29009 8245 29043 8279
rect 30389 8245 30423 8279
rect 32413 8245 32447 8279
rect 34253 8245 34287 8279
rect 37105 8245 37139 8279
rect 2053 8041 2087 8075
rect 3065 8041 3099 8075
rect 3433 8041 3467 8075
rect 3709 8041 3743 8075
rect 6653 8041 6687 8075
rect 7665 8041 7699 8075
rect 8033 8041 8067 8075
rect 8401 8041 8435 8075
rect 10517 8041 10551 8075
rect 10885 8041 10919 8075
rect 11897 8041 11931 8075
rect 15025 8041 15059 8075
rect 15669 8041 15703 8075
rect 16221 8041 16255 8075
rect 18981 8041 19015 8075
rect 19809 8041 19843 8075
rect 22109 8041 22143 8075
rect 23673 8041 23707 8075
rect 24317 8041 24351 8075
rect 25881 8041 25915 8075
rect 26893 8041 26927 8075
rect 27445 8041 27479 8075
rect 27813 8041 27847 8075
rect 33425 8041 33459 8075
rect 34345 8041 34379 8075
rect 35909 8041 35943 8075
rect 1685 7973 1719 8007
rect 2466 7973 2500 8007
rect 4261 7973 4295 8007
rect 4813 7973 4847 8007
rect 7107 7973 7141 8007
rect 11298 7973 11332 8007
rect 12909 7973 12943 8007
rect 13461 7973 13495 8007
rect 16497 7973 16531 8007
rect 17141 7973 17175 8007
rect 17233 7973 17267 8007
rect 17785 7973 17819 8007
rect 21281 7973 21315 8007
rect 21833 7973 21867 8007
rect 22845 7973 22879 8007
rect 28089 7973 28123 8007
rect 28641 7973 28675 8007
rect 32499 7973 32533 8007
rect 35081 7973 35115 8007
rect 2145 7905 2179 7939
rect 5641 7905 5675 7939
rect 6745 7905 6779 7939
rect 8493 7905 8527 7939
rect 10000 7905 10034 7939
rect 10977 7905 11011 7939
rect 12541 7905 12575 7939
rect 15301 7905 15335 7939
rect 18613 7905 18647 7939
rect 19533 7905 19567 7939
rect 24869 7905 24903 7939
rect 25421 7905 25455 7939
rect 30481 7905 30515 7939
rect 31033 7905 31067 7939
rect 33920 7905 33954 7939
rect 36461 7905 36495 7939
rect 4169 7837 4203 7871
rect 10103 7837 10137 7871
rect 12173 7837 12207 7871
rect 12817 7837 12851 7871
rect 20729 7837 20763 7871
rect 21189 7837 21223 7871
rect 22753 7837 22787 7871
rect 23397 7837 23431 7871
rect 24777 7837 24811 7871
rect 25605 7837 25639 7871
rect 26525 7837 26559 7871
rect 28549 7837 28583 7871
rect 29193 7837 29227 7871
rect 31217 7837 31251 7871
rect 32137 7837 32171 7871
rect 34989 7837 35023 7871
rect 35633 7837 35667 7871
rect 5825 7769 5859 7803
rect 16865 7769 16899 7803
rect 34023 7769 34057 7803
rect 36645 7769 36679 7803
rect 5273 7701 5307 7735
rect 6285 7701 6319 7735
rect 8677 7701 8711 7735
rect 18337 7701 18371 7735
rect 29469 7701 29503 7735
rect 33057 7701 33091 7735
rect 34805 7701 34839 7735
rect 3157 7497 3191 7531
rect 4905 7497 4939 7531
rect 7757 7497 7791 7531
rect 9965 7497 9999 7531
rect 11529 7497 11563 7531
rect 13461 7497 13495 7531
rect 15485 7497 15519 7531
rect 17417 7497 17451 7531
rect 18981 7497 19015 7531
rect 20913 7497 20947 7531
rect 21281 7497 21315 7531
rect 21557 7497 21591 7531
rect 24869 7497 24903 7531
rect 26985 7497 27019 7531
rect 27629 7497 27663 7531
rect 28641 7497 28675 7531
rect 32505 7497 32539 7531
rect 33057 7497 33091 7531
rect 34253 7497 34287 7531
rect 36277 7497 36311 7531
rect 3801 7429 3835 7463
rect 4169 7429 4203 7463
rect 5089 7429 5123 7463
rect 13829 7429 13863 7463
rect 22385 7429 22419 7463
rect 27951 7429 27985 7463
rect 30665 7429 30699 7463
rect 36001 7429 36035 7463
rect 5273 7361 5307 7395
rect 6285 7361 6319 7395
rect 6837 7361 6871 7395
rect 10609 7361 10643 7395
rect 14289 7361 14323 7395
rect 16037 7361 16071 7395
rect 16681 7361 16715 7395
rect 18061 7361 18095 7395
rect 19993 7361 20027 7395
rect 21833 7361 21867 7395
rect 23765 7361 23799 7395
rect 24133 7361 24167 7395
rect 26065 7361 26099 7395
rect 27261 7361 27295 7395
rect 29377 7361 29411 7395
rect 31401 7361 31435 7395
rect 33333 7361 33367 7395
rect 34989 7361 35023 7395
rect 36553 7361 36587 7395
rect 36829 7361 36863 7395
rect 2237 7293 2271 7327
rect 3433 7293 3467 7327
rect 3985 7293 4019 7327
rect 4537 7293 4571 7327
rect 5089 7293 5123 7327
rect 8125 7293 8159 7327
rect 8861 7293 8895 7327
rect 9045 7293 9079 7327
rect 12541 7293 12575 7327
rect 14657 7293 14691 7327
rect 14933 7293 14967 7327
rect 25329 7293 25363 7327
rect 27880 7293 27914 7327
rect 28273 7293 28307 7327
rect 30849 7293 30883 7327
rect 31309 7293 31343 7327
rect 2486 7225 2520 7259
rect 5365 7225 5399 7259
rect 5917 7225 5951 7259
rect 6653 7225 6687 7259
rect 7199 7225 7233 7259
rect 8493 7225 8527 7259
rect 10517 7225 10551 7259
rect 10971 7225 11005 7259
rect 15117 7225 15151 7259
rect 16129 7225 16163 7259
rect 17877 7225 17911 7259
rect 18423 7225 18457 7259
rect 20314 7225 20348 7259
rect 21925 7225 21959 7259
rect 22845 7225 22879 7259
rect 23857 7225 23891 7259
rect 26386 7225 26420 7259
rect 29469 7225 29503 7259
rect 30021 7225 30055 7259
rect 33425 7225 33459 7259
rect 33977 7225 34011 7259
rect 35081 7225 35115 7259
rect 35633 7225 35667 7259
rect 36645 7225 36679 7259
rect 1777 7157 1811 7191
rect 2145 7157 2179 7191
rect 8677 7157 8711 7191
rect 11805 7157 11839 7191
rect 12173 7157 12207 7191
rect 12909 7157 12943 7191
rect 15853 7157 15887 7191
rect 17141 7157 17175 7191
rect 19349 7157 19383 7191
rect 19809 7157 19843 7191
rect 23397 7157 23431 7191
rect 25881 7157 25915 7191
rect 29101 7157 29135 7191
rect 30297 7157 30331 7191
rect 32229 7157 32263 7191
rect 34713 7157 34747 7191
rect 1685 6953 1719 6987
rect 2145 6953 2179 6987
rect 3157 6953 3191 6987
rect 4353 6953 4387 6987
rect 5641 6953 5675 6987
rect 6009 6953 6043 6987
rect 7665 6953 7699 6987
rect 10609 6953 10643 6987
rect 11989 6953 12023 6987
rect 14473 6953 14507 6987
rect 15761 6953 15795 6987
rect 16313 6953 16347 6987
rect 18153 6953 18187 6987
rect 18613 6953 18647 6987
rect 19993 6953 20027 6987
rect 22661 6953 22695 6987
rect 23213 6953 23247 6987
rect 24961 6953 24995 6987
rect 26065 6953 26099 6987
rect 26939 6953 26973 6987
rect 27721 6953 27755 6987
rect 28733 6953 28767 6987
rect 29285 6953 29319 6987
rect 30481 6953 30515 6987
rect 31125 6953 31159 6987
rect 34161 6953 34195 6987
rect 36461 6953 36495 6987
rect 2558 6885 2592 6919
rect 3433 6885 3467 6919
rect 4813 6885 4847 6919
rect 6377 6885 6411 6919
rect 7849 6885 7883 6919
rect 7941 6885 7975 6919
rect 9827 6885 9861 6919
rect 11390 6885 11424 6919
rect 13001 6885 13035 6919
rect 13553 6885 13587 6919
rect 16859 6885 16893 6919
rect 18889 6885 18923 6919
rect 20361 6885 20395 6919
rect 21465 6885 21499 6919
rect 24294 6885 24328 6919
rect 28175 6885 28209 6919
rect 29923 6885 29957 6919
rect 35449 6885 35483 6919
rect 35903 6885 35937 6919
rect 36737 6885 36771 6919
rect 2237 6817 2271 6851
rect 5365 6817 5399 6851
rect 9724 6817 9758 6851
rect 11069 6817 11103 6851
rect 15301 6817 15335 6851
rect 16497 6817 16531 6851
rect 20913 6817 20947 6851
rect 21097 6817 21131 6851
rect 23489 6817 23523 6851
rect 26836 6817 26870 6851
rect 32137 6817 32171 6851
rect 32689 6817 32723 6851
rect 34713 6817 34747 6851
rect 4721 6749 4755 6783
rect 6285 6749 6319 6783
rect 6561 6749 6595 6783
rect 8125 6749 8159 6783
rect 12909 6749 12943 6783
rect 18797 6749 18831 6783
rect 19441 6749 19475 6783
rect 22293 6749 22327 6783
rect 24041 6749 24075 6783
rect 27813 6749 27847 6783
rect 29561 6749 29595 6783
rect 30849 6749 30883 6783
rect 31585 6749 31619 6783
rect 32873 6749 32907 6783
rect 33793 6749 33827 6783
rect 35541 6749 35575 6783
rect 9137 6681 9171 6715
rect 10241 6681 10275 6715
rect 15485 6681 15519 6715
rect 7297 6613 7331 6647
rect 8861 6613 8895 6647
rect 12541 6613 12575 6647
rect 17417 6613 17451 6647
rect 21925 6613 21959 6647
rect 23857 6613 23891 6647
rect 27353 6613 27387 6647
rect 33333 6613 33367 6647
rect 34989 6613 35023 6647
rect 3617 6409 3651 6443
rect 4353 6409 4387 6443
rect 6561 6409 6595 6443
rect 10793 6409 10827 6443
rect 13461 6409 13495 6443
rect 15761 6409 15795 6443
rect 17141 6409 17175 6443
rect 18521 6409 18555 6443
rect 19809 6409 19843 6443
rect 24777 6409 24811 6443
rect 24961 6409 24995 6443
rect 25053 6409 25087 6443
rect 28917 6409 28951 6443
rect 29009 6409 29043 6443
rect 32597 6409 32631 6443
rect 34345 6409 34379 6443
rect 36001 6409 36035 6443
rect 6193 6341 6227 6375
rect 11529 6341 11563 6375
rect 17509 6341 17543 6375
rect 2053 6273 2087 6307
rect 5273 6273 5307 6307
rect 5917 6273 5951 6307
rect 8217 6273 8251 6307
rect 12541 6273 12575 6307
rect 13185 6273 13219 6307
rect 16221 6273 16255 6307
rect 20361 6273 20395 6307
rect 22385 6273 22419 6307
rect 3868 6205 3902 6239
rect 6872 6205 6906 6239
rect 7297 6205 7331 6239
rect 9229 6205 9263 6239
rect 9965 6205 9999 6239
rect 10241 6205 10275 6239
rect 11345 6205 11379 6239
rect 13921 6205 13955 6239
rect 14105 6205 14139 6239
rect 21741 6205 21775 6239
rect 22109 6205 22143 6239
rect 22293 6205 22327 6239
rect 23673 6205 23707 6239
rect 24225 6205 24259 6239
rect 1961 6137 1995 6171
rect 2415 6137 2449 6171
rect 3341 6137 3375 6171
rect 5365 6137 5399 6171
rect 6975 6137 7009 6171
rect 7757 6137 7791 6171
rect 8309 6137 8343 6171
rect 8861 6137 8895 6171
rect 12633 6137 12667 6171
rect 14013 6137 14047 6171
rect 16129 6137 16163 6171
rect 16583 6137 16617 6171
rect 17877 6137 17911 6171
rect 18797 6137 18831 6171
rect 18889 6137 18923 6171
rect 19441 6137 19475 6171
rect 20453 6137 20487 6171
rect 21005 6137 21039 6171
rect 24409 6137 24443 6171
rect 25237 6273 25271 6307
rect 26801 6273 26835 6307
rect 27077 6273 27111 6307
rect 30941 6341 30975 6375
rect 32137 6341 32171 6375
rect 33885 6341 33919 6375
rect 33333 6273 33367 6307
rect 34989 6273 35023 6307
rect 36829 6273 36863 6307
rect 28917 6205 28951 6239
rect 29285 6205 29319 6239
rect 29745 6205 29779 6239
rect 31125 6205 31159 6239
rect 31585 6205 31619 6239
rect 2973 6069 3007 6103
rect 3939 6069 3973 6103
rect 4629 6069 4663 6103
rect 5089 6069 5123 6103
rect 9597 6069 9631 6103
rect 9781 6069 9815 6103
rect 11161 6069 11195 6103
rect 11897 6069 11931 6103
rect 12173 6069 12207 6103
rect 15393 6069 15427 6103
rect 20085 6069 20119 6103
rect 21281 6069 21315 6103
rect 22845 6069 22879 6103
rect 23489 6069 23523 6103
rect 24961 6069 24995 6103
rect 26525 6137 26559 6171
rect 27169 6137 27203 6171
rect 27721 6137 27755 6171
rect 28457 6137 28491 6171
rect 31861 6137 31895 6171
rect 33425 6137 33459 6171
rect 34621 6137 34655 6171
rect 35081 6137 35115 6171
rect 35633 6137 35667 6171
rect 36553 6137 36587 6171
rect 36645 6137 36679 6171
rect 25605 6069 25639 6103
rect 26157 6069 26191 6103
rect 27997 6069 28031 6103
rect 29377 6069 29411 6103
rect 30389 6069 30423 6103
rect 33057 6069 33091 6103
rect 36277 6069 36311 6103
rect 3249 5865 3283 5899
rect 4997 5865 5031 5899
rect 7481 5865 7515 5899
rect 8033 5865 8067 5899
rect 8861 5865 8895 5899
rect 12817 5865 12851 5899
rect 14657 5865 14691 5899
rect 16221 5865 16255 5899
rect 17601 5865 17635 5899
rect 22201 5865 22235 5899
rect 22385 5865 22419 5899
rect 23765 5865 23799 5899
rect 24409 5865 24443 5899
rect 25237 5865 25271 5899
rect 29653 5865 29687 5899
rect 31217 5865 31251 5899
rect 33793 5865 33827 5899
rect 34253 5865 34287 5899
rect 34805 5865 34839 5899
rect 36645 5865 36679 5899
rect 1869 5797 1903 5831
rect 2282 5797 2316 5831
rect 4439 5797 4473 5831
rect 5089 5797 5123 5831
rect 5641 5797 5675 5831
rect 6285 5797 6319 5831
rect 9873 5797 9907 5831
rect 11891 5797 11925 5831
rect 13461 5797 13495 5831
rect 15025 5797 15059 5831
rect 16726 5797 16760 5831
rect 18797 5797 18831 5831
rect 20269 5797 20303 5831
rect 21097 5797 21131 5831
rect 21649 5797 21683 5831
rect 1961 5729 1995 5763
rect 2881 5729 2915 5763
rect 4077 5661 4111 5695
rect 23213 5797 23247 5831
rect 26709 5797 26743 5831
rect 28273 5797 28307 5831
rect 30659 5797 30693 5831
rect 32499 5797 32533 5831
rect 35817 5797 35851 5831
rect 5365 5729 5399 5763
rect 7665 5729 7699 5763
rect 8585 5729 8619 5763
rect 12449 5729 12483 5763
rect 15393 5729 15427 5763
rect 16405 5729 16439 5763
rect 17325 5729 17359 5763
rect 18429 5729 18463 5763
rect 22201 5729 22235 5763
rect 22753 5729 22787 5763
rect 22937 5729 22971 5763
rect 6193 5661 6227 5695
rect 6469 5661 6503 5695
rect 9413 5661 9447 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 11529 5661 11563 5695
rect 13369 5661 13403 5695
rect 17969 5661 18003 5695
rect 18705 5661 18739 5695
rect 19073 5661 19107 5695
rect 21005 5661 21039 5695
rect 24041 5661 24075 5695
rect 26617 5661 26651 5695
rect 27261 5661 27295 5695
rect 28181 5661 28215 5695
rect 28457 5661 28491 5695
rect 30297 5661 30331 5695
rect 32137 5661 32171 5695
rect 33885 5661 33919 5695
rect 35725 5661 35759 5695
rect 36001 5661 36035 5695
rect 13921 5593 13955 5627
rect 15577 5593 15611 5627
rect 35081 5593 35115 5627
rect 5089 5525 5123 5559
rect 10977 5525 11011 5559
rect 11345 5525 11379 5559
rect 14289 5525 14323 5559
rect 15853 5525 15887 5559
rect 19625 5525 19659 5559
rect 20637 5525 20671 5559
rect 21925 5525 21959 5559
rect 24961 5525 24995 5559
rect 29285 5525 29319 5559
rect 33057 5525 33091 5559
rect 35449 5525 35483 5559
rect 1593 5321 1627 5355
rect 5457 5321 5491 5355
rect 6469 5321 6503 5355
rect 7205 5321 7239 5355
rect 8585 5321 8619 5355
rect 8953 5321 8987 5355
rect 10425 5321 10459 5355
rect 12633 5321 12667 5355
rect 16405 5321 16439 5355
rect 17049 5321 17083 5355
rect 22017 5321 22051 5355
rect 23305 5321 23339 5355
rect 23397 5321 23431 5355
rect 26341 5321 26375 5355
rect 28089 5321 28123 5355
rect 28457 5321 28491 5355
rect 31033 5321 31067 5355
rect 34253 5321 34287 5355
rect 35909 5321 35943 5355
rect 6101 5253 6135 5287
rect 11621 5253 11655 5287
rect 11897 5253 11931 5287
rect 13461 5253 13495 5287
rect 21649 5253 21683 5287
rect 4537 5185 4571 5219
rect 4905 5185 4939 5219
rect 7665 5185 7699 5219
rect 9321 5185 9355 5219
rect 1409 5117 1443 5151
rect 1961 5117 1995 5151
rect 2697 5117 2731 5151
rect 3617 5117 3651 5151
rect 9505 5117 9539 5151
rect 9965 5117 9999 5151
rect 10885 5117 10919 5151
rect 11161 5117 11195 5151
rect 11529 5117 11563 5151
rect 12265 5185 12299 5219
rect 14841 5185 14875 5219
rect 15393 5185 15427 5219
rect 15669 5185 15703 5219
rect 19257 5185 19291 5219
rect 21097 5185 21131 5219
rect 23121 5185 23155 5219
rect 2513 5049 2547 5083
rect 3059 5049 3093 5083
rect 4169 5049 4203 5083
rect 4629 5049 4663 5083
rect 7573 5049 7607 5083
rect 8027 5049 8061 5083
rect 10977 5049 11011 5083
rect 11621 5049 11655 5083
rect 12081 5117 12115 5151
rect 12449 5117 12483 5151
rect 12909 5117 12943 5151
rect 13553 5117 13587 5151
rect 14473 5117 14507 5151
rect 15209 5117 15243 5151
rect 16865 5117 16899 5151
rect 18061 5117 18095 5151
rect 18521 5117 18555 5151
rect 24593 5253 24627 5287
rect 33241 5253 33275 5287
rect 36277 5253 36311 5287
rect 26065 5185 26099 5219
rect 26709 5185 26743 5219
rect 26985 5185 27019 5219
rect 27261 5185 27295 5219
rect 29653 5185 29687 5219
rect 32321 5185 32355 5219
rect 33977 5185 34011 5219
rect 34989 5185 35023 5219
rect 35357 5185 35391 5219
rect 36829 5185 36863 5219
rect 23673 5117 23707 5151
rect 30849 5117 30883 5151
rect 31309 5117 31343 5151
rect 33517 5117 33551 5151
rect 13915 5049 13949 5083
rect 15485 5049 15519 5083
rect 19165 5049 19199 5083
rect 19619 5049 19653 5083
rect 21189 5049 21223 5083
rect 23305 5049 23339 5083
rect 23994 5049 24028 5083
rect 24869 5049 24903 5083
rect 27077 5049 27111 5083
rect 29009 5049 29043 5083
rect 29377 5049 29411 5083
rect 29469 5049 29503 5083
rect 30389 5049 30423 5083
rect 31861 5049 31895 5083
rect 32229 5049 32263 5083
rect 32683 5049 32717 5083
rect 35081 5049 35115 5083
rect 36553 5049 36587 5083
rect 36645 5049 36679 5083
rect 9505 4981 9539 5015
rect 12081 4981 12115 5015
rect 17325 4981 17359 5015
rect 17693 4981 17727 5015
rect 18245 4981 18279 5015
rect 20177 4981 20211 5015
rect 20453 4981 20487 5015
rect 20821 4981 20855 5015
rect 22385 4981 22419 5015
rect 22569 4981 22603 5015
rect 25421 4981 25455 5015
rect 30665 4981 30699 5015
rect 34713 4981 34747 5015
rect 1685 4777 1719 4811
rect 3801 4777 3835 4811
rect 5825 4777 5859 4811
rect 7757 4777 7791 4811
rect 8217 4777 8251 4811
rect 12173 4777 12207 4811
rect 12449 4777 12483 4811
rect 12909 4777 12943 4811
rect 14013 4777 14047 4811
rect 14381 4777 14415 4811
rect 18061 4777 18095 4811
rect 19625 4777 19659 4811
rect 21925 4777 21959 4811
rect 24317 4777 24351 4811
rect 24961 4777 24995 4811
rect 26249 4777 26283 4811
rect 29285 4777 29319 4811
rect 32597 4777 32631 4811
rect 32965 4777 32999 4811
rect 34989 4777 35023 4811
rect 36093 4777 36127 4811
rect 36461 4777 36495 4811
rect 2139 4709 2173 4743
rect 4261 4709 4295 4743
rect 5089 4709 5123 4743
rect 9873 4709 9907 4743
rect 10425 4709 10459 4743
rect 11615 4709 11649 4743
rect 13185 4709 13219 4743
rect 13737 4709 13771 4743
rect 16865 4709 16899 4743
rect 19067 4709 19101 4743
rect 20729 4709 20763 4743
rect 21097 4709 21131 4743
rect 21649 4709 21683 4743
rect 24041 4709 24075 4743
rect 24685 4709 24719 4743
rect 26709 4709 26743 4743
rect 28273 4709 28307 4743
rect 33787 4709 33821 4743
rect 35449 4709 35483 4743
rect 6561 4641 6595 4675
rect 6745 4641 6779 4675
rect 8769 4641 8803 4675
rect 15301 4641 15335 4675
rect 15853 4641 15887 4675
rect 18705 4641 18739 4675
rect 20269 4641 20303 4675
rect 23397 4641 23431 4675
rect 23765 4641 23799 4675
rect 24869 4641 24903 4675
rect 25329 4641 25363 4675
rect 30481 4641 30515 4675
rect 31033 4641 31067 4675
rect 31217 4641 31251 4675
rect 1777 4573 1811 4607
rect 3525 4573 3559 4607
rect 4169 4573 4203 4607
rect 7021 4573 7055 4607
rect 7297 4573 7331 4607
rect 7849 4573 7883 4607
rect 9781 4573 9815 4607
rect 11253 4573 11287 4607
rect 13093 4573 13127 4607
rect 15669 4573 15703 4607
rect 16405 4573 16439 4607
rect 17233 4573 17267 4607
rect 21005 4573 21039 4607
rect 26617 4573 26651 4607
rect 28181 4573 28215 4607
rect 28457 4573 28491 4607
rect 32137 4573 32171 4607
rect 33425 4573 33459 4607
rect 35173 4573 35207 4607
rect 3065 4505 3099 4539
rect 4721 4505 4755 4539
rect 27169 4505 27203 4539
rect 2697 4437 2731 4471
rect 9045 4437 9079 4471
rect 9413 4437 9447 4471
rect 10885 4437 10919 4471
rect 15117 4437 15151 4471
rect 16681 4437 16715 4471
rect 17003 4437 17037 4471
rect 17141 4437 17175 4471
rect 17325 4437 17359 4471
rect 18429 4437 18463 4471
rect 19901 4437 19935 4471
rect 31493 4437 31527 4471
rect 34345 4437 34379 4471
rect 2513 4233 2547 4267
rect 5549 4233 5583 4267
rect 6377 4233 6411 4267
rect 7021 4233 7055 4267
rect 9229 4233 9263 4267
rect 16589 4233 16623 4267
rect 17325 4233 17359 4267
rect 18199 4233 18233 4267
rect 19165 4233 19199 4267
rect 20913 4233 20947 4267
rect 21281 4233 21315 4267
rect 23029 4233 23063 4267
rect 24777 4233 24811 4267
rect 25881 4233 25915 4267
rect 27629 4233 27663 4267
rect 28181 4233 28215 4267
rect 30941 4233 30975 4267
rect 32413 4233 32447 4267
rect 34621 4233 34655 4267
rect 35909 4233 35943 4267
rect 36277 4233 36311 4267
rect 36645 4233 36679 4267
rect 2145 4165 2179 4199
rect 3249 4165 3283 4199
rect 3985 4165 4019 4199
rect 5917 4165 5951 4199
rect 11345 4165 11379 4199
rect 11897 4165 11931 4199
rect 12725 4165 12759 4199
rect 16478 4165 16512 4199
rect 18337 4165 18371 4199
rect 21557 4165 21591 4199
rect 23305 4165 23339 4199
rect 24501 4165 24535 4199
rect 30481 4165 30515 4199
rect 33701 4165 33735 4199
rect 35541 4165 35575 4199
rect 2697 4097 2731 4131
rect 4261 4097 4295 4131
rect 7849 4097 7883 4131
rect 16681 4097 16715 4131
rect 17785 4097 17819 4131
rect 18429 4097 18463 4131
rect 18797 4097 18831 4131
rect 26525 4097 26559 4131
rect 31125 4097 31159 4131
rect 34989 4097 35023 4131
rect 1501 4029 1535 4063
rect 5733 4029 5767 4063
rect 6837 4029 6871 4063
rect 7389 4029 7423 4063
rect 9965 4029 9999 4063
rect 10701 4029 10735 4063
rect 11253 4029 11287 4063
rect 11437 4029 11471 4063
rect 13185 4029 13219 4063
rect 13553 4029 13587 4063
rect 13875 4029 13909 4063
rect 14289 4029 14323 4063
rect 15117 4029 15151 4063
rect 15485 4029 15519 4063
rect 17049 4029 17083 4063
rect 19441 4029 19475 4063
rect 19993 4029 20027 4063
rect 21741 4029 21775 4063
rect 22293 4029 22327 4063
rect 24961 4029 24995 4063
rect 26709 4029 26743 4063
rect 29377 4029 29411 4063
rect 29837 4029 29871 4063
rect 32597 4029 32631 4063
rect 33057 4029 33091 4063
rect 36461 4029 36495 4063
rect 37013 4029 37047 4063
rect 37600 4029 37634 4063
rect 38025 4029 38059 4063
rect 2789 3961 2823 3995
rect 3617 3961 3651 3995
rect 4353 3961 4387 3995
rect 4905 3961 4939 3995
rect 7757 3961 7791 3995
rect 8170 3961 8204 3995
rect 9597 3961 9631 3995
rect 14841 3961 14875 3995
rect 14933 3961 14967 3995
rect 15761 3961 15795 3995
rect 16313 3961 16347 3995
rect 18061 3961 18095 3995
rect 20314 3961 20348 3995
rect 25282 3961 25316 3995
rect 27071 3961 27105 3995
rect 30113 3961 30147 3995
rect 31217 3961 31251 3995
rect 31769 3961 31803 3995
rect 33333 3961 33367 3995
rect 35081 3961 35115 3995
rect 37703 3961 37737 3995
rect 1731 3893 1765 3927
rect 5273 3893 5307 3927
rect 8769 3893 8803 3927
rect 10333 3893 10367 3927
rect 12265 3893 12299 3927
rect 13553 3893 13587 3927
rect 16129 3893 16163 3927
rect 19809 3893 19843 3927
rect 22017 3893 22051 3927
rect 23673 3893 23707 3927
rect 26157 3893 26191 3927
rect 28457 3893 28491 3927
rect 29009 3893 29043 3927
rect 33977 3893 34011 3927
rect 2789 3689 2823 3723
rect 3157 3689 3191 3723
rect 3893 3689 3927 3723
rect 4169 3689 4203 3723
rect 5733 3689 5767 3723
rect 6929 3689 6963 3723
rect 7573 3689 7607 3723
rect 9137 3689 9171 3723
rect 9873 3689 9907 3723
rect 11069 3689 11103 3723
rect 13461 3689 13495 3723
rect 14105 3689 14139 3723
rect 14289 3689 14323 3723
rect 18981 3689 19015 3723
rect 22201 3689 22235 3723
rect 22753 3689 22787 3723
rect 23305 3689 23339 3723
rect 25145 3689 25179 3723
rect 25973 3689 26007 3723
rect 26249 3689 26283 3723
rect 28089 3689 28123 3723
rect 30113 3689 30147 3723
rect 31125 3689 31159 3723
rect 34621 3689 34655 3723
rect 1955 3621 1989 3655
rect 8217 3621 8251 3655
rect 13829 3621 13863 3655
rect 16405 3621 16439 3655
rect 18245 3621 18279 3655
rect 19901 3621 19935 3655
rect 20913 3621 20947 3655
rect 24225 3621 24259 3655
rect 24317 3621 24351 3655
rect 26801 3621 26835 3655
rect 27353 3621 27387 3655
rect 28502 3621 28536 3655
rect 30526 3621 30560 3655
rect 34022 3621 34056 3655
rect 35633 3621 35667 3655
rect 4077 3553 4111 3587
rect 4629 3553 4663 3587
rect 5733 3553 5767 3587
rect 6193 3553 6227 3587
rect 9689 3553 9723 3587
rect 11069 3553 11103 3587
rect 11621 3553 11655 3587
rect 11805 3553 11839 3587
rect 12817 3553 12851 3587
rect 14105 3553 14139 3587
rect 15669 3553 15703 3587
rect 15899 3553 15933 3587
rect 17049 3553 17083 3587
rect 17233 3553 17267 3587
rect 19165 3553 19199 3587
rect 19625 3553 19659 3587
rect 21097 3553 21131 3587
rect 22385 3553 22419 3587
rect 30205 3553 30239 3587
rect 32137 3553 32171 3587
rect 32597 3553 32631 3587
rect 33701 3553 33735 3587
rect 1593 3485 1627 3519
rect 8125 3485 8159 3519
rect 10517 3485 10551 3519
rect 12964 3485 12998 3519
rect 13185 3485 13219 3519
rect 16037 3485 16071 3519
rect 16865 3485 16899 3519
rect 17601 3485 17635 3519
rect 17969 3485 18003 3519
rect 21465 3485 21499 3519
rect 24501 3485 24535 3519
rect 26709 3485 26743 3519
rect 28181 3485 28215 3519
rect 32873 3485 32907 3519
rect 35173 3485 35207 3519
rect 35541 3485 35575 3519
rect 8677 3417 8711 3451
rect 15807 3417 15841 3451
rect 17049 3417 17083 3451
rect 17509 3417 17543 3451
rect 20177 3417 20211 3451
rect 20545 3417 20579 3451
rect 29101 3417 29135 3451
rect 36093 3417 36127 3451
rect 2513 3349 2547 3383
rect 5273 3349 5307 3383
rect 7941 3349 7975 3383
rect 9505 3349 9539 3383
rect 12541 3349 12575 3383
rect 13093 3349 13127 3383
rect 14657 3349 14691 3383
rect 15025 3349 15059 3383
rect 15577 3349 15611 3383
rect 17371 3349 17405 3383
rect 18613 3349 18647 3383
rect 21741 3349 21775 3383
rect 25513 3349 25547 3383
rect 29377 3349 29411 3383
rect 31493 3349 31527 3383
rect 1685 3145 1719 3179
rect 3709 3145 3743 3179
rect 4077 3145 4111 3179
rect 6285 3145 6319 3179
rect 8125 3145 8159 3179
rect 9873 3145 9907 3179
rect 10517 3145 10551 3179
rect 12265 3145 12299 3179
rect 13461 3145 13495 3179
rect 17785 3145 17819 3179
rect 20913 3145 20947 3179
rect 21281 3145 21315 3179
rect 21833 3145 21867 3179
rect 23029 3145 23063 3179
rect 23489 3145 23523 3179
rect 24225 3145 24259 3179
rect 26065 3145 26099 3179
rect 28641 3145 28675 3179
rect 30665 3145 30699 3179
rect 31861 3145 31895 3179
rect 32321 3145 32355 3179
rect 34069 3145 34103 3179
rect 34713 3145 34747 3179
rect 35909 3145 35943 3179
rect 36277 3145 36311 3179
rect 3157 3077 3191 3111
rect 4353 3077 4387 3111
rect 14105 3077 14139 3111
rect 16589 3077 16623 3111
rect 17233 3077 17267 3111
rect 18153 3077 18187 3111
rect 24501 3077 24535 3111
rect 24593 3077 24627 3111
rect 27169 3077 27203 3111
rect 30389 3077 30423 3111
rect 33701 3077 33735 3111
rect 35725 3077 35759 3111
rect 2237 3009 2271 3043
rect 2881 3009 2915 3043
rect 5089 3009 5123 3043
rect 10241 3009 10275 3043
rect 11437 3009 11471 3043
rect 11897 3009 11931 3043
rect 16037 3009 16071 3043
rect 18521 3009 18555 3043
rect 23765 3009 23799 3043
rect 4169 2941 4203 2975
rect 5181 2941 5215 2975
rect 5273 2941 5307 2975
rect 5457 2941 5491 2975
rect 6653 2941 6687 2975
rect 6837 2941 6871 2975
rect 7297 2941 7331 2975
rect 8493 2941 8527 2975
rect 8953 2941 8987 2975
rect 10793 2941 10827 2975
rect 12449 2941 12483 2975
rect 12541 2941 12575 2975
rect 12725 2941 12759 2975
rect 14013 2941 14047 2975
rect 14289 2941 14323 2975
rect 15577 2941 15611 2975
rect 15669 2941 15703 2975
rect 15853 2941 15887 2975
rect 18061 2941 18095 2975
rect 18337 2941 18371 2975
rect 19901 2941 19935 2975
rect 20085 2941 20119 2975
rect 22017 2941 22051 2975
rect 22569 2941 22603 2975
rect 26341 3009 26375 3043
rect 26617 3009 26651 3043
rect 30021 3009 30055 3043
rect 31585 3009 31619 3043
rect 33149 3009 33183 3043
rect 34989 3009 35023 3043
rect 35633 3009 35667 3043
rect 24777 2941 24811 2975
rect 28216 2941 28250 2975
rect 30849 2941 30883 2975
rect 31309 2941 31343 2975
rect 32413 2941 32447 2975
rect 32873 2941 32907 2975
rect 36461 3009 36495 3043
rect 37508 2941 37542 2975
rect 37933 2941 37967 2975
rect 2329 2873 2363 2907
rect 5917 2873 5951 2907
rect 15393 2873 15427 2907
rect 19073 2873 19107 2907
rect 19441 2873 19475 2907
rect 22753 2873 22787 2907
rect 24501 2873 24535 2907
rect 25098 2873 25132 2907
rect 26709 2873 26743 2907
rect 27537 2873 27571 2907
rect 28319 2873 28353 2907
rect 29377 2873 29411 2907
rect 29469 2873 29503 2907
rect 35081 2873 35115 2907
rect 35725 2873 35759 2907
rect 37611 2873 37645 2907
rect 2053 2805 2087 2839
rect 4721 2805 4755 2839
rect 6929 2805 6963 2839
rect 8861 2805 8895 2839
rect 9321 2805 9355 2839
rect 12909 2805 12943 2839
rect 13829 2805 13863 2839
rect 14473 2805 14507 2839
rect 15025 2805 15059 2839
rect 19717 2805 19751 2839
rect 25697 2805 25731 2839
rect 28089 2805 28123 2839
rect 29009 2805 29043 2839
rect 2053 2601 2087 2635
rect 5365 2601 5399 2635
rect 6377 2601 6411 2635
rect 7941 2601 7975 2635
rect 9229 2601 9263 2635
rect 9505 2601 9539 2635
rect 10885 2601 10919 2635
rect 13277 2601 13311 2635
rect 14105 2601 14139 2635
rect 15209 2601 15243 2635
rect 16957 2601 16991 2635
rect 17601 2601 17635 2635
rect 20085 2601 20119 2635
rect 21373 2601 21407 2635
rect 25053 2601 25087 2635
rect 25421 2601 25455 2635
rect 26341 2601 26375 2635
rect 28825 2601 28859 2635
rect 29561 2601 29595 2635
rect 32597 2601 32631 2635
rect 34069 2601 34103 2635
rect 34989 2601 35023 2635
rect 35909 2601 35943 2635
rect 2237 2533 2271 2567
rect 2329 2533 2363 2567
rect 2881 2533 2915 2567
rect 8861 2533 8895 2567
rect 9965 2533 9999 2567
rect 11253 2533 11287 2567
rect 12633 2533 12667 2567
rect 18337 2533 18371 2567
rect 19717 2533 19751 2567
rect 21741 2533 21775 2567
rect 22109 2533 22143 2567
rect 23121 2533 23155 2567
rect 27353 2533 27387 2567
rect 28181 2533 28215 2567
rect 29101 2533 29135 2567
rect 30481 2533 30515 2567
rect 30941 2533 30975 2567
rect 31769 2533 31803 2567
rect 4721 2465 4755 2499
rect 4905 2465 4939 2499
rect 5181 2465 5215 2499
rect 6745 2465 6779 2499
rect 6929 2465 6963 2499
rect 7665 2465 7699 2499
rect 8401 2465 8435 2499
rect 8585 2465 8619 2499
rect 11380 2465 11414 2499
rect 14197 2465 14231 2499
rect 15577 2465 15611 2499
rect 16589 2465 16623 2499
rect 17049 2465 17083 2499
rect 18061 2465 18095 2499
rect 18429 2465 18463 2499
rect 19901 2465 19935 2499
rect 21189 2465 21223 2499
rect 22385 2465 22419 2499
rect 22937 2465 22971 2499
rect 23857 2465 23891 2499
rect 24225 2465 24259 2499
rect 24501 2465 24535 2499
rect 25640 2465 25674 2499
rect 27445 2465 27479 2499
rect 27997 2465 28031 2499
rect 29745 2465 29779 2499
rect 30297 2465 30331 2499
rect 31344 2465 31378 2499
rect 33660 2465 33694 2499
rect 35516 2465 35550 2499
rect 36528 2465 36562 2499
rect 36921 2465 36955 2499
rect 3157 2397 3191 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 12081 2397 12115 2431
rect 13001 2397 13035 2431
rect 13829 2397 13863 2431
rect 20913 2397 20947 2431
rect 23397 2397 23431 2431
rect 24777 2397 24811 2431
rect 31447 2397 31481 2431
rect 31953 2397 31987 2431
rect 33747 2397 33781 2431
rect 1685 2329 1719 2363
rect 4997 2329 5031 2363
rect 5917 2329 5951 2363
rect 7113 2329 7147 2363
rect 12449 2329 12483 2363
rect 17233 2329 17267 2363
rect 20545 2329 20579 2363
rect 26617 2329 26651 2363
rect 32137 2329 32171 2363
rect 33057 2329 33091 2363
rect 35587 2329 35621 2363
rect 4445 2261 4479 2295
rect 11483 2261 11517 2295
rect 12771 2261 12805 2295
rect 12909 2261 12943 2295
rect 13645 2261 13679 2295
rect 13829 2261 13863 2295
rect 14381 2261 14415 2295
rect 14841 2261 14875 2295
rect 15761 2261 15795 2295
rect 25743 2261 25777 2295
rect 31953 2261 31987 2295
rect 36599 2261 36633 2295
<< metal1 >>
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 106 12928 112 12980
rect 164 12968 170 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 164 12940 1593 12968
rect 164 12928 170 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 35621 12971 35679 12977
rect 35621 12937 35633 12971
rect 35667 12968 35679 12971
rect 39574 12968 39580 12980
rect 35667 12940 39580 12968
rect 35667 12937 35679 12940
rect 35621 12931 35679 12937
rect 39574 12928 39580 12940
rect 39632 12928 39638 12980
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12733 1455 12767
rect 1397 12727 1455 12733
rect 2568 12767 2626 12773
rect 2568 12733 2580 12767
rect 2614 12764 2626 12767
rect 2777 12767 2835 12773
rect 2777 12764 2789 12767
rect 2614 12736 2789 12764
rect 2614 12733 2626 12736
rect 2568 12727 2626 12733
rect 2777 12733 2789 12736
rect 2823 12733 2835 12767
rect 2777 12727 2835 12733
rect 4960 12767 5018 12773
rect 4960 12733 4972 12767
rect 5006 12764 5018 12767
rect 12989 12767 13047 12773
rect 5006 12736 5488 12764
rect 5006 12733 5018 12736
rect 4960 12727 5018 12733
rect 1412 12696 1440 12727
rect 2041 12699 2099 12705
rect 2041 12696 2053 12699
rect 1412 12668 2053 12696
rect 2041 12665 2053 12668
rect 2087 12696 2099 12699
rect 5350 12696 5356 12708
rect 2087 12668 5356 12696
rect 2087 12665 2099 12668
rect 2041 12659 2099 12665
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 5460 12640 5488 12736
rect 12989 12733 13001 12767
rect 13035 12764 13047 12767
rect 13449 12767 13507 12773
rect 13449 12764 13461 12767
rect 13035 12736 13461 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 13449 12733 13461 12736
rect 13495 12764 13507 12767
rect 16758 12764 16764 12776
rect 13495 12736 16764 12764
rect 13495 12733 13507 12736
rect 13449 12727 13507 12733
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 32214 12724 32220 12776
rect 32272 12764 32278 12776
rect 35437 12767 35495 12773
rect 35437 12764 35449 12767
rect 32272 12736 35449 12764
rect 32272 12724 32278 12736
rect 35437 12733 35449 12736
rect 35483 12764 35495 12767
rect 35989 12767 36047 12773
rect 35989 12764 36001 12767
rect 35483 12736 36001 12764
rect 35483 12733 35495 12736
rect 35437 12727 35495 12733
rect 35989 12733 36001 12736
rect 36035 12733 36047 12767
rect 35989 12727 36047 12733
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 2639 12631 2697 12637
rect 2639 12628 2651 12631
rect 1636 12600 2651 12628
rect 1636 12588 1642 12600
rect 2639 12597 2651 12600
rect 2685 12597 2697 12631
rect 2639 12591 2697 12597
rect 2777 12631 2835 12637
rect 2777 12597 2789 12631
rect 2823 12628 2835 12631
rect 3053 12631 3111 12637
rect 3053 12628 3065 12631
rect 2823 12600 3065 12628
rect 2823 12597 2835 12600
rect 2777 12591 2835 12597
rect 3053 12597 3065 12600
rect 3099 12628 3111 12631
rect 3786 12628 3792 12640
rect 3099 12600 3792 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 5031 12631 5089 12637
rect 5031 12597 5043 12631
rect 5077 12628 5089 12631
rect 5166 12628 5172 12640
rect 5077 12600 5172 12628
rect 5077 12597 5089 12600
rect 5031 12591 5089 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 5442 12628 5448 12640
rect 5403 12600 5448 12628
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 11882 12588 11888 12640
rect 11940 12628 11946 12640
rect 13173 12631 13231 12637
rect 13173 12628 13185 12631
rect 11940 12600 13185 12628
rect 11940 12588 11946 12600
rect 13173 12597 13185 12600
rect 13219 12597 13231 12631
rect 13173 12591 13231 12597
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1026 12384 1032 12436
rect 1084 12424 1090 12436
rect 1581 12427 1639 12433
rect 1581 12424 1593 12427
rect 1084 12396 1593 12424
rect 1084 12384 1090 12396
rect 1581 12393 1593 12396
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 5350 12316 5356 12368
rect 5408 12356 5414 12368
rect 5408 12328 11351 12356
rect 5408 12316 5414 12328
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 2498 12288 2504 12300
rect 2459 12260 2504 12288
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 4111 12291 4169 12297
rect 4111 12257 4123 12291
rect 4157 12257 4169 12291
rect 4111 12251 4169 12257
rect 5972 12291 6030 12297
rect 5972 12257 5984 12291
rect 6018 12288 6030 12291
rect 6178 12288 6184 12300
rect 6018 12260 6184 12288
rect 6018 12257 6030 12260
rect 5972 12251 6030 12257
rect 106 12112 112 12164
rect 164 12152 170 12164
rect 2685 12155 2743 12161
rect 2685 12152 2697 12155
rect 164 12124 2697 12152
rect 164 12112 170 12124
rect 2685 12121 2697 12124
rect 2731 12121 2743 12155
rect 4126 12152 4154 12251
rect 6178 12248 6184 12260
rect 6236 12248 6242 12300
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10502 12288 10508 12300
rect 10275 12260 10508 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 11323 12297 11351 12328
rect 11308 12291 11366 12297
rect 11308 12257 11320 12291
rect 11354 12288 11366 12291
rect 12250 12288 12256 12300
rect 11354 12260 12256 12288
rect 11354 12257 11366 12260
rect 11308 12251 11366 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13446 12288 13452 12300
rect 13127 12260 13452 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 4614 12152 4620 12164
rect 4126 12124 4620 12152
rect 2685 12115 2743 12121
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12084 2099 12087
rect 2130 12084 2136 12096
rect 2087 12056 2136 12084
rect 2087 12053 2099 12056
rect 2041 12047 2099 12053
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 2314 12084 2320 12096
rect 2275 12056 2320 12084
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 4203 12087 4261 12093
rect 4203 12053 4215 12087
rect 4249 12084 4261 12087
rect 4338 12084 4344 12096
rect 4249 12056 4344 12084
rect 4249 12053 4261 12056
rect 4203 12047 4261 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 6043 12087 6101 12093
rect 6043 12053 6055 12087
rect 6089 12084 6101 12087
rect 7466 12084 7472 12096
rect 6089 12056 7472 12084
rect 6089 12053 6101 12056
rect 6043 12047 6101 12053
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 10410 12084 10416 12096
rect 10371 12056 10416 12084
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 11379 12087 11437 12093
rect 11379 12053 11391 12087
rect 11425 12084 11437 12087
rect 11790 12084 11796 12096
rect 11425 12056 11796 12084
rect 11425 12053 11437 12056
rect 11379 12047 11437 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 14090 12084 14096 12096
rect 13311 12056 14096 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 14274 12084 14280 12096
rect 14235 12056 14280 12084
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 2961 11883 3019 11889
rect 2961 11880 2973 11883
rect 2556 11852 2973 11880
rect 2556 11840 2562 11852
rect 2961 11849 2973 11852
rect 3007 11880 3019 11883
rect 5442 11880 5448 11892
rect 3007 11852 5448 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 14090 11880 14096 11892
rect 5592 11852 8524 11880
rect 14051 11852 14096 11880
rect 5592 11840 5598 11852
rect 14 11772 20 11824
rect 72 11812 78 11824
rect 3605 11815 3663 11821
rect 3605 11812 3617 11815
rect 72 11784 3617 11812
rect 72 11772 78 11784
rect 3605 11781 3617 11784
rect 3651 11781 3663 11815
rect 3605 11775 3663 11781
rect 3694 11772 3700 11824
rect 3752 11812 3758 11824
rect 6641 11815 6699 11821
rect 6641 11812 6653 11815
rect 3752 11784 6653 11812
rect 3752 11772 3758 11784
rect 6641 11781 6653 11784
rect 6687 11781 6699 11815
rect 6641 11775 6699 11781
rect 1394 11704 1400 11756
rect 1452 11744 1458 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1452 11716 1685 11744
rect 1452 11704 1458 11716
rect 1673 11713 1685 11716
rect 1719 11744 1731 11747
rect 7098 11744 7104 11756
rect 1719 11716 7104 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 8496 11744 8524 11852
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 10413 11815 10471 11821
rect 10413 11781 10425 11815
rect 10459 11812 10471 11815
rect 15470 11812 15476 11824
rect 10459 11784 15476 11812
rect 10459 11781 10471 11784
rect 10413 11775 10471 11781
rect 15470 11772 15476 11784
rect 15528 11772 15534 11824
rect 8496 11716 11351 11744
rect 2130 11676 2136 11688
rect 2091 11648 2136 11676
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 2314 11676 2320 11688
rect 2275 11648 2320 11676
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3375 11648 3433 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3421 11645 3433 11648
rect 3467 11676 3479 11679
rect 4706 11676 4712 11688
rect 3467 11648 4712 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 4890 11676 4896 11688
rect 4854 11648 4896 11676
rect 4890 11636 4896 11648
rect 4948 11685 4954 11688
rect 4948 11679 5002 11685
rect 4948 11645 4956 11679
rect 4990 11676 5002 11679
rect 5353 11679 5411 11685
rect 5353 11676 5365 11679
rect 4990 11648 5365 11676
rect 4990 11645 5002 11648
rect 4948 11639 5002 11645
rect 5353 11645 5365 11648
rect 5399 11676 5411 11679
rect 5534 11676 5540 11688
rect 5399 11648 5540 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 4948 11636 4954 11639
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 6876 11679 6934 11685
rect 6876 11676 6888 11679
rect 6687 11648 6888 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 6876 11645 6888 11648
rect 6922 11676 6934 11679
rect 10229 11679 10287 11685
rect 6922 11648 7420 11676
rect 6922 11645 6934 11648
rect 6876 11639 6934 11645
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 5031 11611 5089 11617
rect 5031 11608 5043 11611
rect 4120 11580 5043 11608
rect 4120 11568 4126 11580
rect 5031 11577 5043 11580
rect 5077 11577 5089 11611
rect 5031 11571 5089 11577
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 6963 11611 7021 11617
rect 6963 11608 6975 11611
rect 5500 11580 6975 11608
rect 5500 11568 5506 11580
rect 6963 11577 6975 11580
rect 7009 11577 7021 11611
rect 6963 11571 7021 11577
rect 7392 11552 7420 11648
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 10594 11676 10600 11688
rect 10275 11648 10600 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 10594 11636 10600 11648
rect 10652 11676 10658 11688
rect 11323 11685 11351 11716
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10652 11648 11069 11676
rect 10652 11636 10658 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11308 11679 11366 11685
rect 11308 11645 11320 11679
rect 11354 11676 11366 11679
rect 11354 11648 11836 11676
rect 11354 11645 11366 11648
rect 11308 11639 11366 11645
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2133 11543 2191 11549
rect 2133 11540 2145 11543
rect 2096 11512 2145 11540
rect 2096 11500 2102 11512
rect 2133 11509 2145 11512
rect 2179 11509 2191 11543
rect 2133 11503 2191 11509
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 4614 11540 4620 11552
rect 4203 11512 4620 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6178 11540 6184 11552
rect 6043 11512 6184 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 7374 11540 7380 11552
rect 7335 11512 7380 11540
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 10560 11512 10701 11540
rect 10560 11500 10566 11512
rect 10689 11509 10701 11512
rect 10735 11509 10747 11543
rect 10689 11503 10747 11509
rect 11379 11543 11437 11549
rect 11379 11509 11391 11543
rect 11425 11540 11437 11543
rect 11514 11540 11520 11552
rect 11425 11512 11520 11540
rect 11425 11509 11437 11512
rect 11379 11503 11437 11509
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 11808 11549 11836 11648
rect 13354 11636 13360 11688
rect 13412 11676 13418 11688
rect 14274 11676 14280 11688
rect 13412 11648 14280 11676
rect 13412 11636 13418 11648
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14737 11679 14795 11685
rect 14737 11645 14749 11679
rect 14783 11645 14795 11679
rect 14737 11639 14795 11645
rect 12161 11611 12219 11617
rect 12161 11577 12173 11611
rect 12207 11608 12219 11611
rect 12250 11608 12256 11620
rect 12207 11580 12256 11608
rect 12207 11577 12219 11580
rect 12161 11571 12219 11577
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 14090 11568 14096 11620
rect 14148 11608 14154 11620
rect 14752 11608 14780 11639
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 18484 11679 18542 11685
rect 18484 11676 18496 11679
rect 17368 11648 18496 11676
rect 17368 11636 17374 11648
rect 18484 11645 18496 11648
rect 18530 11676 18542 11679
rect 19242 11676 19248 11688
rect 18530 11648 19248 11676
rect 18530 11645 18542 11648
rect 18484 11639 18542 11645
rect 19242 11636 19248 11648
rect 19300 11636 19306 11688
rect 19740 11679 19798 11685
rect 19740 11676 19752 11679
rect 19622 11648 19752 11676
rect 15010 11608 15016 11620
rect 14148 11580 14780 11608
rect 14971 11580 15016 11608
rect 14148 11568 14154 11580
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 15746 11568 15752 11620
rect 15804 11608 15810 11620
rect 19622 11608 19650 11648
rect 19740 11645 19752 11648
rect 19786 11676 19798 11679
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 19786 11648 20177 11676
rect 19786 11645 19798 11648
rect 19740 11639 19798 11645
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 15804 11580 19650 11608
rect 19843 11611 19901 11617
rect 15804 11568 15810 11580
rect 19843 11577 19855 11611
rect 19889 11608 19901 11611
rect 22002 11608 22008 11620
rect 19889 11580 22008 11608
rect 19889 11577 19901 11580
rect 19843 11571 19901 11577
rect 22002 11568 22008 11580
rect 22060 11568 22066 11620
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 12066 11540 12072 11552
rect 11839 11512 12072 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12434 11540 12440 11552
rect 12395 11512 12440 11540
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13446 11540 13452 11552
rect 13219 11512 13452 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 18555 11543 18613 11549
rect 18555 11509 18567 11543
rect 18601 11540 18613 11543
rect 18782 11540 18788 11552
rect 18601 11512 18788 11540
rect 18601 11509 18613 11512
rect 18555 11503 18613 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 18969 11543 19027 11549
rect 18969 11509 18981 11543
rect 19015 11540 19027 11543
rect 19242 11540 19248 11552
rect 19015 11512 19248 11540
rect 19015 11509 19027 11512
rect 18969 11503 19027 11509
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 16991 11339 17049 11345
rect 16991 11305 17003 11339
rect 17037 11336 17049 11339
rect 19518 11336 19524 11348
rect 17037 11308 19524 11336
rect 17037 11305 17049 11308
rect 16991 11299 17049 11305
rect 19518 11296 19524 11308
rect 19576 11296 19582 11348
rect 35618 11336 35624 11348
rect 35579 11308 35624 11336
rect 35618 11296 35624 11308
rect 35676 11296 35682 11348
rect 4706 11228 4712 11280
rect 4764 11268 4770 11280
rect 4764 11240 7282 11268
rect 4764 11228 4770 11240
rect 1762 11160 1768 11212
rect 1820 11200 1826 11212
rect 1857 11203 1915 11209
rect 1857 11200 1869 11203
rect 1820 11172 1869 11200
rect 1820 11160 1826 11172
rect 1857 11169 1869 11172
rect 1903 11169 1915 11203
rect 2314 11200 2320 11212
rect 2275 11172 2320 11200
rect 1857 11163 1915 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4100 11203 4158 11209
rect 4100 11200 4112 11203
rect 3936 11172 4112 11200
rect 3936 11160 3942 11172
rect 4100 11169 4112 11172
rect 4146 11169 4158 11203
rect 4100 11163 4158 11169
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 5144 11203 5202 11209
rect 5144 11200 5156 11203
rect 4663 11172 5156 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 5144 11169 5156 11172
rect 5190 11200 5202 11203
rect 5258 11200 5264 11212
rect 5190 11172 5264 11200
rect 5190 11169 5202 11172
rect 5144 11163 5202 11169
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 6086 11200 6092 11212
rect 6047 11172 6092 11200
rect 6086 11160 6092 11172
rect 6144 11160 6150 11212
rect 7098 11200 7104 11212
rect 7059 11172 7104 11200
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7254 11200 7282 11240
rect 8180 11203 8238 11209
rect 8180 11200 8192 11203
rect 7254 11172 8192 11200
rect 8180 11169 8192 11172
rect 8226 11200 8238 11203
rect 8570 11200 8576 11212
rect 8226 11172 8576 11200
rect 8226 11169 8238 11172
rect 8180 11163 8238 11169
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10756 11203 10814 11209
rect 10756 11169 10768 11203
rect 10802 11200 10814 11203
rect 11238 11200 11244 11212
rect 10802 11172 11244 11200
rect 10802 11169 10814 11172
rect 10756 11163 10814 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11756 11172 11805 11200
rect 11756 11160 11762 11172
rect 11793 11169 11805 11172
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 13630 11200 13636 11212
rect 13587 11172 13636 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14090 11200 14096 11212
rect 14051 11172 14096 11200
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 16888 11203 16946 11209
rect 16888 11200 16900 11203
rect 16724 11172 16900 11200
rect 16724 11160 16730 11172
rect 16888 11169 16900 11172
rect 16934 11169 16946 11203
rect 16888 11163 16946 11169
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 18506 11200 18512 11212
rect 18371 11172 18512 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 19426 11200 19432 11212
rect 19387 11172 19432 11200
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 22072 11203 22130 11209
rect 22072 11169 22084 11203
rect 22118 11200 22130 11203
rect 22646 11200 22652 11212
rect 22118 11172 22652 11200
rect 22118 11169 22130 11172
rect 22072 11163 22130 11169
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 26672 11203 26730 11209
rect 26672 11169 26684 11203
rect 26718 11200 26730 11203
rect 26970 11200 26976 11212
rect 26718 11172 26976 11200
rect 26718 11169 26730 11172
rect 26672 11163 26730 11169
rect 26970 11160 26976 11172
rect 27028 11160 27034 11212
rect 34146 11160 34152 11212
rect 34204 11200 34210 11212
rect 34400 11203 34458 11209
rect 34400 11200 34412 11203
rect 34204 11172 34412 11200
rect 34204 11160 34210 11172
rect 34400 11169 34412 11172
rect 34446 11200 34458 11203
rect 34606 11200 34612 11212
rect 34446 11172 34612 11200
rect 34446 11169 34458 11172
rect 34400 11163 34458 11169
rect 34606 11160 34612 11172
rect 34664 11160 34670 11212
rect 35434 11200 35440 11212
rect 35395 11172 35440 11200
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2280 11104 2421 11132
rect 2280 11092 2286 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 12802 11132 12808 11144
rect 12483 11104 12808 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 15194 11132 15200 11144
rect 14415 11104 15200 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15654 11132 15660 11144
rect 15615 11104 15660 11132
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 3602 11024 3608 11076
rect 3660 11064 3666 11076
rect 5215 11067 5273 11073
rect 5215 11064 5227 11067
rect 3660 11036 5227 11064
rect 3660 11024 3666 11036
rect 5215 11033 5227 11036
rect 5261 11033 5273 11067
rect 5215 11027 5273 11033
rect 6454 11024 6460 11076
rect 6512 11064 6518 11076
rect 8251 11067 8309 11073
rect 8251 11064 8263 11067
rect 6512 11036 8263 11064
rect 6512 11024 6518 11036
rect 8251 11033 8263 11036
rect 8297 11033 8309 11067
rect 8251 11027 8309 11033
rect 9861 11067 9919 11073
rect 9861 11033 9873 11067
rect 9907 11064 9919 11067
rect 12158 11064 12164 11076
rect 9907 11036 12164 11064
rect 9907 11033 9919 11036
rect 9861 11027 9919 11033
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 1762 10996 1768 11008
rect 1723 10968 1768 10996
rect 1762 10956 1768 10968
rect 1820 10956 1826 11008
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 4203 10999 4261 11005
rect 4203 10996 4215 10999
rect 3568 10968 4215 10996
rect 3568 10956 3574 10968
rect 4203 10965 4215 10968
rect 4249 10965 4261 10999
rect 4203 10959 4261 10965
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 6227 10999 6285 11005
rect 6227 10996 6239 10999
rect 4856 10968 6239 10996
rect 4856 10956 4862 10968
rect 6227 10965 6239 10968
rect 6273 10965 6285 10999
rect 6227 10959 6285 10965
rect 6362 10956 6368 11008
rect 6420 10996 6426 11008
rect 7239 10999 7297 11005
rect 7239 10996 7251 10999
rect 6420 10968 7251 10996
rect 6420 10956 6426 10968
rect 7239 10965 7251 10968
rect 7285 10965 7297 10999
rect 7239 10959 7297 10965
rect 10827 10999 10885 11005
rect 10827 10965 10839 10999
rect 10873 10996 10885 10999
rect 13078 10996 13084 11008
rect 10873 10968 13084 10996
rect 10873 10965 10885 10968
rect 10827 10959 10885 10965
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 18555 10999 18613 11005
rect 18555 10965 18567 10999
rect 18601 10996 18613 10999
rect 18966 10996 18972 11008
rect 18601 10968 18972 10996
rect 18601 10965 18613 10968
rect 18555 10959 18613 10965
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 19567 10999 19625 11005
rect 19567 10965 19579 10999
rect 19613 10996 19625 10999
rect 19794 10996 19800 11008
rect 19613 10968 19800 10996
rect 19613 10965 19625 10968
rect 19567 10959 19625 10965
rect 19794 10956 19800 10968
rect 19852 10956 19858 11008
rect 22143 10999 22201 11005
rect 22143 10965 22155 10999
rect 22189 10996 22201 10999
rect 24486 10996 24492 11008
rect 22189 10968 24492 10996
rect 22189 10965 22201 10968
rect 22143 10959 22201 10965
rect 24486 10956 24492 10968
rect 24544 10956 24550 11008
rect 26743 10999 26801 11005
rect 26743 10965 26755 10999
rect 26789 10996 26801 10999
rect 29086 10996 29092 11008
rect 26789 10968 29092 10996
rect 26789 10965 26801 10968
rect 26743 10959 26801 10965
rect 29086 10956 29092 10968
rect 29144 10956 29150 11008
rect 34471 10999 34529 11005
rect 34471 10965 34483 10999
rect 34517 10996 34529 10999
rect 36170 10996 36176 11008
rect 34517 10968 36176 10996
rect 34517 10965 34529 10968
rect 34471 10959 34529 10965
rect 36170 10956 36176 10968
rect 36228 10956 36234 11008
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 934 10752 940 10804
rect 992 10792 998 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 992 10764 1593 10792
rect 992 10752 998 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 4522 10792 4528 10804
rect 4483 10764 4528 10792
rect 1581 10755 1639 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5258 10792 5264 10804
rect 5215 10764 5264 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5859 10795 5917 10801
rect 5859 10761 5871 10795
rect 5905 10792 5917 10795
rect 6270 10792 6276 10804
rect 5905 10764 6276 10792
rect 5905 10761 5917 10764
rect 5859 10755 5917 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 10468 10764 15301 10792
rect 10468 10752 10474 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 18506 10792 18512 10804
rect 18467 10764 18512 10792
rect 15289 10755 15347 10761
rect 11606 10684 11612 10736
rect 11664 10724 11670 10736
rect 13725 10727 13783 10733
rect 13725 10724 13737 10727
rect 11664 10696 13737 10724
rect 11664 10684 11670 10696
rect 13725 10693 13737 10696
rect 13771 10724 13783 10727
rect 14090 10724 14096 10736
rect 13771 10696 14096 10724
rect 13771 10693 13783 10696
rect 13725 10687 13783 10693
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 2685 10659 2743 10665
rect 2685 10656 2697 10659
rect 2188 10628 2697 10656
rect 2188 10616 2194 10628
rect 2685 10625 2697 10628
rect 2731 10656 2743 10659
rect 2731 10628 3372 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3344 10600 3372 10628
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7558 10656 7564 10668
rect 7156 10628 7564 10656
rect 7156 10616 7162 10628
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8570 10656 8576 10668
rect 8483 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10656 8634 10668
rect 11238 10656 11244 10668
rect 8628 10628 11244 10656
rect 8628 10616 8634 10628
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11394 10628 11805 10656
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 1412 10520 1440 10551
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 2777 10591 2835 10597
rect 2777 10588 2789 10591
rect 2556 10560 2789 10588
rect 2556 10548 2562 10560
rect 2777 10557 2789 10560
rect 2823 10557 2835 10591
rect 3326 10588 3332 10600
rect 3287 10560 3332 10588
rect 2777 10551 2835 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 5258 10588 5264 10600
rect 4387 10560 5264 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 5626 10588 5632 10600
rect 5587 10560 5632 10588
rect 5626 10548 5632 10560
rect 5684 10588 5690 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 5684 10560 6561 10588
rect 5684 10548 5690 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8067 10560 8892 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 2041 10523 2099 10529
rect 2041 10520 2053 10523
rect 1412 10492 2053 10520
rect 2041 10489 2053 10492
rect 2087 10520 2099 10523
rect 3970 10520 3976 10532
rect 2087 10492 3976 10520
rect 2087 10489 2099 10492
rect 2041 10483 2099 10489
rect 3970 10480 3976 10492
rect 4028 10480 4034 10532
rect 8864 10464 8892 10560
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 11394 10597 11422 10628
rect 11793 10625 11805 10628
rect 11839 10656 11851 10659
rect 12894 10656 12900 10668
rect 11839 10628 12900 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 14108 10656 14136 10684
rect 14108 10628 14596 10656
rect 10356 10591 10414 10597
rect 10356 10588 10368 10591
rect 9548 10560 10368 10588
rect 9548 10548 9554 10560
rect 10356 10557 10368 10560
rect 10402 10588 10414 10591
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10402 10560 10793 10588
rect 10402 10557 10414 10560
rect 10356 10551 10414 10557
rect 10781 10557 10793 10560
rect 10827 10588 10839 10591
rect 11368 10591 11426 10597
rect 11368 10588 11380 10591
rect 10827 10560 11380 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 11368 10557 11380 10560
rect 11414 10557 11426 10591
rect 11368 10551 11426 10557
rect 11471 10591 11529 10597
rect 11471 10557 11483 10591
rect 11517 10588 11529 10591
rect 12250 10588 12256 10600
rect 11517 10560 12256 10588
rect 11517 10557 11529 10560
rect 11471 10551 11529 10557
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12452 10560 12541 10588
rect 10459 10523 10517 10529
rect 10459 10489 10471 10523
rect 10505 10520 10517 10523
rect 12342 10520 12348 10532
rect 10505 10492 12348 10520
rect 10505 10489 10517 10492
rect 10459 10483 10517 10489
rect 12342 10480 12348 10492
rect 12400 10480 12406 10532
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 2869 10455 2927 10461
rect 2869 10452 2881 10455
rect 2832 10424 2881 10452
rect 2832 10412 2838 10424
rect 2869 10421 2881 10424
rect 2915 10421 2927 10455
rect 2869 10415 2927 10421
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 3936 10424 4077 10452
rect 3936 10412 3942 10424
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 6086 10452 6092 10464
rect 4580 10424 6092 10452
rect 4580 10412 4586 10424
rect 6086 10412 6092 10424
rect 6144 10452 6150 10464
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 6144 10424 6193 10452
rect 6144 10412 6150 10424
rect 6181 10421 6193 10424
rect 6227 10421 6239 10455
rect 6181 10415 6239 10421
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10452 7067 10455
rect 7282 10452 7288 10464
rect 7055 10424 7288 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8846 10452 8852 10464
rect 8807 10424 8852 10452
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9306 10452 9312 10464
rect 9267 10424 9312 10452
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9732 10424 9873 10452
rect 9732 10412 9738 10424
rect 9861 10421 9873 10424
rect 9907 10452 9919 10455
rect 10226 10452 10232 10464
rect 9907 10424 10232 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 11238 10452 11244 10464
rect 11199 10424 11244 10452
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 12124 10424 12173 10452
rect 12124 10412 12130 10424
rect 12161 10421 12173 10424
rect 12207 10452 12219 10455
rect 12452 10452 12480 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 14182 10588 14188 10600
rect 14143 10560 14188 10588
rect 12529 10551 12587 10557
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 14568 10597 14596 10628
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10557 14611 10591
rect 15304 10588 15332 10755
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 22646 10792 22652 10804
rect 22607 10764 22652 10792
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 26234 10792 26240 10804
rect 26195 10764 26240 10792
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 35345 10795 35403 10801
rect 35345 10761 35357 10795
rect 35391 10792 35403 10795
rect 35434 10792 35440 10804
rect 35391 10764 35440 10792
rect 35391 10761 35403 10764
rect 35345 10755 35403 10761
rect 35434 10752 35440 10764
rect 35492 10752 35498 10804
rect 35618 10724 35624 10736
rect 35579 10696 35624 10724
rect 35618 10684 35624 10696
rect 35676 10684 35682 10736
rect 17678 10656 17684 10668
rect 15856 10628 17684 10656
rect 15856 10597 15884 10628
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 18877 10659 18935 10665
rect 18877 10656 18889 10659
rect 17972 10628 18889 10656
rect 17972 10600 18000 10628
rect 18877 10625 18889 10628
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 19300 10628 21097 10656
rect 19300 10616 19306 10628
rect 15841 10591 15899 10597
rect 15841 10588 15853 10591
rect 15304 10560 15853 10588
rect 14553 10551 14611 10557
rect 15841 10557 15853 10560
rect 15887 10557 15899 10591
rect 15841 10551 15899 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 16482 10588 16488 10600
rect 16439 10560 16488 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 14826 10520 14832 10532
rect 14787 10492 14832 10520
rect 14826 10480 14832 10492
rect 14884 10480 14890 10532
rect 15749 10523 15807 10529
rect 15749 10489 15761 10523
rect 15795 10520 15807 10523
rect 16408 10520 16436 10551
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 17954 10588 17960 10600
rect 17915 10560 17960 10588
rect 17954 10548 17960 10560
rect 18012 10548 18018 10600
rect 18322 10548 18328 10600
rect 18380 10588 18386 10600
rect 19096 10591 19154 10597
rect 19096 10588 19108 10591
rect 18380 10560 19108 10588
rect 18380 10548 18386 10560
rect 19096 10557 19108 10560
rect 19142 10588 19154 10591
rect 19889 10591 19947 10597
rect 19889 10588 19901 10591
rect 19142 10560 19901 10588
rect 19142 10557 19154 10560
rect 19096 10551 19154 10557
rect 19889 10557 19901 10560
rect 19935 10588 19947 10591
rect 20254 10588 20260 10600
rect 19935 10560 20260 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20254 10548 20260 10560
rect 20312 10548 20318 10600
rect 20891 10597 20919 10628
rect 21085 10625 21097 10628
rect 21131 10625 21143 10659
rect 28074 10656 28080 10668
rect 21085 10619 21143 10625
rect 22296 10628 28080 10656
rect 22296 10597 22324 10628
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 35342 10616 35348 10668
rect 35400 10616 35406 10668
rect 20860 10591 20919 10597
rect 20860 10557 20872 10591
rect 20906 10560 20919 10591
rect 21856 10591 21914 10597
rect 21856 10588 21868 10591
rect 20951 10560 21868 10588
rect 20906 10557 20918 10560
rect 20860 10551 20918 10557
rect 16574 10520 16580 10532
rect 15795 10492 16436 10520
rect 16535 10492 16580 10520
rect 15795 10489 15807 10492
rect 15749 10483 15807 10489
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 18598 10480 18604 10532
rect 18656 10520 18662 10532
rect 19199 10523 19257 10529
rect 19199 10520 19211 10523
rect 18656 10492 19211 10520
rect 18656 10480 18662 10492
rect 19199 10489 19211 10492
rect 19245 10489 19257 10523
rect 20951 10520 20979 10560
rect 21856 10557 21868 10560
rect 21902 10588 21914 10591
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 21902 10560 22293 10588
rect 21902 10557 21914 10560
rect 21856 10551 21914 10557
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 25038 10548 25044 10600
rect 25096 10588 25102 10600
rect 25752 10591 25810 10597
rect 25752 10588 25764 10591
rect 25096 10560 25764 10588
rect 25096 10548 25102 10560
rect 25752 10557 25764 10560
rect 25798 10588 25810 10591
rect 26234 10588 26240 10600
rect 25798 10560 26240 10588
rect 25798 10557 25810 10560
rect 25752 10551 25810 10557
rect 26234 10548 26240 10560
rect 26292 10548 26298 10600
rect 26602 10548 26608 10600
rect 26660 10588 26666 10600
rect 26732 10591 26790 10597
rect 26732 10588 26744 10591
rect 26660 10560 26744 10588
rect 26660 10548 26666 10560
rect 26732 10557 26744 10560
rect 26778 10588 26790 10591
rect 27157 10591 27215 10597
rect 27157 10588 27169 10591
rect 26778 10560 27169 10588
rect 26778 10557 26790 10560
rect 26732 10551 26790 10557
rect 27157 10557 27169 10560
rect 27203 10557 27215 10591
rect 27157 10551 27215 10557
rect 27776 10591 27834 10597
rect 27776 10557 27788 10591
rect 27822 10588 27834 10591
rect 27982 10588 27988 10600
rect 27822 10560 27988 10588
rect 27822 10557 27834 10560
rect 27776 10551 27834 10557
rect 27982 10548 27988 10560
rect 28040 10588 28046 10600
rect 28169 10591 28227 10597
rect 28169 10588 28181 10591
rect 28040 10560 28181 10588
rect 28040 10548 28046 10560
rect 28169 10557 28181 10560
rect 28215 10557 28227 10591
rect 28169 10551 28227 10557
rect 33296 10591 33354 10597
rect 33296 10557 33308 10591
rect 33342 10588 33354 10591
rect 35360 10588 35388 10616
rect 35437 10591 35495 10597
rect 35437 10588 35449 10591
rect 33342 10560 33732 10588
rect 35360 10560 35449 10588
rect 33342 10557 33354 10560
rect 33296 10551 33354 10557
rect 19199 10483 19257 10489
rect 19536 10492 20979 10520
rect 21085 10523 21143 10529
rect 19536 10464 19564 10492
rect 21085 10489 21097 10523
rect 21131 10520 21143 10523
rect 21361 10523 21419 10529
rect 21361 10520 21373 10523
rect 21131 10492 21373 10520
rect 21131 10489 21143 10492
rect 21085 10483 21143 10489
rect 21361 10489 21373 10492
rect 21407 10520 21419 10523
rect 23014 10520 23020 10532
rect 21407 10492 23020 10520
rect 21407 10489 21419 10492
rect 21361 10483 21419 10489
rect 23014 10480 23020 10492
rect 23072 10480 23078 10532
rect 26835 10523 26893 10529
rect 26835 10489 26847 10523
rect 26881 10520 26893 10523
rect 28626 10520 28632 10532
rect 26881 10492 28632 10520
rect 26881 10489 26893 10492
rect 26835 10483 26893 10489
rect 28626 10480 28632 10492
rect 28684 10480 28690 10532
rect 33704 10464 33732 10560
rect 35437 10557 35449 10560
rect 35483 10588 35495 10591
rect 35989 10591 36047 10597
rect 35989 10588 36001 10591
rect 35483 10560 36001 10588
rect 35483 10557 35495 10560
rect 35437 10551 35495 10557
rect 35989 10557 36001 10560
rect 36035 10557 36047 10591
rect 35989 10551 36047 10557
rect 12710 10452 12716 10464
rect 12207 10424 12480 10452
rect 12671 10424 12716 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 16724 10424 16865 10452
rect 16724 10412 16730 10424
rect 16853 10421 16865 10424
rect 16899 10421 16911 10455
rect 16853 10415 16911 10421
rect 17126 10412 17132 10464
rect 17184 10452 17190 10464
rect 18187 10455 18245 10461
rect 18187 10452 18199 10455
rect 17184 10424 18199 10452
rect 17184 10412 17190 10424
rect 18187 10421 18199 10424
rect 18233 10421 18245 10455
rect 19518 10452 19524 10464
rect 19479 10424 19524 10452
rect 18187 10415 18245 10421
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 20070 10412 20076 10464
rect 20128 10452 20134 10464
rect 20947 10455 21005 10461
rect 20947 10452 20959 10455
rect 20128 10424 20959 10452
rect 20128 10412 20134 10424
rect 20947 10421 20959 10424
rect 20993 10421 21005 10455
rect 20947 10415 21005 10421
rect 21959 10455 22017 10461
rect 21959 10421 21971 10455
rect 22005 10452 22017 10455
rect 22094 10452 22100 10464
rect 22005 10424 22100 10452
rect 22005 10421 22017 10424
rect 21959 10415 22017 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 25823 10455 25881 10461
rect 25823 10421 25835 10455
rect 25869 10452 25881 10455
rect 25958 10452 25964 10464
rect 25869 10424 25964 10452
rect 25869 10421 25881 10424
rect 25823 10415 25881 10421
rect 25958 10412 25964 10424
rect 26016 10412 26022 10464
rect 26605 10455 26663 10461
rect 26605 10421 26617 10455
rect 26651 10452 26663 10455
rect 26970 10452 26976 10464
rect 26651 10424 26976 10452
rect 26651 10421 26663 10424
rect 26605 10415 26663 10421
rect 26970 10412 26976 10424
rect 27028 10412 27034 10464
rect 27246 10412 27252 10464
rect 27304 10452 27310 10464
rect 27847 10455 27905 10461
rect 27847 10452 27859 10455
rect 27304 10424 27859 10452
rect 27304 10412 27310 10424
rect 27847 10421 27859 10424
rect 27893 10421 27905 10455
rect 27847 10415 27905 10421
rect 33042 10412 33048 10464
rect 33100 10452 33106 10464
rect 33367 10455 33425 10461
rect 33367 10452 33379 10455
rect 33100 10424 33379 10452
rect 33100 10412 33106 10424
rect 33367 10421 33379 10424
rect 33413 10421 33425 10455
rect 33686 10452 33692 10464
rect 33647 10424 33692 10452
rect 33367 10415 33425 10421
rect 33686 10412 33692 10424
rect 33744 10412 33750 10464
rect 34425 10455 34483 10461
rect 34425 10421 34437 10455
rect 34471 10452 34483 10455
rect 34606 10452 34612 10464
rect 34471 10424 34612 10452
rect 34471 10421 34483 10424
rect 34425 10415 34483 10421
rect 34606 10412 34612 10424
rect 34664 10452 34670 10464
rect 35158 10452 35164 10464
rect 34664 10424 35164 10452
rect 34664 10412 34670 10424
rect 35158 10412 35164 10424
rect 35216 10412 35222 10464
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 3510 10248 3516 10260
rect 3471 10220 3516 10248
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 4157 10251 4215 10257
rect 4157 10217 4169 10251
rect 4203 10217 4215 10251
rect 6730 10248 6736 10260
rect 6691 10220 6736 10248
rect 4157 10211 4215 10217
rect 3142 10140 3148 10192
rect 3200 10180 3206 10192
rect 4172 10180 4200 10211
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 13262 10248 13268 10260
rect 6972 10220 13268 10248
rect 6972 10208 6978 10220
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13446 10248 13452 10260
rect 13407 10220 13452 10248
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 14090 10248 14096 10260
rect 14051 10220 14096 10248
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 27157 10251 27215 10257
rect 27157 10217 27169 10251
rect 27203 10248 27215 10251
rect 27246 10248 27252 10260
rect 27203 10220 27252 10248
rect 27203 10217 27215 10220
rect 27157 10211 27215 10217
rect 27246 10208 27252 10220
rect 27304 10208 27310 10260
rect 35434 10248 35440 10260
rect 33923 10220 35440 10248
rect 4430 10180 4436 10192
rect 3200 10152 4200 10180
rect 4343 10152 4436 10180
rect 3200 10140 3206 10152
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1762 10072 1768 10124
rect 1820 10112 1826 10124
rect 1857 10115 1915 10121
rect 1857 10112 1869 10115
rect 1820 10084 1869 10112
rect 1820 10072 1826 10084
rect 1857 10081 1869 10084
rect 1903 10112 1915 10115
rect 2406 10112 2412 10124
rect 1903 10084 2412 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 4356 10121 4384 10152
rect 4430 10140 4436 10152
rect 4488 10180 4494 10192
rect 6822 10180 6828 10192
rect 4488 10152 6828 10180
rect 4488 10140 4494 10152
rect 6822 10140 6828 10152
rect 6880 10180 6886 10192
rect 10594 10180 10600 10192
rect 6880 10152 10600 10180
rect 6880 10140 6886 10152
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 12986 10180 12992 10192
rect 12728 10152 12992 10180
rect 2996 10115 3054 10121
rect 2996 10112 3008 10115
rect 2740 10084 3008 10112
rect 2740 10072 2746 10084
rect 2996 10081 3008 10084
rect 3042 10081 3054 10115
rect 2996 10075 3054 10081
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10081 4399 10115
rect 4341 10075 4399 10081
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 5696 10115 5754 10121
rect 5696 10081 5708 10115
rect 5742 10112 5754 10115
rect 5994 10112 6000 10124
rect 5742 10084 6000 10112
rect 5742 10081 5754 10084
rect 5696 10075 5754 10081
rect 1946 10044 1952 10056
rect 1907 10016 1952 10044
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 2314 10004 2320 10056
rect 2372 10044 2378 10056
rect 2501 10047 2559 10053
rect 2501 10044 2513 10047
rect 2372 10016 2513 10044
rect 2372 10004 2378 10016
rect 2501 10013 2513 10016
rect 2547 10044 2559 10047
rect 3878 10044 3884 10056
rect 2547 10016 3884 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 3878 10004 3884 10016
rect 3936 10044 3942 10056
rect 4540 10044 4568 10075
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 6914 10112 6920 10124
rect 6875 10084 6920 10112
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 8640 10115 8698 10121
rect 8640 10081 8652 10115
rect 8686 10112 8698 10115
rect 9398 10112 9404 10124
rect 8686 10084 9404 10112
rect 8686 10081 8698 10084
rect 8640 10075 8698 10081
rect 6546 10044 6552 10056
rect 3936 10016 6552 10044
rect 3936 10004 3942 10016
rect 6546 10004 6552 10016
rect 6604 10044 6610 10056
rect 7116 10044 7144 10075
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10284 10084 10517 10112
rect 10284 10072 10290 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10112 11023 10115
rect 11606 10112 11612 10124
rect 11011 10084 11612 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 11054 10044 11060 10056
rect 6604 10016 7144 10044
rect 11015 10016 11060 10044
rect 6604 10004 6610 10016
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 8711 9979 8769 9985
rect 8711 9945 8723 9979
rect 8757 9976 8769 9979
rect 12618 9976 12624 9988
rect 8757 9948 12624 9976
rect 8757 9945 8769 9948
rect 8711 9939 8769 9945
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 2777 9911 2835 9917
rect 2777 9908 2789 9911
rect 2556 9880 2789 9908
rect 2556 9868 2562 9880
rect 2777 9877 2789 9880
rect 2823 9877 2835 9911
rect 2777 9871 2835 9877
rect 3099 9911 3157 9917
rect 3099 9877 3111 9911
rect 3145 9908 3157 9911
rect 3234 9908 3240 9920
rect 3145 9880 3240 9908
rect 3145 9877 3157 9880
rect 3099 9871 3157 9877
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 5767 9911 5825 9917
rect 5767 9908 5779 9911
rect 4672 9880 5779 9908
rect 4672 9868 4678 9880
rect 5767 9877 5779 9880
rect 5813 9877 5825 9911
rect 11698 9908 11704 9920
rect 11659 9880 11704 9908
rect 5767 9871 5825 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 12526 9908 12532 9920
rect 12487 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 12728 9908 12756 10152
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 27430 10180 27436 10192
rect 27391 10152 27436 10180
rect 27430 10140 27436 10152
rect 27488 10140 27494 10192
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 13262 10112 13268 10124
rect 12851 10084 13268 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 16482 10121 16488 10124
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10112 16175 10115
rect 16439 10115 16488 10121
rect 16163 10084 16252 10112
rect 16163 10081 16175 10084
rect 16117 10075 16175 10081
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12912 10016 13185 10044
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 12912 9976 12940 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 12860 9948 12940 9976
rect 12970 9979 13028 9985
rect 12860 9936 12866 9948
rect 12970 9945 12982 9979
rect 13016 9976 13028 9979
rect 13016 9948 13216 9976
rect 13016 9945 13028 9948
rect 12970 9939 13028 9945
rect 13188 9920 13216 9948
rect 15470 9936 15476 9988
rect 15528 9976 15534 9988
rect 16224 9976 16252 10084
rect 16439 10081 16451 10115
rect 16485 10081 16488 10115
rect 16439 10075 16488 10081
rect 16482 10072 16488 10075
rect 16540 10112 16546 10124
rect 17770 10112 17776 10124
rect 16540 10084 16712 10112
rect 17731 10084 17776 10112
rect 16540 10072 16546 10084
rect 16298 10004 16304 10056
rect 16356 10044 16362 10056
rect 16684 10044 16712 10084
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 18233 10115 18291 10121
rect 18233 10112 18245 10115
rect 17920 10084 18245 10112
rect 17920 10072 17926 10084
rect 18233 10081 18245 10084
rect 18279 10081 18291 10115
rect 19334 10112 19340 10124
rect 19295 10084 19340 10112
rect 18233 10075 18291 10081
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20936 10115 20994 10121
rect 20936 10112 20948 10115
rect 20864 10084 20948 10112
rect 20864 10072 20870 10084
rect 20936 10081 20948 10084
rect 20982 10081 20994 10115
rect 20936 10075 20994 10081
rect 21980 10115 22038 10121
rect 21980 10081 21992 10115
rect 22026 10112 22038 10115
rect 22370 10112 22376 10124
rect 22026 10084 22376 10112
rect 22026 10081 22038 10084
rect 21980 10075 22038 10081
rect 22370 10072 22376 10084
rect 22428 10072 22434 10124
rect 22922 10112 22928 10124
rect 22883 10084 22928 10112
rect 22922 10072 22928 10084
rect 22980 10072 22986 10124
rect 24394 10112 24400 10124
rect 24355 10084 24400 10112
rect 24394 10072 24400 10084
rect 24452 10072 24458 10124
rect 25409 10115 25467 10121
rect 25409 10081 25421 10115
rect 25455 10112 25467 10115
rect 25498 10112 25504 10124
rect 25455 10084 25504 10112
rect 25455 10081 25467 10084
rect 25409 10075 25467 10081
rect 25498 10072 25504 10084
rect 25556 10072 25562 10124
rect 28718 10072 28724 10124
rect 28776 10112 28782 10124
rect 33502 10121 33508 10124
rect 28848 10115 28906 10121
rect 28848 10112 28860 10115
rect 28776 10084 28860 10112
rect 28776 10072 28782 10084
rect 28848 10081 28860 10084
rect 28894 10081 28906 10115
rect 33480 10115 33508 10121
rect 33480 10112 33492 10115
rect 33415 10084 33492 10112
rect 28848 10075 28906 10081
rect 33480 10081 33492 10084
rect 33560 10112 33566 10124
rect 33923 10112 33951 10220
rect 35434 10208 35440 10220
rect 35492 10208 35498 10260
rect 35621 10251 35679 10257
rect 35621 10217 35633 10251
rect 35667 10248 35679 10251
rect 35710 10248 35716 10260
rect 35667 10220 35716 10248
rect 35667 10217 35679 10220
rect 35621 10211 35679 10217
rect 35710 10208 35716 10220
rect 35768 10208 35774 10260
rect 33560 10084 33951 10112
rect 34476 10115 34534 10121
rect 33480 10075 33508 10081
rect 33502 10072 33508 10075
rect 33560 10072 33566 10084
rect 34476 10081 34488 10115
rect 34522 10112 34534 10115
rect 34698 10112 34704 10124
rect 34522 10084 34704 10112
rect 34522 10081 34534 10084
rect 34476 10075 34534 10081
rect 34698 10072 34704 10084
rect 34756 10072 34762 10124
rect 35437 10115 35495 10121
rect 35437 10081 35449 10115
rect 35483 10112 35495 10115
rect 35894 10112 35900 10124
rect 35483 10084 35900 10112
rect 35483 10081 35495 10084
rect 35437 10075 35495 10081
rect 35894 10072 35900 10084
rect 35952 10072 35958 10124
rect 36078 10072 36084 10124
rect 36136 10112 36142 10124
rect 36576 10115 36634 10121
rect 36576 10112 36588 10115
rect 36136 10084 36588 10112
rect 36136 10072 36142 10084
rect 36556 10081 36588 10084
rect 36622 10081 36634 10115
rect 36556 10075 36634 10081
rect 17880 10044 17908 10072
rect 18506 10044 18512 10056
rect 16356 10016 16401 10044
rect 16684 10016 17908 10044
rect 18467 10016 18512 10044
rect 16356 10004 16362 10016
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 21453 10047 21511 10053
rect 21453 10013 21465 10047
rect 21499 10044 21511 10047
rect 21542 10044 21548 10056
rect 21499 10016 21548 10044
rect 21499 10013 21511 10016
rect 21453 10007 21511 10013
rect 21542 10004 21548 10016
rect 21600 10004 21606 10056
rect 27154 10004 27160 10056
rect 27212 10044 27218 10056
rect 27341 10047 27399 10053
rect 27341 10044 27353 10047
rect 27212 10016 27353 10044
rect 27212 10004 27218 10016
rect 27341 10013 27353 10016
rect 27387 10013 27399 10047
rect 27341 10007 27399 10013
rect 27985 10047 28043 10053
rect 27985 10013 27997 10047
rect 28031 10044 28043 10047
rect 29178 10044 29184 10056
rect 28031 10016 29184 10044
rect 28031 10013 28043 10016
rect 27985 10007 28043 10013
rect 29178 10004 29184 10016
rect 29236 10004 29242 10056
rect 34563 10047 34621 10053
rect 34563 10013 34575 10047
rect 34609 10044 34621 10047
rect 36556 10044 36584 10075
rect 37458 10044 37464 10056
rect 34609 10016 35525 10044
rect 36556 10016 37464 10044
rect 34609 10013 34621 10016
rect 34563 10007 34621 10013
rect 18230 9976 18236 9988
rect 15528 9948 18236 9976
rect 15528 9936 15534 9948
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 27062 9936 27068 9988
rect 27120 9976 27126 9988
rect 28951 9979 29009 9985
rect 28951 9976 28963 9979
rect 27120 9948 28963 9976
rect 27120 9936 27126 9948
rect 28951 9945 28963 9948
rect 28997 9945 29009 9979
rect 28951 9939 29009 9945
rect 33551 9979 33609 9985
rect 33551 9945 33563 9979
rect 33597 9976 33609 9979
rect 35342 9976 35348 9988
rect 33597 9948 35348 9976
rect 33597 9945 33609 9948
rect 33551 9939 33609 9945
rect 35342 9936 35348 9948
rect 35400 9936 35406 9988
rect 35497 9976 35525 10016
rect 37458 10004 37464 10016
rect 37516 10004 37522 10056
rect 36538 9976 36544 9988
rect 35497 9948 36544 9976
rect 36538 9936 36544 9948
rect 36596 9936 36602 9988
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 12728 9880 13093 9908
rect 13081 9877 13093 9880
rect 13127 9877 13139 9911
rect 13081 9871 13139 9877
rect 13170 9868 13176 9920
rect 13228 9868 13234 9920
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 14553 9911 14611 9917
rect 14553 9908 14565 9911
rect 14240 9880 14565 9908
rect 14240 9868 14246 9880
rect 14553 9877 14565 9880
rect 14599 9908 14611 9911
rect 15286 9908 15292 9920
rect 14599 9880 15292 9908
rect 14599 9877 14611 9880
rect 14553 9871 14611 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 19475 9911 19533 9917
rect 19475 9877 19487 9911
rect 19521 9908 19533 9911
rect 19702 9908 19708 9920
rect 19521 9880 19708 9908
rect 19521 9877 19533 9880
rect 19475 9871 19533 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 20162 9908 20168 9920
rect 19935 9880 20168 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 21039 9911 21097 9917
rect 21039 9877 21051 9911
rect 21085 9908 21097 9911
rect 21266 9908 21272 9920
rect 21085 9880 21272 9908
rect 21085 9877 21097 9880
rect 21039 9871 21097 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 21729 9911 21787 9917
rect 21729 9908 21741 9911
rect 21508 9880 21741 9908
rect 21508 9868 21514 9880
rect 21729 9877 21741 9880
rect 21775 9877 21787 9911
rect 21729 9871 21787 9877
rect 21818 9868 21824 9920
rect 21876 9908 21882 9920
rect 22051 9911 22109 9917
rect 22051 9908 22063 9911
rect 21876 9880 22063 9908
rect 21876 9868 21882 9880
rect 22051 9877 22063 9880
rect 22097 9877 22109 9911
rect 22051 9871 22109 9877
rect 23109 9911 23167 9917
rect 23109 9877 23121 9911
rect 23155 9908 23167 9911
rect 23382 9908 23388 9920
rect 23155 9880 23388 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 23382 9868 23388 9880
rect 23440 9908 23446 9920
rect 24121 9911 24179 9917
rect 24121 9908 24133 9911
rect 23440 9880 24133 9908
rect 23440 9868 23446 9880
rect 24121 9877 24133 9880
rect 24167 9877 24179 9911
rect 24121 9871 24179 9877
rect 24581 9911 24639 9917
rect 24581 9877 24593 9911
rect 24627 9908 24639 9911
rect 24762 9908 24768 9920
rect 24627 9880 24768 9908
rect 24627 9877 24639 9880
rect 24581 9871 24639 9877
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 25547 9911 25605 9917
rect 25547 9877 25559 9911
rect 25593 9908 25605 9911
rect 28166 9908 28172 9920
rect 25593 9880 28172 9908
rect 25593 9877 25605 9880
rect 25547 9871 25605 9877
rect 28166 9868 28172 9880
rect 28224 9868 28230 9920
rect 35434 9868 35440 9920
rect 35492 9908 35498 9920
rect 36679 9911 36737 9917
rect 36679 9908 36691 9911
rect 35492 9880 36691 9908
rect 35492 9868 35498 9880
rect 36679 9877 36691 9880
rect 36725 9877 36737 9911
rect 36679 9871 36737 9877
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 4065 9707 4123 9713
rect 4065 9704 4077 9707
rect 3936 9676 4077 9704
rect 3936 9664 3942 9676
rect 4065 9673 4077 9676
rect 4111 9673 4123 9707
rect 6546 9704 6552 9716
rect 6507 9676 6552 9704
rect 4065 9667 4123 9673
rect 6546 9664 6552 9676
rect 6604 9704 6610 9716
rect 8202 9704 8208 9716
rect 6604 9676 8208 9704
rect 6604 9664 6610 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 10226 9704 10232 9716
rect 10187 9676 10232 9704
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 11517 9707 11575 9713
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11606 9704 11612 9716
rect 11563 9676 11612 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 3970 9596 3976 9648
rect 4028 9636 4034 9648
rect 5994 9636 6000 9648
rect 4028 9608 6000 9636
rect 4028 9596 4034 9608
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 6273 9639 6331 9645
rect 6273 9605 6285 9639
rect 6319 9636 6331 9639
rect 6914 9636 6920 9648
rect 6319 9608 6920 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 3510 9568 3516 9580
rect 3099 9540 3516 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 3878 9568 3884 9580
rect 3752 9540 3884 9568
rect 3752 9528 3758 9540
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 5684 9540 7205 9568
rect 5684 9528 5690 9540
rect 7193 9537 7205 9540
rect 7239 9568 7251 9571
rect 7558 9568 7564 9580
rect 7239 9540 7564 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8220 9568 8248 9664
rect 8662 9568 8668 9580
rect 8220 9540 8668 9568
rect 8662 9528 8668 9540
rect 8720 9568 8726 9580
rect 9953 9571 10011 9577
rect 8720 9540 8892 9568
rect 8720 9528 8726 9540
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 1670 9500 1676 9512
rect 1627 9472 1676 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2406 9500 2412 9512
rect 1995 9472 2412 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 2498 9460 2504 9512
rect 2556 9500 2562 9512
rect 2556 9472 2912 9500
rect 2556 9460 2562 9472
rect 2130 9432 2136 9444
rect 2091 9404 2136 9432
rect 2130 9392 2136 9404
rect 2188 9392 2194 9444
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 2777 9367 2835 9373
rect 2777 9364 2789 9367
rect 2740 9336 2789 9364
rect 2740 9324 2746 9336
rect 2777 9333 2789 9336
rect 2823 9333 2835 9367
rect 2884 9364 2912 9472
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 4154 9500 4160 9512
rect 3844 9472 4160 9500
rect 3844 9460 3850 9472
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 5074 9500 5080 9512
rect 4479 9472 5080 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5902 9500 5908 9512
rect 5307 9472 5908 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8864 9509 8892 9540
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 9999 9540 10732 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10704 9512 10732 9540
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 8849 9463 8907 9469
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10744 9472 10977 9500
rect 10744 9460 10750 9472
rect 10965 9469 10977 9472
rect 11011 9500 11023 9503
rect 11532 9500 11560 9667
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11790 9704 11796 9716
rect 11751 9676 11796 9704
rect 11790 9664 11796 9676
rect 11848 9704 11854 9716
rect 15470 9704 15476 9716
rect 11848 9676 12572 9704
rect 15431 9676 15476 9704
rect 11848 9664 11854 9676
rect 12544 9577 12572 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 15841 9707 15899 9713
rect 15841 9673 15853 9707
rect 15887 9704 15899 9707
rect 16482 9704 16488 9716
rect 15887 9676 16488 9704
rect 15887 9673 15899 9676
rect 15841 9667 15899 9673
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 17494 9704 17500 9716
rect 17407 9676 17500 9704
rect 17494 9664 17500 9676
rect 17552 9704 17558 9716
rect 17770 9704 17776 9716
rect 17552 9676 17776 9704
rect 17552 9664 17558 9676
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 19334 9704 19340 9716
rect 19295 9676 19340 9704
rect 19334 9664 19340 9676
rect 19392 9704 19398 9716
rect 20806 9704 20812 9716
rect 19392 9676 20812 9704
rect 19392 9664 19398 9676
rect 20806 9664 20812 9676
rect 20864 9704 20870 9716
rect 20901 9707 20959 9713
rect 20901 9704 20913 9707
rect 20864 9676 20913 9704
rect 20864 9664 20870 9676
rect 20901 9673 20913 9676
rect 20947 9704 20959 9707
rect 21634 9704 21640 9716
rect 20947 9676 21640 9704
rect 20947 9673 20959 9676
rect 20901 9667 20959 9673
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 22370 9704 22376 9716
rect 22331 9676 22376 9704
rect 22370 9664 22376 9676
rect 22428 9674 22434 9716
rect 22428 9664 22508 9674
rect 26602 9664 26608 9716
rect 26660 9704 26666 9716
rect 32214 9704 32220 9716
rect 26660 9676 32220 9704
rect 26660 9664 26666 9676
rect 13170 9596 13176 9648
rect 13228 9636 13234 9648
rect 22388 9646 22508 9664
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 13228 9608 13461 9636
rect 13228 9596 13234 9608
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 22480 9636 22508 9646
rect 25498 9636 25504 9648
rect 13449 9599 13507 9605
rect 18426 9608 22324 9636
rect 22480 9608 24256 9636
rect 25459 9608 25504 9636
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 13722 9568 13728 9580
rect 12768 9540 13728 9568
rect 12768 9528 12774 9540
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15712 9540 16037 9568
rect 15712 9528 15718 9540
rect 16025 9537 16037 9540
rect 16071 9568 16083 9571
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 16071 9540 16957 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 16945 9537 16957 9540
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 11011 9472 11560 9500
rect 13173 9503 13231 9509
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 13173 9469 13185 9503
rect 13219 9500 13231 9503
rect 13538 9500 13544 9512
rect 13219 9472 13544 9500
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 3145 9435 3203 9441
rect 3145 9401 3157 9435
rect 3191 9432 3203 9435
rect 3418 9432 3424 9444
rect 3191 9404 3424 9432
rect 3191 9401 3203 9404
rect 3145 9395 3203 9401
rect 3418 9392 3424 9404
rect 3476 9392 3482 9444
rect 3694 9432 3700 9444
rect 3607 9404 3700 9432
rect 3694 9392 3700 9404
rect 3752 9432 3758 9444
rect 6917 9435 6975 9441
rect 6917 9432 6929 9435
rect 3752 9404 6929 9432
rect 3752 9392 3758 9404
rect 6917 9401 6929 9404
rect 6963 9401 6975 9435
rect 6917 9395 6975 9401
rect 3970 9364 3976 9376
rect 2884 9336 3976 9364
rect 2777 9327 2835 9333
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 5721 9367 5779 9373
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 5994 9364 6000 9376
rect 5767 9336 6000 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6932 9364 6960 9395
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7064 9404 7109 9432
rect 7064 9392 7070 9404
rect 12526 9392 12532 9444
rect 12584 9432 12590 9444
rect 12621 9435 12679 9441
rect 12621 9432 12633 9435
rect 12584 9404 12633 9432
rect 12584 9392 12590 9404
rect 12621 9401 12633 9404
rect 12667 9401 12679 9435
rect 12621 9395 12679 9401
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 13814 9432 13820 9444
rect 13320 9404 13820 9432
rect 13320 9392 13326 9404
rect 13814 9392 13820 9404
rect 13872 9432 13878 9444
rect 14277 9435 14335 9441
rect 13872 9404 13965 9432
rect 13872 9392 13878 9404
rect 14277 9401 14289 9435
rect 14323 9432 14335 9435
rect 15028 9432 15056 9463
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 18288 9472 18337 9500
rect 18288 9460 18294 9472
rect 18325 9469 18337 9472
rect 18371 9500 18383 9503
rect 18426 9500 18454 9608
rect 20530 9528 20536 9580
rect 20588 9568 20594 9580
rect 21729 9571 21787 9577
rect 21729 9568 21741 9571
rect 20588 9540 21741 9568
rect 20588 9528 20594 9540
rect 21729 9537 21741 9540
rect 21775 9537 21787 9571
rect 22296 9568 22324 9608
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 22296 9540 23949 9568
rect 21729 9531 21787 9537
rect 23937 9537 23949 9540
rect 23983 9568 23995 9571
rect 24228 9568 24256 9608
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 27338 9596 27344 9648
rect 27396 9636 27402 9648
rect 29411 9639 29469 9645
rect 29411 9636 29423 9639
rect 27396 9608 29423 9636
rect 27396 9596 27402 9608
rect 29411 9605 29423 9608
rect 29457 9605 29469 9639
rect 29411 9599 29469 9605
rect 23983 9540 24164 9568
rect 24228 9540 26439 9568
rect 23983 9537 23995 9540
rect 23937 9531 23995 9537
rect 24136 9512 24164 9540
rect 18371 9472 18454 9500
rect 18601 9503 18659 9509
rect 18371 9469 18383 9472
rect 18325 9463 18383 9469
rect 18601 9469 18613 9503
rect 18647 9500 18659 9503
rect 18874 9500 18880 9512
rect 18647 9472 18880 9500
rect 18647 9469 18659 9472
rect 18601 9463 18659 9469
rect 18874 9460 18880 9472
rect 18932 9460 18938 9512
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 19978 9500 19984 9512
rect 19935 9472 19984 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 20162 9500 20168 9512
rect 20123 9472 20168 9500
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 24118 9500 24124 9512
rect 24031 9472 24124 9500
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 26411 9509 26439 9540
rect 27246 9528 27252 9580
rect 27304 9568 27310 9580
rect 27433 9571 27491 9577
rect 27433 9568 27445 9571
rect 27304 9540 27445 9568
rect 27304 9528 27310 9540
rect 27433 9537 27445 9540
rect 27479 9537 27491 9571
rect 27433 9531 27491 9537
rect 24581 9503 24639 9509
rect 24581 9469 24593 9503
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 26396 9503 26454 9509
rect 26396 9469 26408 9503
rect 26442 9500 26454 9503
rect 29340 9503 29398 9509
rect 26442 9472 26924 9500
rect 26442 9469 26454 9472
rect 26396 9463 26454 9469
rect 14323 9404 15700 9432
rect 14323 9401 14335 9404
rect 14277 9395 14335 9401
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 6932 9336 7849 9364
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 8352 9336 8493 9364
rect 8352 9324 8358 9336
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 9398 9364 9404 9376
rect 9359 9336 9404 9364
rect 8481 9327 8539 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 10502 9364 10508 9376
rect 10463 9336 10508 9364
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 12253 9367 12311 9373
rect 12253 9333 12265 9367
rect 12299 9364 12311 9367
rect 12710 9364 12716 9376
rect 12299 9336 12716 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 12710 9324 12716 9336
rect 12768 9364 12774 9376
rect 12986 9364 12992 9376
rect 12768 9336 12992 9364
rect 12768 9324 12774 9336
rect 12986 9324 12992 9336
rect 13044 9364 13050 9376
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 13044 9336 14657 9364
rect 13044 9324 13050 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 15672 9364 15700 9404
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 16666 9432 16672 9444
rect 16172 9404 16217 9432
rect 16627 9404 16672 9432
rect 16172 9392 16178 9404
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 21450 9432 21456 9444
rect 21411 9404 21456 9432
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 21542 9392 21548 9444
rect 21600 9432 21606 9444
rect 23658 9432 23664 9444
rect 21600 9404 21645 9432
rect 23446 9404 23664 9432
rect 21600 9392 21606 9404
rect 23446 9376 23474 9404
rect 23658 9392 23664 9404
rect 23716 9432 23722 9444
rect 24596 9432 24624 9463
rect 24854 9432 24860 9444
rect 23716 9404 24624 9432
rect 24815 9404 24860 9432
rect 23716 9392 23722 9404
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 26896 9376 26924 9472
rect 29340 9469 29352 9503
rect 29386 9500 29398 9503
rect 29822 9500 29828 9512
rect 29386 9472 29828 9500
rect 29386 9469 29398 9472
rect 29340 9463 29398 9469
rect 29822 9460 29828 9472
rect 29880 9460 29886 9512
rect 30282 9500 30288 9512
rect 30243 9472 30288 9500
rect 30282 9460 30288 9472
rect 30340 9500 30346 9512
rect 31839 9509 31867 9676
rect 32214 9664 32220 9676
rect 32272 9664 32278 9716
rect 33502 9704 33508 9716
rect 33463 9676 33508 9704
rect 33502 9664 33508 9676
rect 33560 9664 33566 9716
rect 35526 9704 35532 9716
rect 35487 9676 35532 9704
rect 35526 9664 35532 9676
rect 35584 9664 35590 9716
rect 35894 9704 35900 9716
rect 35855 9676 35900 9704
rect 35894 9664 35900 9676
rect 35952 9664 35958 9716
rect 36633 9707 36691 9713
rect 36633 9673 36645 9707
rect 36679 9704 36691 9707
rect 37642 9704 37648 9716
rect 36679 9676 37648 9704
rect 36679 9673 36691 9676
rect 36633 9667 36691 9673
rect 37642 9664 37648 9676
rect 37700 9664 37706 9716
rect 33594 9528 33600 9580
rect 33652 9568 33658 9580
rect 33689 9571 33747 9577
rect 33689 9568 33701 9571
rect 33652 9540 33701 9568
rect 33652 9528 33658 9540
rect 33689 9537 33701 9540
rect 33735 9568 33747 9571
rect 34333 9571 34391 9577
rect 34333 9568 34345 9571
rect 33735 9540 34345 9568
rect 33735 9537 33747 9540
rect 33689 9531 33747 9537
rect 34333 9537 34345 9540
rect 34379 9568 34391 9571
rect 35526 9568 35532 9580
rect 34379 9540 35532 9568
rect 34379 9537 34391 9540
rect 34333 9531 34391 9537
rect 35526 9528 35532 9540
rect 35584 9528 35590 9580
rect 30745 9503 30803 9509
rect 30745 9500 30757 9503
rect 30340 9472 30757 9500
rect 30340 9460 30346 9472
rect 30745 9469 30757 9472
rect 30791 9469 30803 9503
rect 30745 9463 30803 9469
rect 31808 9503 31867 9509
rect 31808 9469 31820 9503
rect 31854 9472 31867 9503
rect 32804 9503 32862 9509
rect 31854 9469 31866 9472
rect 31808 9463 31866 9469
rect 32804 9469 32816 9503
rect 32850 9469 32862 9503
rect 35345 9503 35403 9509
rect 35345 9500 35357 9503
rect 32804 9463 32862 9469
rect 35176 9472 35357 9500
rect 27249 9435 27307 9441
rect 27249 9401 27261 9435
rect 27295 9432 27307 9435
rect 27430 9432 27436 9444
rect 27295 9404 27436 9432
rect 27295 9401 27307 9404
rect 27249 9395 27307 9401
rect 27430 9392 27436 9404
rect 27488 9432 27494 9444
rect 27525 9435 27583 9441
rect 27525 9432 27537 9435
rect 27488 9404 27537 9432
rect 27488 9392 27494 9404
rect 27525 9401 27537 9404
rect 27571 9401 27583 9435
rect 28074 9432 28080 9444
rect 28035 9404 28080 9432
rect 27525 9395 27583 9401
rect 15930 9364 15936 9376
rect 15672 9336 15936 9364
rect 14645 9327 14703 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 17862 9364 17868 9376
rect 17823 9336 17868 9364
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18138 9364 18144 9376
rect 18099 9336 18144 9364
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 19886 9364 19892 9376
rect 19847 9336 19892 9364
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 22462 9324 22468 9376
rect 22520 9364 22526 9376
rect 22922 9364 22928 9376
rect 22520 9336 22928 9364
rect 22520 9324 22526 9336
rect 22922 9324 22928 9336
rect 22980 9324 22986 9376
rect 23382 9324 23388 9376
rect 23440 9336 23474 9376
rect 26467 9367 26525 9373
rect 23440 9324 23446 9336
rect 26467 9333 26479 9367
rect 26513 9364 26525 9367
rect 26694 9364 26700 9376
rect 26513 9336 26700 9364
rect 26513 9333 26525 9336
rect 26467 9327 26525 9333
rect 26694 9324 26700 9336
rect 26752 9324 26758 9376
rect 26878 9364 26884 9376
rect 26839 9336 26884 9364
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 27540 9364 27568 9395
rect 28074 9392 28080 9404
rect 28132 9392 28138 9444
rect 31895 9435 31953 9441
rect 31895 9401 31907 9435
rect 31941 9432 31953 9435
rect 32398 9432 32404 9444
rect 31941 9404 32404 9432
rect 31941 9401 31953 9404
rect 31895 9395 31953 9401
rect 32398 9392 32404 9404
rect 32456 9392 32462 9444
rect 32819 9432 32847 9463
rect 35176 9441 35204 9472
rect 35345 9469 35357 9472
rect 35391 9469 35403 9503
rect 36446 9500 36452 9512
rect 36407 9472 36452 9500
rect 35345 9463 35403 9469
rect 36446 9460 36452 9472
rect 36504 9500 36510 9512
rect 37001 9503 37059 9509
rect 37001 9500 37013 9503
rect 36504 9472 37013 9500
rect 36504 9460 36510 9472
rect 37001 9469 37013 9472
rect 37047 9469 37059 9503
rect 37001 9463 37059 9469
rect 35161 9435 35219 9441
rect 35161 9432 35173 9435
rect 32600 9404 35173 9432
rect 32600 9376 32628 9404
rect 35161 9401 35173 9404
rect 35207 9401 35219 9435
rect 35161 9395 35219 9401
rect 28353 9367 28411 9373
rect 28353 9364 28365 9367
rect 27540 9336 28365 9364
rect 28353 9333 28365 9336
rect 28399 9333 28411 9367
rect 28353 9327 28411 9333
rect 28718 9324 28724 9376
rect 28776 9364 28782 9376
rect 28813 9367 28871 9373
rect 28813 9364 28825 9367
rect 28776 9336 28825 9364
rect 28776 9324 28782 9336
rect 28813 9333 28825 9336
rect 28859 9333 28871 9367
rect 28813 9327 28871 9333
rect 30469 9367 30527 9373
rect 30469 9333 30481 9367
rect 30515 9364 30527 9367
rect 30650 9364 30656 9376
rect 30515 9336 30656 9364
rect 30515 9333 30527 9336
rect 30469 9327 30527 9333
rect 30650 9324 30656 9336
rect 30708 9324 30714 9376
rect 32582 9364 32588 9376
rect 32543 9336 32588 9364
rect 32582 9324 32588 9336
rect 32640 9324 32646 9376
rect 32907 9367 32965 9373
rect 32907 9333 32919 9367
rect 32953 9364 32965 9367
rect 33226 9364 33232 9376
rect 32953 9336 33232 9364
rect 32953 9333 32965 9336
rect 32907 9327 32965 9333
rect 33226 9324 33232 9336
rect 33284 9324 33290 9376
rect 33502 9324 33508 9376
rect 33560 9364 33566 9376
rect 33919 9367 33977 9373
rect 33919 9364 33931 9367
rect 33560 9336 33931 9364
rect 33560 9324 33566 9336
rect 33919 9333 33931 9336
rect 33965 9333 33977 9367
rect 34698 9364 34704 9376
rect 34659 9336 34704 9364
rect 33919 9327 33977 9333
rect 34698 9324 34704 9336
rect 34756 9324 34762 9376
rect 37458 9364 37464 9376
rect 37419 9336 37464 9364
rect 37458 9324 37464 9336
rect 37516 9324 37522 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1728 9132 1961 9160
rect 1728 9120 1734 9132
rect 1949 9129 1961 9132
rect 1995 9160 2007 9163
rect 2498 9160 2504 9172
rect 1995 9132 2504 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 3418 9160 3424 9172
rect 3379 9132 3424 9160
rect 3418 9120 3424 9132
rect 3476 9120 3482 9172
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 4890 9160 4896 9172
rect 3568 9132 4896 9160
rect 3568 9120 3574 9132
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 5592 9132 8201 9160
rect 5592 9120 5598 9132
rect 2314 9092 2320 9104
rect 2275 9064 2320 9092
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 2593 9095 2651 9101
rect 2593 9061 2605 9095
rect 2639 9092 2651 9095
rect 2866 9092 2872 9104
rect 2639 9064 2872 9092
rect 2639 9061 2651 9064
rect 2593 9055 2651 9061
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3694 9092 3700 9104
rect 3191 9064 3700 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3694 9052 3700 9064
rect 3752 9052 3758 9104
rect 4246 9092 4252 9104
rect 4207 9064 4252 9092
rect 4246 9052 4252 9064
rect 4304 9052 4310 9104
rect 7374 9092 7380 9104
rect 7335 9064 7380 9092
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 1464 9027 1522 9033
rect 1464 8993 1476 9027
rect 1510 9024 1522 9027
rect 1670 9024 1676 9036
rect 1510 8996 1676 9024
rect 1510 8993 1522 8996
rect 1464 8987 1522 8993
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 5718 9024 5724 9036
rect 5675 8996 5724 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 5902 9024 5908 9036
rect 5863 8996 5908 9024
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 8173 9024 8201 9132
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 10652 9132 11069 9160
rect 10652 9120 10658 9132
rect 11057 9129 11069 9132
rect 11103 9129 11115 9163
rect 11514 9160 11520 9172
rect 11475 9132 11520 9160
rect 11057 9123 11115 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 15654 9160 15660 9172
rect 15615 9132 15660 9160
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16209 9163 16267 9169
rect 16209 9160 16221 9163
rect 16172 9132 16221 9160
rect 16172 9120 16178 9132
rect 16209 9129 16221 9132
rect 16255 9160 16267 9163
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16255 9132 16497 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 16485 9123 16543 9129
rect 18141 9163 18199 9169
rect 18141 9129 18153 9163
rect 18187 9160 18199 9163
rect 18230 9160 18236 9172
rect 18187 9132 18236 9160
rect 18187 9129 18199 9132
rect 18141 9123 18199 9129
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 18690 9160 18696 9172
rect 18651 9132 18696 9160
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 20070 9160 20076 9172
rect 20031 9132 20076 9160
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 21450 9120 21456 9172
rect 21508 9160 21514 9172
rect 23891 9163 23949 9169
rect 23891 9160 23903 9163
rect 21508 9132 23903 9160
rect 21508 9120 21514 9132
rect 23891 9129 23903 9132
rect 23937 9129 23949 9163
rect 24394 9160 24400 9172
rect 24355 9132 24400 9160
rect 23891 9123 23949 9129
rect 24394 9120 24400 9132
rect 24452 9120 24458 9172
rect 26694 9120 26700 9172
rect 26752 9160 26758 9172
rect 28261 9163 28319 9169
rect 28261 9160 28273 9163
rect 26752 9132 28273 9160
rect 26752 9120 26758 9132
rect 27724 9104 27752 9132
rect 28261 9129 28273 9132
rect 28307 9129 28319 9163
rect 28626 9160 28632 9172
rect 28587 9132 28632 9160
rect 28261 9123 28319 9129
rect 28626 9120 28632 9132
rect 28684 9120 28690 9172
rect 33042 9120 33048 9172
rect 33100 9160 33106 9172
rect 33318 9160 33324 9172
rect 33100 9132 33324 9160
rect 33100 9120 33106 9132
rect 33318 9120 33324 9132
rect 33376 9120 33382 9172
rect 34698 9120 34704 9172
rect 34756 9160 34762 9172
rect 38654 9160 38660 9172
rect 34756 9132 38660 9160
rect 34756 9120 34762 9132
rect 38654 9120 38660 9132
rect 38712 9120 38718 9172
rect 11793 9095 11851 9101
rect 11793 9061 11805 9095
rect 11839 9092 11851 9095
rect 11882 9092 11888 9104
rect 11839 9064 11888 9092
rect 11839 9061 11851 9064
rect 11793 9055 11851 9061
rect 11882 9052 11888 9064
rect 11940 9092 11946 9104
rect 13357 9095 13415 9101
rect 13357 9092 13369 9095
rect 11940 9064 13369 9092
rect 11940 9052 11946 9064
rect 13357 9061 13369 9064
rect 13403 9092 13415 9095
rect 13446 9092 13452 9104
rect 13403 9064 13452 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 17221 9095 17279 9101
rect 17221 9061 17233 9095
rect 17267 9092 17279 9095
rect 17402 9092 17408 9104
rect 17267 9064 17408 9092
rect 17267 9061 17279 9064
rect 17221 9055 17279 9061
rect 17402 9052 17408 9064
rect 17460 9052 17466 9104
rect 18046 9052 18052 9104
rect 18104 9092 18110 9104
rect 18509 9095 18567 9101
rect 18509 9092 18521 9095
rect 18104 9064 18521 9092
rect 18104 9052 18110 9064
rect 18509 9061 18521 9064
rect 18555 9092 18567 9095
rect 18874 9092 18880 9104
rect 18555 9064 18880 9092
rect 18555 9061 18567 9064
rect 18509 9055 18567 9061
rect 18874 9052 18880 9064
rect 18932 9092 18938 9104
rect 21266 9092 21272 9104
rect 18932 9064 19196 9092
rect 21227 9064 21272 9092
rect 18932 9052 18938 9064
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 8173 8996 10057 9024
rect 10045 8993 10057 8996
rect 10091 9024 10103 9027
rect 10410 9024 10416 9036
rect 10091 8996 10416 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10686 9024 10692 9036
rect 10551 8996 10692 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 14826 8984 14832 9036
rect 14884 9024 14890 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14884 8996 15301 9024
rect 14884 8984 14890 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 19168 9033 19196 9064
rect 21266 9052 21272 9064
rect 21324 9052 21330 9104
rect 21358 9052 21364 9104
rect 21416 9092 21422 9104
rect 27338 9092 27344 9104
rect 21416 9064 21461 9092
rect 27299 9064 27344 9092
rect 21416 9052 21422 9064
rect 27338 9052 27344 9064
rect 27396 9052 27402 9104
rect 27433 9095 27491 9101
rect 27433 9061 27445 9095
rect 27479 9092 27491 9095
rect 27522 9092 27528 9104
rect 27479 9064 27528 9092
rect 27479 9061 27491 9064
rect 27433 9055 27491 9061
rect 27522 9052 27528 9064
rect 27580 9052 27586 9104
rect 27706 9052 27712 9104
rect 27764 9052 27770 9104
rect 28994 9092 29000 9104
rect 28955 9064 29000 9092
rect 28994 9052 29000 9064
rect 29052 9052 29058 9104
rect 34057 9095 34115 9101
rect 34057 9061 34069 9095
rect 34103 9092 34115 9095
rect 34146 9092 34152 9104
rect 34103 9064 34152 9092
rect 34103 9061 34115 9064
rect 34057 9055 34115 9061
rect 34146 9052 34152 9064
rect 34204 9052 34210 9104
rect 35618 9092 35624 9104
rect 35579 9064 35624 9092
rect 35618 9052 35624 9064
rect 35676 9052 35682 9104
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 17828 8996 18613 9024
rect 17828 8984 17834 8996
rect 18601 8993 18613 8996
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 9024 19211 9027
rect 20162 9024 20168 9036
rect 19199 8996 20168 9024
rect 19199 8993 19211 8996
rect 19153 8987 19211 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 3602 8956 3608 8968
rect 2547 8928 3608 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4798 8956 4804 8968
rect 4203 8928 4804 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 6086 8956 6092 8968
rect 5040 8928 5764 8956
rect 6047 8928 6092 8956
rect 5040 8916 5046 8928
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 4614 8888 4620 8900
rect 3108 8860 4620 8888
rect 3108 8848 3114 8860
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 5736 8897 5764 8928
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 7282 8956 7288 8968
rect 7243 8928 7288 8956
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 7558 8956 7564 8968
rect 7519 8928 7564 8956
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 10594 8956 10600 8968
rect 10555 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 11698 8956 11704 8968
rect 11659 8928 11704 8956
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 11974 8956 11980 8968
rect 11935 8928 11980 8956
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 13078 8916 13084 8968
rect 13136 8956 13142 8968
rect 13265 8959 13323 8965
rect 13265 8956 13277 8959
rect 13136 8928 13277 8956
rect 13136 8916 13142 8928
rect 13265 8925 13277 8928
rect 13311 8925 13323 8959
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13265 8919 13323 8925
rect 13538 8916 13544 8928
rect 13596 8956 13602 8968
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 13596 8928 13814 8956
rect 13596 8916 13602 8928
rect 4709 8891 4767 8897
rect 4709 8857 4721 8891
rect 4755 8888 4767 8891
rect 5721 8891 5779 8897
rect 4755 8860 5304 8888
rect 4755 8857 4767 8860
rect 4709 8851 4767 8857
rect 5276 8832 5304 8860
rect 5721 8857 5733 8891
rect 5767 8857 5779 8891
rect 5721 8851 5779 8857
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 8570 8888 8576 8900
rect 8527 8860 8576 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 8570 8848 8576 8860
rect 8628 8888 8634 8900
rect 9030 8888 9036 8900
rect 8628 8860 9036 8888
rect 8628 8848 8634 8860
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 11606 8848 11612 8900
rect 11664 8888 11670 8900
rect 13630 8888 13636 8900
rect 11664 8860 13636 8888
rect 11664 8848 11670 8860
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 13786 8888 13814 8928
rect 16868 8928 17141 8956
rect 16868 8897 16896 8928
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17405 8959 17463 8965
rect 17405 8925 17417 8959
rect 17451 8925 17463 8959
rect 18616 8956 18644 8987
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 22738 9024 22744 9036
rect 22699 8996 22744 9024
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 23820 9027 23878 9033
rect 23820 8993 23832 9027
rect 23866 9024 23878 9027
rect 23934 9024 23940 9036
rect 23866 8996 23940 9024
rect 23866 8993 23878 8996
rect 23820 8987 23878 8993
rect 23934 8984 23940 8996
rect 23992 8984 23998 9036
rect 24118 8984 24124 9036
rect 24176 9024 24182 9036
rect 24857 9027 24915 9033
rect 24857 9024 24869 9027
rect 24176 8996 24869 9024
rect 24176 8984 24182 8996
rect 24857 8993 24869 8996
rect 24903 9024 24915 9027
rect 25222 9024 25228 9036
rect 24903 8996 25228 9024
rect 24903 8993 24915 8996
rect 24857 8987 24915 8993
rect 25222 8984 25228 8996
rect 25280 8984 25286 9036
rect 25406 9024 25412 9036
rect 25367 8996 25412 9024
rect 25406 8984 25412 8996
rect 25464 8984 25470 9036
rect 30374 9024 30380 9036
rect 30335 8996 30380 9024
rect 30374 8984 30380 8996
rect 30432 8984 30438 9036
rect 32306 9024 32312 9036
rect 32267 8996 32312 9024
rect 32306 8984 32312 8996
rect 32364 8984 32370 9036
rect 32674 9024 32680 9036
rect 32635 8996 32680 9024
rect 32674 8984 32680 8996
rect 32732 8984 32738 9036
rect 19242 8956 19248 8968
rect 18616 8928 19248 8956
rect 17405 8919 17463 8925
rect 16853 8891 16911 8897
rect 16853 8888 16865 8891
rect 13786 8860 16865 8888
rect 16853 8857 16865 8860
rect 16899 8857 16911 8891
rect 16853 8851 16911 8857
rect 1535 8823 1593 8829
rect 1535 8789 1547 8823
rect 1581 8820 1593 8823
rect 1762 8820 1768 8832
rect 1581 8792 1768 8820
rect 1581 8789 1593 8792
rect 1535 8783 1593 8789
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 4430 8820 4436 8832
rect 3927 8792 4436 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 5258 8820 5264 8832
rect 5219 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 8849 8823 8907 8829
rect 8849 8820 8861 8823
rect 8812 8792 8861 8820
rect 8812 8780 8818 8792
rect 8849 8789 8861 8792
rect 8895 8789 8907 8823
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 8849 8783 8907 8789
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13648 8820 13676 8848
rect 16298 8820 16304 8832
rect 13648 8792 16304 8820
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17420 8820 17448 8919
rect 19242 8916 19248 8928
rect 19300 8956 19306 8968
rect 21726 8956 21732 8968
rect 19300 8928 21732 8956
rect 19300 8916 19306 8928
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 21913 8959 21971 8965
rect 21913 8925 21925 8959
rect 21959 8956 21971 8959
rect 22186 8956 22192 8968
rect 21959 8928 22192 8956
rect 21959 8925 21971 8928
rect 21913 8919 21971 8925
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 25590 8956 25596 8968
rect 25551 8928 25596 8956
rect 25590 8916 25596 8928
rect 25648 8916 25654 8968
rect 27985 8959 28043 8965
rect 27985 8925 27997 8959
rect 28031 8956 28043 8959
rect 28074 8956 28080 8968
rect 28031 8928 28080 8956
rect 28031 8925 28043 8928
rect 27985 8919 28043 8925
rect 28074 8916 28080 8928
rect 28132 8956 28138 8968
rect 28534 8956 28540 8968
rect 28132 8928 28540 8956
rect 28132 8916 28138 8928
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 28626 8916 28632 8968
rect 28684 8956 28690 8968
rect 28905 8959 28963 8965
rect 28905 8956 28917 8959
rect 28684 8928 28917 8956
rect 28684 8916 28690 8928
rect 28905 8925 28917 8928
rect 28951 8925 28963 8959
rect 29178 8956 29184 8968
rect 29139 8928 29184 8956
rect 28905 8919 28963 8925
rect 29178 8916 29184 8928
rect 29236 8916 29242 8968
rect 32858 8956 32864 8968
rect 32819 8928 32864 8956
rect 32858 8916 32864 8928
rect 32916 8916 32922 8968
rect 33226 8916 33232 8968
rect 33284 8956 33290 8968
rect 33962 8956 33968 8968
rect 33284 8928 33968 8956
rect 33284 8916 33290 8928
rect 33962 8916 33968 8928
rect 34020 8916 34026 8968
rect 34054 8916 34060 8968
rect 34112 8956 34118 8968
rect 34241 8959 34299 8965
rect 34241 8956 34253 8959
rect 34112 8928 34253 8956
rect 34112 8916 34118 8928
rect 34241 8925 34253 8928
rect 34287 8925 34299 8959
rect 34241 8919 34299 8925
rect 35342 8916 35348 8968
rect 35400 8956 35406 8968
rect 35529 8959 35587 8965
rect 35529 8956 35541 8959
rect 35400 8928 35541 8956
rect 35400 8916 35406 8928
rect 35529 8925 35541 8928
rect 35575 8956 35587 8959
rect 36262 8956 36268 8968
rect 35575 8928 36268 8956
rect 35575 8925 35587 8928
rect 35529 8919 35587 8925
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 19705 8891 19763 8897
rect 19705 8857 19717 8891
rect 19751 8888 19763 8891
rect 19978 8888 19984 8900
rect 19751 8860 19984 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 19978 8848 19984 8860
rect 20036 8888 20042 8900
rect 23382 8888 23388 8900
rect 20036 8860 23388 8888
rect 20036 8848 20042 8860
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 26694 8848 26700 8900
rect 26752 8888 26758 8900
rect 30515 8891 30573 8897
rect 30515 8888 30527 8891
rect 26752 8860 30527 8888
rect 26752 8848 26758 8860
rect 30515 8857 30527 8860
rect 30561 8857 30573 8891
rect 30515 8851 30573 8857
rect 36081 8891 36139 8897
rect 36081 8857 36093 8891
rect 36127 8888 36139 8891
rect 36814 8888 36820 8900
rect 36127 8860 36820 8888
rect 36127 8857 36139 8860
rect 36081 8851 36139 8857
rect 36814 8848 36820 8860
rect 36872 8848 36878 8900
rect 16724 8792 17448 8820
rect 16724 8780 16730 8792
rect 21450 8780 21456 8832
rect 21508 8820 21514 8832
rect 22281 8823 22339 8829
rect 22281 8820 22293 8823
rect 21508 8792 22293 8820
rect 21508 8780 21514 8792
rect 22281 8789 22293 8792
rect 22327 8820 22339 8823
rect 22879 8823 22937 8829
rect 22879 8820 22891 8823
rect 22327 8792 22891 8820
rect 22327 8789 22339 8792
rect 22281 8783 22339 8789
rect 22879 8789 22891 8792
rect 22925 8789 22937 8823
rect 22879 8783 22937 8789
rect 23106 8780 23112 8832
rect 23164 8820 23170 8832
rect 24394 8820 24400 8832
rect 23164 8792 24400 8820
rect 23164 8780 23170 8792
rect 24394 8780 24400 8792
rect 24452 8780 24458 8832
rect 27154 8820 27160 8832
rect 27115 8792 27160 8820
rect 27154 8780 27160 8792
rect 27212 8780 27218 8832
rect 31297 8823 31355 8829
rect 31297 8789 31309 8823
rect 31343 8820 31355 8823
rect 31386 8820 31392 8832
rect 31343 8792 31392 8820
rect 31343 8789 31355 8792
rect 31297 8783 31355 8789
rect 31386 8780 31392 8792
rect 31444 8780 31450 8832
rect 33134 8780 33140 8832
rect 33192 8820 33198 8832
rect 33229 8823 33287 8829
rect 33229 8820 33241 8823
rect 33192 8792 33241 8820
rect 33192 8780 33198 8792
rect 33229 8789 33241 8792
rect 33275 8789 33287 8823
rect 33229 8783 33287 8789
rect 33318 8780 33324 8832
rect 33376 8820 33382 8832
rect 33597 8823 33655 8829
rect 33597 8820 33609 8823
rect 33376 8792 33609 8820
rect 33376 8780 33382 8792
rect 33597 8789 33609 8792
rect 33643 8789 33655 8823
rect 34974 8820 34980 8832
rect 34935 8792 34980 8820
rect 33597 8783 33655 8789
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2406 8576 2412 8588
rect 2464 8616 2470 8628
rect 4157 8619 4215 8625
rect 2464 8588 3832 8616
rect 2464 8576 2470 8588
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 3694 8548 3700 8560
rect 3651 8520 3700 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 3694 8508 3700 8520
rect 3752 8508 3758 8560
rect 3804 8548 3832 8588
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4246 8616 4252 8628
rect 4203 8588 4252 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4798 8616 4804 8628
rect 4571 8588 4804 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 7374 8576 7380 8628
rect 7432 8616 7438 8628
rect 8018 8616 8024 8628
rect 7432 8588 8024 8616
rect 7432 8576 7438 8588
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8662 8616 8668 8628
rect 8623 8588 8668 8616
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10686 8616 10692 8628
rect 10183 8588 10692 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11514 8616 11520 8628
rect 11394 8588 11520 8616
rect 4430 8548 4436 8560
rect 3804 8520 4436 8548
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 7282 8508 7288 8560
rect 7340 8548 7346 8560
rect 8297 8551 8355 8557
rect 8297 8548 8309 8551
rect 7340 8520 8309 8548
rect 7340 8508 7346 8520
rect 8297 8517 8309 8520
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8480 1547 8483
rect 1578 8480 1584 8492
rect 1535 8452 1584 8480
rect 1535 8449 1547 8452
rect 1489 8443 1547 8449
rect 1578 8440 1584 8452
rect 1636 8480 1642 8492
rect 1854 8480 1860 8492
rect 1636 8452 1860 8480
rect 1636 8440 1642 8452
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 5258 8480 5264 8492
rect 2179 8452 5264 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5626 8480 5632 8492
rect 5587 8452 5632 8480
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 8680 8480 8708 8576
rect 10410 8548 10416 8560
rect 10371 8520 10416 8548
rect 10410 8508 10416 8520
rect 10468 8508 10474 8560
rect 10873 8483 10931 8489
rect 8680 8452 9352 8480
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7147 8384 8156 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 3050 8344 3056 8356
rect 1636 8316 1681 8344
rect 3011 8316 3056 8344
rect 1636 8304 1642 8316
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8313 3203 8347
rect 5350 8344 5356 8356
rect 5311 8316 5356 8344
rect 3145 8307 3203 8313
rect 2866 8276 2872 8288
rect 2827 8248 2872 8276
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3160 8276 3188 8307
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 7422 8347 7480 8353
rect 7422 8344 7434 8347
rect 7300 8316 7434 8344
rect 7300 8288 7328 8316
rect 7422 8313 7434 8316
rect 7468 8313 7480 8347
rect 8128 8344 8156 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9324 8421 9352 8452
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11394 8480 11422 8588
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 17083 8619 17141 8625
rect 17083 8585 17095 8619
rect 17129 8616 17141 8619
rect 19610 8616 19616 8628
rect 17129 8588 19616 8616
rect 17129 8585 17141 8588
rect 17083 8579 17141 8585
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 21324 8588 22385 8616
rect 21324 8576 21330 8588
rect 22373 8585 22385 8588
rect 22419 8585 22431 8619
rect 22738 8616 22744 8628
rect 22699 8588 22744 8616
rect 22373 8579 22431 8585
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 23934 8616 23940 8628
rect 23895 8588 23940 8616
rect 23934 8576 23940 8588
rect 23992 8576 23998 8628
rect 25222 8576 25228 8628
rect 25280 8616 25286 8628
rect 25317 8619 25375 8625
rect 25317 8616 25329 8619
rect 25280 8588 25329 8616
rect 25280 8576 25286 8588
rect 25317 8585 25329 8588
rect 25363 8585 25375 8619
rect 25317 8579 25375 8585
rect 26789 8619 26847 8625
rect 26789 8585 26801 8619
rect 26835 8616 26847 8619
rect 27798 8616 27804 8628
rect 26835 8588 27804 8616
rect 26835 8585 26847 8588
rect 26789 8579 26847 8585
rect 27798 8576 27804 8588
rect 27856 8616 27862 8628
rect 28721 8619 28779 8625
rect 28721 8616 28733 8619
rect 27856 8588 28733 8616
rect 27856 8576 27862 8588
rect 28721 8585 28733 8588
rect 28767 8616 28779 8619
rect 28994 8616 29000 8628
rect 28767 8588 29000 8616
rect 28767 8585 28779 8588
rect 28721 8579 28779 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 32674 8576 32680 8628
rect 32732 8616 32738 8628
rect 32769 8619 32827 8625
rect 32769 8616 32781 8619
rect 32732 8588 32781 8616
rect 32732 8576 32738 8588
rect 32769 8585 32781 8588
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 34057 8619 34115 8625
rect 34057 8585 34069 8619
rect 34103 8616 34115 8619
rect 35618 8616 35624 8628
rect 34103 8588 35624 8616
rect 34103 8585 34115 8588
rect 34057 8579 34115 8585
rect 35618 8576 35624 8588
rect 35676 8616 35682 8628
rect 35989 8619 36047 8625
rect 35989 8616 36001 8619
rect 35676 8588 36001 8616
rect 35676 8576 35682 8588
rect 35989 8585 36001 8588
rect 36035 8585 36047 8619
rect 36262 8616 36268 8628
rect 36223 8588 36268 8616
rect 35989 8579 36047 8585
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 36630 8616 36636 8628
rect 36591 8588 36636 8616
rect 36630 8576 36636 8588
rect 36688 8576 36694 8628
rect 13078 8508 13084 8560
rect 13136 8548 13142 8560
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13136 8520 13829 8548
rect 13136 8508 13142 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 17770 8508 17776 8560
rect 17828 8548 17834 8560
rect 18877 8551 18935 8557
rect 18877 8548 18889 8551
rect 17828 8520 18889 8548
rect 17828 8508 17834 8520
rect 18877 8517 18889 8520
rect 18923 8548 18935 8551
rect 19058 8548 19064 8560
rect 18923 8520 19064 8548
rect 18923 8517 18935 8520
rect 18877 8511 18935 8517
rect 19058 8508 19064 8520
rect 19116 8508 19122 8560
rect 19242 8548 19248 8560
rect 19203 8520 19248 8548
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 20254 8508 20260 8560
rect 20312 8548 20318 8560
rect 28442 8548 28448 8560
rect 20312 8520 28448 8548
rect 20312 8508 20318 8520
rect 28442 8508 28448 8520
rect 28500 8508 28506 8560
rect 35529 8551 35587 8557
rect 35529 8548 35541 8551
rect 34072 8520 35541 8548
rect 34072 8492 34100 8520
rect 35529 8517 35541 8520
rect 35575 8548 35587 8551
rect 35894 8548 35900 8560
rect 35575 8520 35900 8548
rect 35575 8517 35587 8520
rect 35529 8511 35587 8517
rect 35894 8508 35900 8520
rect 35952 8508 35958 8560
rect 10919 8452 11422 8480
rect 11517 8483 11575 8489
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11974 8480 11980 8492
rect 11563 8452 11980 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 11974 8440 11980 8452
rect 12032 8480 12038 8492
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 12032 8452 12817 8480
rect 12032 8440 12038 8452
rect 12805 8449 12817 8452
rect 12851 8480 12863 8483
rect 16482 8480 16488 8492
rect 12851 8452 16488 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 18046 8480 18052 8492
rect 17911 8452 18052 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 19702 8480 19708 8492
rect 18371 8452 19708 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20070 8480 20076 8492
rect 19935 8452 20076 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 21450 8480 21456 8492
rect 21411 8452 21456 8480
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 27706 8480 27712 8492
rect 21784 8452 24348 8480
rect 27667 8452 27712 8480
rect 21784 8440 21790 8452
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8720 8384 8861 8412
rect 8720 8372 8726 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 14036 8415 14094 8421
rect 14036 8381 14048 8415
rect 14082 8381 14094 8415
rect 15194 8412 15200 8424
rect 15155 8384 15200 8412
rect 14036 8375 14094 8381
rect 10962 8344 10968 8356
rect 8128 8316 8984 8344
rect 10923 8316 10968 8344
rect 7422 8307 7480 8313
rect 8956 8288 8984 8316
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 12342 8304 12348 8356
rect 12400 8344 12406 8356
rect 12529 8347 12587 8353
rect 12529 8344 12541 8347
rect 12400 8316 12541 8344
rect 12400 8304 12406 8316
rect 12529 8313 12541 8316
rect 12575 8313 12587 8347
rect 12529 8307 12587 8313
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8344 12679 8347
rect 12894 8344 12900 8356
rect 12667 8316 12900 8344
rect 12667 8313 12679 8316
rect 12621 8307 12679 8313
rect 3418 8276 3424 8288
rect 3160 8248 3424 8276
rect 3418 8236 3424 8248
rect 3476 8276 3482 8288
rect 4246 8276 4252 8288
rect 3476 8248 4252 8276
rect 3476 8236 3482 8248
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4982 8276 4988 8288
rect 4943 8248 4988 8276
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 6181 8279 6239 8285
rect 6181 8276 6193 8279
rect 5776 8248 6193 8276
rect 5776 8236 5782 8248
rect 6181 8245 6193 8248
rect 6227 8245 6239 8279
rect 6181 8239 6239 8245
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 7282 8276 7288 8288
rect 6687 8248 7288 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8938 8276 8944 8288
rect 8899 8248 8944 8276
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 11885 8279 11943 8285
rect 11885 8245 11897 8279
rect 11931 8276 11943 8279
rect 11974 8276 11980 8288
rect 11931 8248 11980 8276
rect 11931 8245 11943 8248
rect 11885 8239 11943 8245
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 12253 8279 12311 8285
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12636 8276 12664 8307
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 12299 8248 12664 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 13078 8236 13084 8288
rect 13136 8276 13142 8288
rect 14051 8276 14079 8375
rect 15194 8372 15200 8384
rect 15252 8412 15258 8424
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 15252 8384 16773 8412
rect 15252 8372 15258 8384
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 16761 8375 16819 8381
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 16980 8415 17038 8421
rect 16980 8412 16992 8415
rect 16908 8384 16992 8412
rect 16908 8372 16914 8384
rect 16980 8381 16992 8384
rect 17026 8381 17038 8415
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 16980 8375 17038 8381
rect 20640 8384 21189 8412
rect 14139 8347 14197 8353
rect 14139 8313 14151 8347
rect 14185 8344 14197 8347
rect 14642 8344 14648 8356
rect 14185 8316 14648 8344
rect 14185 8313 14197 8316
rect 14139 8307 14197 8313
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 18414 8344 18420 8356
rect 18375 8316 18420 8344
rect 18414 8304 18420 8316
rect 18472 8304 18478 8356
rect 19981 8347 20039 8353
rect 19981 8313 19993 8347
rect 20027 8313 20039 8347
rect 19981 8307 20039 8313
rect 14553 8279 14611 8285
rect 14553 8276 14565 8279
rect 13136 8248 14565 8276
rect 13136 8236 13142 8248
rect 14553 8245 14565 8248
rect 14599 8276 14611 8279
rect 14734 8276 14740 8288
rect 14599 8248 14740 8276
rect 14599 8245 14611 8248
rect 14553 8239 14611 8245
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 15105 8279 15163 8285
rect 15105 8245 15117 8279
rect 15151 8276 15163 8279
rect 15565 8279 15623 8285
rect 15565 8276 15577 8279
rect 15151 8248 15577 8276
rect 15151 8245 15163 8248
rect 15105 8239 15163 8245
rect 15565 8245 15577 8248
rect 15611 8276 15623 8279
rect 15654 8276 15660 8288
rect 15611 8248 15660 8276
rect 15611 8245 15623 8248
rect 15565 8239 15623 8245
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 16114 8276 16120 8288
rect 16075 8248 16120 8276
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 16485 8279 16543 8285
rect 16485 8245 16497 8279
rect 16531 8276 16543 8279
rect 16942 8276 16948 8288
rect 16531 8248 16948 8276
rect 16531 8245 16543 8248
rect 16485 8239 16543 8245
rect 16942 8236 16948 8248
rect 17000 8236 17006 8288
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 19610 8276 19616 8288
rect 19571 8248 19616 8276
rect 19610 8236 19616 8248
rect 19668 8276 19674 8288
rect 19996 8276 20024 8307
rect 20640 8276 20668 8384
rect 21177 8381 21189 8384
rect 21223 8412 21235 8415
rect 21266 8412 21272 8424
rect 21223 8384 21272 8412
rect 21223 8381 21235 8384
rect 21177 8375 21235 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 23382 8372 23388 8424
rect 23440 8412 23446 8424
rect 23492 8412 23520 8452
rect 24320 8424 24348 8452
rect 27706 8440 27712 8452
rect 27764 8440 27770 8492
rect 29178 8440 29184 8492
rect 29236 8480 29242 8492
rect 29641 8483 29699 8489
rect 29641 8480 29653 8483
rect 29236 8452 29653 8480
rect 29236 8440 29242 8452
rect 29641 8449 29653 8452
rect 29687 8449 29699 8483
rect 33318 8480 33324 8492
rect 33279 8452 33324 8480
rect 29641 8443 29699 8449
rect 33318 8440 33324 8452
rect 33376 8440 33382 8492
rect 33965 8483 34023 8489
rect 33965 8449 33977 8483
rect 34011 8480 34023 8483
rect 34054 8480 34060 8492
rect 34011 8452 34060 8480
rect 34011 8449 34023 8452
rect 33965 8443 34023 8449
rect 34054 8440 34060 8452
rect 34112 8440 34118 8492
rect 34974 8480 34980 8492
rect 34887 8452 34980 8480
rect 34974 8440 34980 8452
rect 35032 8480 35038 8492
rect 37691 8483 37749 8489
rect 37691 8480 37703 8483
rect 35032 8452 37703 8480
rect 35032 8440 35038 8452
rect 37691 8449 37703 8452
rect 37737 8449 37749 8483
rect 37691 8443 37749 8449
rect 24302 8412 24308 8424
rect 23440 8384 23520 8412
rect 24263 8384 24308 8412
rect 23440 8372 23446 8384
rect 24302 8372 24308 8384
rect 24360 8372 24366 8424
rect 24762 8412 24768 8424
rect 24723 8384 24768 8412
rect 24762 8372 24768 8384
rect 24820 8372 24826 8424
rect 25041 8415 25099 8421
rect 25041 8381 25053 8415
rect 25087 8412 25099 8415
rect 25866 8412 25872 8424
rect 25087 8384 25872 8412
rect 25087 8381 25099 8384
rect 25041 8375 25099 8381
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 31205 8415 31263 8421
rect 31205 8381 31217 8415
rect 31251 8412 31263 8415
rect 31386 8412 31392 8424
rect 31251 8384 31392 8412
rect 31251 8381 31263 8384
rect 31205 8375 31263 8381
rect 31386 8372 31392 8384
rect 31444 8372 31450 8424
rect 32125 8415 32183 8421
rect 32125 8381 32137 8415
rect 32171 8412 32183 8415
rect 33134 8412 33140 8424
rect 32171 8384 33140 8412
rect 32171 8381 32183 8384
rect 32125 8375 32183 8381
rect 33106 8372 33140 8384
rect 33192 8372 33198 8424
rect 36449 8415 36507 8421
rect 36449 8381 36461 8415
rect 36495 8412 36507 8415
rect 37604 8415 37662 8421
rect 36495 8384 37136 8412
rect 36495 8381 36507 8384
rect 36449 8375 36507 8381
rect 21542 8344 21548 8356
rect 20824 8316 21548 8344
rect 20824 8288 20852 8316
rect 21542 8304 21548 8316
rect 21600 8304 21606 8356
rect 22097 8347 22155 8353
rect 22097 8313 22109 8347
rect 22143 8344 22155 8347
rect 22186 8344 22192 8356
rect 22143 8316 22192 8344
rect 22143 8313 22155 8316
rect 22097 8307 22155 8313
rect 22186 8304 22192 8316
rect 22244 8304 22250 8356
rect 23477 8347 23535 8353
rect 23477 8313 23489 8347
rect 23523 8344 23535 8347
rect 24780 8344 24808 8372
rect 23523 8316 24808 8344
rect 26231 8347 26289 8353
rect 23523 8313 23535 8316
rect 23477 8307 23535 8313
rect 26231 8313 26243 8347
rect 26277 8313 26289 8347
rect 27798 8344 27804 8356
rect 27759 8316 27804 8344
rect 26231 8307 26289 8313
rect 20806 8276 20812 8288
rect 19668 8248 20668 8276
rect 20767 8248 20812 8276
rect 19668 8236 19674 8248
rect 20806 8236 20812 8248
rect 20864 8236 20870 8288
rect 25777 8279 25835 8285
rect 25777 8245 25789 8279
rect 25823 8276 25835 8279
rect 26252 8276 26280 8307
rect 27798 8304 27804 8316
rect 27856 8304 27862 8356
rect 28353 8347 28411 8353
rect 28353 8313 28365 8347
rect 28399 8344 28411 8347
rect 28534 8344 28540 8356
rect 28399 8316 28540 8344
rect 28399 8313 28411 8316
rect 28353 8307 28411 8313
rect 28534 8304 28540 8316
rect 28592 8304 28598 8356
rect 29362 8344 29368 8356
rect 29323 8316 29368 8344
rect 29362 8304 29368 8316
rect 29420 8304 29426 8356
rect 29457 8347 29515 8353
rect 29457 8313 29469 8347
rect 29503 8313 29515 8347
rect 29457 8307 29515 8313
rect 31113 8347 31171 8353
rect 31113 8313 31125 8347
rect 31159 8344 31171 8347
rect 31526 8347 31584 8353
rect 31526 8344 31538 8347
rect 31159 8316 31538 8344
rect 31159 8313 31171 8316
rect 31113 8307 31171 8313
rect 31526 8313 31538 8316
rect 31572 8344 31584 8347
rect 32582 8344 32588 8356
rect 31572 8316 32588 8344
rect 31572 8313 31584 8316
rect 31526 8307 31584 8313
rect 26786 8276 26792 8288
rect 25823 8248 26792 8276
rect 25823 8245 25835 8248
rect 25777 8239 25835 8245
rect 26786 8236 26792 8248
rect 26844 8236 26850 8288
rect 26970 8236 26976 8288
rect 27028 8276 27034 8288
rect 27249 8279 27307 8285
rect 27249 8276 27261 8279
rect 27028 8248 27261 8276
rect 27028 8236 27034 8248
rect 27249 8245 27261 8248
rect 27295 8276 27307 8279
rect 27522 8276 27528 8288
rect 27295 8248 27528 8276
rect 27295 8245 27307 8248
rect 27249 8239 27307 8245
rect 27522 8236 27528 8248
rect 27580 8276 27586 8288
rect 28997 8279 29055 8285
rect 28997 8276 29009 8279
rect 27580 8248 29009 8276
rect 27580 8236 27586 8248
rect 28997 8245 29009 8248
rect 29043 8276 29055 8279
rect 29472 8276 29500 8307
rect 32582 8304 32588 8316
rect 32640 8304 32646 8356
rect 33106 8344 33134 8372
rect 33413 8347 33471 8353
rect 33413 8344 33425 8347
rect 33106 8316 33425 8344
rect 33413 8313 33425 8316
rect 33459 8344 33471 8347
rect 34057 8347 34115 8353
rect 34057 8344 34069 8347
rect 33459 8316 34069 8344
rect 33459 8313 33471 8316
rect 33413 8307 33471 8313
rect 34057 8313 34069 8316
rect 34103 8313 34115 8347
rect 34057 8307 34115 8313
rect 34606 8304 34612 8356
rect 34664 8344 34670 8356
rect 34701 8347 34759 8353
rect 34701 8344 34713 8347
rect 34664 8316 34713 8344
rect 34664 8304 34670 8316
rect 34701 8313 34713 8316
rect 34747 8344 34759 8347
rect 35069 8347 35127 8353
rect 35069 8344 35081 8347
rect 34747 8316 35081 8344
rect 34747 8313 34759 8316
rect 34701 8307 34759 8313
rect 35069 8313 35081 8316
rect 35115 8313 35127 8347
rect 35069 8307 35127 8313
rect 30374 8276 30380 8288
rect 29043 8248 29500 8276
rect 30335 8248 30380 8276
rect 29043 8245 29055 8248
rect 28997 8239 29055 8245
rect 30374 8236 30380 8248
rect 30432 8236 30438 8288
rect 32306 8236 32312 8288
rect 32364 8276 32370 8288
rect 32401 8279 32459 8285
rect 32401 8276 32413 8279
rect 32364 8248 32413 8276
rect 32364 8236 32370 8248
rect 32401 8245 32413 8248
rect 32447 8245 32459 8279
rect 34238 8276 34244 8288
rect 34199 8248 34244 8276
rect 32401 8239 32459 8245
rect 34238 8236 34244 8248
rect 34296 8236 34302 8288
rect 34514 8236 34520 8288
rect 34572 8276 34578 8288
rect 36464 8276 36492 8375
rect 37108 8285 37136 8384
rect 37604 8381 37616 8415
rect 37650 8412 37662 8415
rect 38010 8412 38016 8424
rect 37650 8384 38016 8412
rect 37650 8381 37662 8384
rect 37604 8375 37662 8381
rect 38010 8372 38016 8384
rect 38068 8372 38074 8424
rect 34572 8248 36492 8276
rect 37093 8279 37151 8285
rect 34572 8236 34578 8248
rect 37093 8245 37105 8279
rect 37139 8276 37151 8279
rect 37366 8276 37372 8288
rect 37139 8248 37372 8276
rect 37139 8245 37151 8248
rect 37093 8239 37151 8245
rect 37366 8236 37372 8248
rect 37424 8236 37430 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 2041 8075 2099 8081
rect 2041 8072 2053 8075
rect 1636 8044 2053 8072
rect 1636 8032 1642 8044
rect 2041 8041 2053 8044
rect 2087 8072 2099 8075
rect 2866 8072 2872 8084
rect 2087 8044 2872 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 3418 8072 3424 8084
rect 3099 8044 3424 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 3697 8075 3755 8081
rect 3697 8072 3709 8075
rect 3660 8044 3709 8072
rect 3660 8032 3666 8044
rect 3697 8041 3709 8044
rect 3743 8041 3755 8075
rect 3697 8035 3755 8041
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 6730 8072 6736 8084
rect 6687 8044 6736 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 6972 8044 7665 8072
rect 6972 8032 6978 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 8018 8072 8024 8084
rect 7979 8044 8024 8072
rect 7653 8035 7711 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8938 8072 8944 8084
rect 8435 8044 8944 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 10594 8072 10600 8084
rect 10551 8044 10600 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 10962 8072 10968 8084
rect 10919 8044 10968 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 10962 8032 10968 8044
rect 11020 8072 11026 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11020 8044 11897 8072
rect 11020 8032 11026 8044
rect 11885 8041 11897 8044
rect 11931 8072 11943 8075
rect 12526 8072 12532 8084
rect 11931 8044 12532 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15654 8072 15660 8084
rect 15615 8044 15660 8072
rect 15013 8035 15071 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 17402 8072 17408 8084
rect 16255 8044 17408 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 18969 8075 19027 8081
rect 18969 8041 18981 8075
rect 19015 8072 19027 8075
rect 19242 8072 19248 8084
rect 19015 8044 19248 8072
rect 19015 8041 19027 8044
rect 18969 8035 19027 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 19797 8075 19855 8081
rect 19797 8072 19809 8075
rect 19760 8044 19809 8072
rect 19760 8032 19766 8044
rect 19797 8041 19809 8044
rect 19843 8041 19855 8075
rect 22094 8072 22100 8084
rect 22055 8044 22100 8072
rect 19797 8035 19855 8041
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 23661 8075 23719 8081
rect 23661 8072 23673 8075
rect 22244 8044 23673 8072
rect 22244 8032 22250 8044
rect 23661 8041 23673 8044
rect 23707 8072 23719 8075
rect 23750 8072 23756 8084
rect 23707 8044 23756 8072
rect 23707 8041 23719 8044
rect 23661 8035 23719 8041
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 24302 8072 24308 8084
rect 24263 8044 24308 8072
rect 24302 8032 24308 8044
rect 24360 8032 24366 8084
rect 25866 8072 25872 8084
rect 25827 8044 25872 8072
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 26786 8032 26792 8084
rect 26844 8072 26850 8084
rect 26881 8075 26939 8081
rect 26881 8072 26893 8075
rect 26844 8044 26893 8072
rect 26844 8032 26850 8044
rect 26881 8041 26893 8044
rect 26927 8041 26939 8075
rect 27430 8072 27436 8084
rect 27391 8044 27436 8072
rect 26881 8035 26939 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 27801 8075 27859 8081
rect 27801 8041 27813 8075
rect 27847 8072 27859 8075
rect 27982 8072 27988 8084
rect 27847 8044 27988 8072
rect 27847 8041 27859 8044
rect 27801 8035 27859 8041
rect 27982 8032 27988 8044
rect 28040 8032 28046 8084
rect 33413 8075 33471 8081
rect 28178 8044 30512 8072
rect 1670 8004 1676 8016
rect 1631 7976 1676 8004
rect 1670 7964 1676 7976
rect 1728 7964 1734 8016
rect 2314 7964 2320 8016
rect 2372 8004 2378 8016
rect 2454 8007 2512 8013
rect 2454 8004 2466 8007
rect 2372 7976 2466 8004
rect 2372 7964 2378 7976
rect 2454 7973 2466 7976
rect 2500 7973 2512 8007
rect 4246 8004 4252 8016
rect 4207 7976 4252 8004
rect 2454 7967 2512 7973
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 4801 8007 4859 8013
rect 4801 7973 4813 8007
rect 4847 8004 4859 8007
rect 5258 8004 5264 8016
rect 4847 7976 5264 8004
rect 4847 7973 4859 7976
rect 4801 7967 4859 7973
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2222 7936 2228 7948
rect 2179 7908 2228 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 6748 7945 6776 8032
rect 7095 8007 7153 8013
rect 7095 7973 7107 8007
rect 7141 8004 7153 8007
rect 7282 8004 7288 8016
rect 7141 7976 7288 8004
rect 7141 7973 7153 7976
rect 7095 7967 7153 7973
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 5629 7939 5687 7945
rect 5629 7936 5641 7939
rect 4948 7908 5641 7936
rect 4948 7896 4954 7908
rect 5629 7905 5641 7908
rect 5675 7936 5687 7939
rect 6733 7939 6791 7945
rect 5675 7908 6408 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4338 7868 4344 7880
rect 4203 7840 4344 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 6380 7812 6408 7908
rect 6733 7905 6745 7939
rect 6779 7905 6791 7939
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 6733 7899 6791 7905
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 9988 7939 10046 7945
rect 9988 7905 10000 7939
rect 10034 7905 10046 7939
rect 10612 7936 10640 8032
rect 11146 7964 11152 8016
rect 11204 8004 11210 8016
rect 11286 8007 11344 8013
rect 11286 8004 11298 8007
rect 11204 7976 11298 8004
rect 11204 7964 11210 7976
rect 11286 7973 11298 7976
rect 11332 7973 11344 8007
rect 12894 8004 12900 8016
rect 12855 7976 12900 8004
rect 11286 7967 11344 7973
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 13449 8007 13507 8013
rect 13449 7973 13461 8007
rect 13495 8004 13507 8007
rect 13538 8004 13544 8016
rect 13495 7976 13544 8004
rect 13495 7973 13507 7976
rect 13449 7967 13507 7973
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 16482 8004 16488 8016
rect 16443 7976 16488 8004
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 17126 8004 17132 8016
rect 17087 7976 17132 8004
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 17770 8004 17776 8016
rect 17276 7976 17321 8004
rect 17731 7976 17776 8004
rect 17276 7964 17282 7976
rect 17770 7964 17776 7976
rect 17828 7964 17834 8016
rect 21266 8004 21272 8016
rect 21227 7976 21272 8004
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 21821 8007 21879 8013
rect 21821 7973 21833 8007
rect 21867 8004 21879 8007
rect 22204 8004 22232 8032
rect 22830 8004 22836 8016
rect 21867 7976 22232 8004
rect 22791 7976 22836 8004
rect 21867 7973 21879 7976
rect 21821 7967 21879 7973
rect 22830 7964 22836 7976
rect 22888 7964 22894 8016
rect 25222 7964 25228 8016
rect 25280 8004 25286 8016
rect 25280 7976 25589 8004
rect 25280 7964 25286 7976
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 10612 7908 10977 7936
rect 9988 7899 10046 7905
rect 10965 7905 10977 7908
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 10003 7812 10031 7899
rect 12342 7896 12348 7948
rect 12400 7936 12406 7948
rect 12529 7939 12587 7945
rect 12529 7936 12541 7939
rect 12400 7908 12541 7936
rect 12400 7896 12406 7908
rect 12529 7905 12541 7908
rect 12575 7905 12587 7939
rect 12529 7899 12587 7905
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 15068 7908 15301 7936
rect 15068 7896 15074 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 18601 7939 18659 7945
rect 18601 7905 18613 7939
rect 18647 7936 18659 7939
rect 18690 7936 18696 7948
rect 18647 7908 18696 7936
rect 18647 7905 18659 7908
rect 18601 7899 18659 7905
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 20806 7936 20812 7948
rect 19567 7908 20812 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 20806 7896 20812 7908
rect 20864 7896 20870 7948
rect 24670 7896 24676 7948
rect 24728 7936 24734 7948
rect 24857 7939 24915 7945
rect 24857 7936 24869 7939
rect 24728 7908 24869 7936
rect 24728 7896 24734 7908
rect 24857 7905 24869 7908
rect 24903 7905 24915 7939
rect 25406 7936 25412 7948
rect 25367 7908 25412 7936
rect 24857 7899 24915 7905
rect 25406 7896 25412 7908
rect 25464 7896 25470 7948
rect 25561 7936 25589 7976
rect 27338 7964 27344 8016
rect 27396 8004 27402 8016
rect 28077 8007 28135 8013
rect 28077 8004 28089 8007
rect 27396 7976 28089 8004
rect 27396 7964 27402 7976
rect 28077 7973 28089 7976
rect 28123 7973 28135 8007
rect 28077 7967 28135 7973
rect 28178 7936 28206 8044
rect 28626 8004 28632 8016
rect 28587 7976 28632 8004
rect 28626 7964 28632 7976
rect 28684 7964 28690 8016
rect 30484 7948 30512 8044
rect 33413 8041 33425 8075
rect 33459 8072 33471 8075
rect 33502 8072 33508 8084
rect 33459 8044 33508 8072
rect 33459 8041 33471 8044
rect 33413 8035 33471 8041
rect 33502 8032 33508 8044
rect 33560 8032 33566 8084
rect 33962 8032 33968 8084
rect 34020 8072 34026 8084
rect 34333 8075 34391 8081
rect 34333 8072 34345 8075
rect 34020 8044 34345 8072
rect 34020 8032 34026 8044
rect 34333 8041 34345 8044
rect 34379 8041 34391 8075
rect 34333 8035 34391 8041
rect 34422 8032 34428 8084
rect 34480 8072 34486 8084
rect 35894 8072 35900 8084
rect 34480 8044 35525 8072
rect 35855 8044 35900 8072
rect 34480 8032 34486 8044
rect 32487 8007 32545 8013
rect 32487 7973 32499 8007
rect 32533 8004 32545 8007
rect 32582 8004 32588 8016
rect 32533 7976 32588 8004
rect 32533 7973 32545 7976
rect 32487 7967 32545 7973
rect 32582 7964 32588 7976
rect 32640 7964 32646 8016
rect 33042 7964 33048 8016
rect 33100 8004 33106 8016
rect 34238 8004 34244 8016
rect 33100 7976 34244 8004
rect 33100 7964 33106 7976
rect 34238 7964 34244 7976
rect 34296 7964 34302 8016
rect 34698 7964 34704 8016
rect 34756 8004 34762 8016
rect 35069 8007 35127 8013
rect 35069 8004 35081 8007
rect 34756 7976 35081 8004
rect 34756 7964 34762 7976
rect 35069 7973 35081 7976
rect 35115 7973 35127 8007
rect 35497 8004 35525 8044
rect 35894 8032 35900 8044
rect 35952 8032 35958 8084
rect 38010 8004 38016 8016
rect 35497 7976 38016 8004
rect 35069 7967 35127 7973
rect 38010 7964 38016 7976
rect 38068 7964 38074 8016
rect 30466 7936 30472 7948
rect 25561 7908 28206 7936
rect 30427 7908 30472 7936
rect 30466 7896 30472 7908
rect 30524 7896 30530 7948
rect 31021 7939 31079 7945
rect 31021 7905 31033 7939
rect 31067 7936 31079 7939
rect 31294 7936 31300 7948
rect 31067 7908 31300 7936
rect 31067 7905 31079 7908
rect 31021 7899 31079 7905
rect 31294 7896 31300 7908
rect 31352 7896 31358 7948
rect 33908 7939 33966 7945
rect 33908 7936 33920 7939
rect 33106 7908 33920 7936
rect 10091 7871 10149 7877
rect 10091 7837 10103 7871
rect 10137 7868 10149 7871
rect 11698 7868 11704 7880
rect 10137 7840 11704 7868
rect 10137 7837 10149 7840
rect 10091 7831 10149 7837
rect 11698 7828 11704 7840
rect 11756 7868 11762 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11756 7840 12173 7868
rect 11756 7828 11762 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 12676 7840 12817 7868
rect 12676 7828 12682 7840
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 19978 7868 19984 7880
rect 14792 7840 19984 7868
rect 14792 7828 14798 7840
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20763 7840 21189 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 21177 7837 21189 7840
rect 21223 7868 21235 7871
rect 21818 7868 21824 7880
rect 21223 7840 21824 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 21818 7828 21824 7840
rect 21876 7828 21882 7880
rect 22738 7868 22744 7880
rect 22699 7840 22744 7868
rect 22738 7828 22744 7840
rect 22796 7828 22802 7880
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7868 23443 7871
rect 24118 7868 24124 7880
rect 23431 7840 24124 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 24118 7828 24124 7840
rect 24176 7828 24182 7880
rect 24762 7868 24768 7880
rect 24675 7840 24768 7868
rect 24762 7828 24768 7840
rect 24820 7868 24826 7880
rect 25424 7868 25452 7896
rect 24820 7840 25452 7868
rect 25593 7871 25651 7877
rect 24820 7828 24826 7840
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 26513 7871 26571 7877
rect 26513 7868 26525 7871
rect 25639 7840 26525 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 26513 7837 26525 7840
rect 26559 7868 26571 7871
rect 27614 7868 27620 7880
rect 26559 7840 27620 7868
rect 26559 7837 26571 7840
rect 26513 7831 26571 7837
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 28534 7868 28540 7880
rect 28495 7840 28540 7868
rect 28534 7828 28540 7840
rect 28592 7828 28598 7880
rect 29181 7871 29239 7877
rect 29181 7837 29193 7871
rect 29227 7868 29239 7871
rect 30006 7868 30012 7880
rect 29227 7840 30012 7868
rect 29227 7837 29239 7840
rect 29181 7831 29239 7837
rect 30006 7828 30012 7840
rect 30064 7828 30070 7880
rect 31205 7871 31263 7877
rect 31205 7837 31217 7871
rect 31251 7868 31263 7871
rect 32125 7871 32183 7877
rect 32125 7868 32137 7871
rect 31251 7840 32137 7868
rect 31251 7837 31263 7840
rect 31205 7831 31263 7837
rect 32125 7837 32137 7840
rect 32171 7868 32183 7871
rect 32490 7868 32496 7880
rect 32171 7840 32496 7868
rect 32171 7837 32183 7840
rect 32125 7831 32183 7837
rect 32490 7828 32496 7840
rect 32548 7828 32554 7880
rect 5810 7800 5816 7812
rect 5771 7772 5816 7800
rect 5810 7760 5816 7772
rect 5868 7760 5874 7812
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 9122 7800 9128 7812
rect 6420 7772 9128 7800
rect 6420 7760 6426 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9950 7800 9956 7812
rect 9898 7772 9956 7800
rect 9950 7760 9956 7772
rect 10008 7800 10031 7812
rect 13078 7800 13084 7812
rect 10008 7772 13084 7800
rect 10008 7760 10014 7772
rect 13078 7760 13084 7772
rect 13136 7760 13142 7812
rect 16850 7800 16856 7812
rect 13786 7772 16856 7800
rect 5258 7732 5264 7744
rect 5219 7704 5264 7732
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6273 7735 6331 7741
rect 6273 7732 6285 7735
rect 5960 7704 6285 7732
rect 5960 7692 5966 7704
rect 6273 7701 6285 7704
rect 6319 7732 6331 7735
rect 6638 7732 6644 7744
rect 6319 7704 6644 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 8662 7732 8668 7744
rect 8623 7704 8668 7732
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 13786 7732 13814 7772
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 24578 7760 24584 7812
rect 24636 7800 24642 7812
rect 30282 7800 30288 7812
rect 24636 7772 30288 7800
rect 24636 7760 24642 7772
rect 30282 7760 30288 7772
rect 30340 7760 30346 7812
rect 30374 7760 30380 7812
rect 30432 7800 30438 7812
rect 33106 7800 33134 7908
rect 33908 7905 33920 7908
rect 33954 7936 33966 7939
rect 34146 7936 34152 7948
rect 33954 7908 34152 7936
rect 33954 7905 33966 7908
rect 33908 7899 33966 7905
rect 34146 7896 34152 7908
rect 34204 7896 34210 7948
rect 36446 7936 36452 7948
rect 36407 7908 36452 7936
rect 36446 7896 36452 7908
rect 36504 7896 36510 7948
rect 34974 7868 34980 7880
rect 34935 7840 34980 7868
rect 34974 7828 34980 7840
rect 35032 7828 35038 7880
rect 35618 7868 35624 7880
rect 35579 7840 35624 7868
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 30432 7772 33134 7800
rect 34011 7803 34069 7809
rect 30432 7760 30438 7772
rect 34011 7769 34023 7803
rect 34057 7800 34069 7803
rect 36354 7800 36360 7812
rect 34057 7772 36360 7800
rect 34057 7769 34069 7772
rect 34011 7763 34069 7769
rect 36354 7760 36360 7772
rect 36412 7760 36418 7812
rect 36630 7800 36636 7812
rect 36591 7772 36636 7800
rect 36630 7760 36636 7772
rect 36688 7760 36694 7812
rect 13596 7704 13814 7732
rect 18325 7735 18383 7741
rect 13596 7692 13602 7704
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18414 7732 18420 7744
rect 18371 7704 18420 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18414 7692 18420 7704
rect 18472 7732 18478 7744
rect 18874 7732 18880 7744
rect 18472 7704 18880 7732
rect 18472 7692 18478 7704
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 27522 7692 27528 7744
rect 27580 7732 27586 7744
rect 29362 7732 29368 7744
rect 27580 7704 29368 7732
rect 27580 7692 27586 7704
rect 29362 7692 29368 7704
rect 29420 7732 29426 7744
rect 29457 7735 29515 7741
rect 29457 7732 29469 7735
rect 29420 7704 29469 7732
rect 29420 7692 29426 7704
rect 29457 7701 29469 7704
rect 29503 7701 29515 7735
rect 33042 7732 33048 7744
rect 33003 7704 33048 7732
rect 29457 7695 29515 7701
rect 33042 7692 33048 7704
rect 33100 7692 33106 7744
rect 34793 7735 34851 7741
rect 34793 7701 34805 7735
rect 34839 7732 34851 7735
rect 34974 7732 34980 7744
rect 34839 7704 34980 7732
rect 34839 7701 34851 7704
rect 34793 7695 34851 7701
rect 34974 7692 34980 7704
rect 35032 7732 35038 7744
rect 36814 7732 36820 7744
rect 35032 7704 36820 7732
rect 35032 7692 35038 7704
rect 36814 7692 36820 7704
rect 36872 7692 36878 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3326 7528 3332 7540
rect 3191 7500 3332 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3326 7488 3332 7500
rect 3384 7528 3390 7540
rect 4246 7528 4252 7540
rect 3384 7500 4252 7528
rect 3384 7488 3390 7500
rect 4246 7488 4252 7500
rect 4304 7528 4310 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 4304 7500 4905 7528
rect 4304 7488 4310 7500
rect 4893 7497 4905 7500
rect 4939 7497 4951 7531
rect 4893 7491 4951 7497
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 5316 7500 7757 7528
rect 5316 7488 5322 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 9950 7528 9956 7540
rect 9911 7500 9956 7528
rect 7745 7491 7803 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 12894 7528 12900 7540
rect 11563 7500 12900 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 12894 7488 12900 7500
rect 12952 7528 12958 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 12952 7500 13461 7528
rect 12952 7488 12958 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 15473 7531 15531 7537
rect 15473 7497 15485 7531
rect 15519 7528 15531 7531
rect 15654 7528 15660 7540
rect 15519 7500 15660 7528
rect 15519 7497 15531 7500
rect 15473 7491 15531 7497
rect 15654 7488 15660 7500
rect 15712 7528 15718 7540
rect 16942 7528 16948 7540
rect 15712 7500 16948 7528
rect 15712 7488 15718 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17405 7531 17463 7537
rect 17405 7528 17417 7531
rect 17184 7500 17417 7528
rect 17184 7488 17190 7500
rect 17405 7497 17417 7500
rect 17451 7497 17463 7531
rect 17405 7491 17463 7497
rect 18969 7531 19027 7537
rect 18969 7497 18981 7531
rect 19015 7528 19027 7531
rect 19610 7528 19616 7540
rect 19015 7500 19616 7528
rect 19015 7497 19027 7500
rect 18969 7491 19027 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 20901 7531 20959 7537
rect 20901 7497 20913 7531
rect 20947 7528 20959 7531
rect 21266 7528 21272 7540
rect 20947 7500 21272 7528
rect 20947 7497 20959 7500
rect 20901 7491 20959 7497
rect 21266 7488 21272 7500
rect 21324 7528 21330 7540
rect 21545 7531 21603 7537
rect 21545 7528 21557 7531
rect 21324 7500 21557 7528
rect 21324 7488 21330 7500
rect 21545 7497 21557 7500
rect 21591 7528 21603 7531
rect 21910 7528 21916 7540
rect 21591 7500 21916 7528
rect 21591 7497 21603 7500
rect 21545 7491 21603 7497
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 24857 7531 24915 7537
rect 24857 7528 24869 7531
rect 24728 7500 24869 7528
rect 24728 7488 24734 7500
rect 24857 7497 24869 7500
rect 24903 7497 24915 7531
rect 26970 7528 26976 7540
rect 26931 7500 26976 7528
rect 24857 7491 24915 7497
rect 26970 7488 26976 7500
rect 27028 7488 27034 7540
rect 27614 7528 27620 7540
rect 27575 7500 27620 7528
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 28626 7528 28632 7540
rect 28587 7500 28632 7528
rect 28626 7488 28632 7500
rect 28684 7488 28690 7540
rect 32490 7528 32496 7540
rect 32451 7500 32496 7528
rect 32490 7488 32496 7500
rect 32548 7488 32554 7540
rect 33042 7528 33048 7540
rect 33003 7500 33048 7528
rect 33042 7488 33048 7500
rect 33100 7488 33106 7540
rect 34146 7488 34152 7540
rect 34204 7528 34210 7540
rect 34241 7531 34299 7537
rect 34241 7528 34253 7531
rect 34204 7500 34253 7528
rect 34204 7488 34210 7500
rect 34241 7497 34253 7500
rect 34287 7528 34299 7531
rect 36265 7531 36323 7537
rect 36265 7528 36277 7531
rect 34287 7500 36277 7528
rect 34287 7497 34299 7500
rect 34241 7491 34299 7497
rect 36265 7497 36277 7500
rect 36311 7528 36323 7531
rect 36446 7528 36452 7540
rect 36311 7500 36452 7528
rect 36311 7497 36323 7500
rect 36265 7491 36323 7497
rect 36446 7488 36452 7500
rect 36504 7488 36510 7540
rect 2222 7420 2228 7472
rect 2280 7460 2286 7472
rect 3789 7463 3847 7469
rect 3789 7460 3801 7463
rect 2280 7432 3801 7460
rect 2280 7420 2286 7432
rect 3789 7429 3801 7432
rect 3835 7429 3847 7463
rect 3789 7423 3847 7429
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 4157 7463 4215 7469
rect 4157 7460 4169 7463
rect 3936 7432 4169 7460
rect 3936 7420 3942 7432
rect 4157 7429 4169 7432
rect 4203 7429 4215 7463
rect 4157 7423 4215 7429
rect 5077 7463 5135 7469
rect 5077 7429 5089 7463
rect 5123 7460 5135 7463
rect 9490 7460 9496 7472
rect 5123 7432 9496 7460
rect 5123 7429 5135 7432
rect 5077 7423 5135 7429
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 12618 7420 12624 7472
rect 12676 7460 12682 7472
rect 13817 7463 13875 7469
rect 13817 7460 13829 7463
rect 12676 7432 13829 7460
rect 12676 7420 12682 7432
rect 13817 7429 13829 7432
rect 13863 7429 13875 7463
rect 17770 7460 17776 7472
rect 13817 7423 13875 7429
rect 15856 7432 17776 7460
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 1728 7364 4016 7392
rect 1728 7352 1734 7364
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 3142 7324 3148 7336
rect 2271 7296 3148 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 3142 7284 3148 7296
rect 3200 7324 3206 7336
rect 3988 7333 4016 7364
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 4120 7364 5273 7392
rect 4120 7352 4126 7364
rect 5261 7361 5273 7364
rect 5307 7392 5319 7395
rect 5994 7392 6000 7404
rect 5307 7364 6000 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6273 7395 6331 7401
rect 6273 7361 6285 7395
rect 6319 7392 6331 7395
rect 6362 7392 6368 7404
rect 6319 7364 6368 7392
rect 6319 7361 6331 7364
rect 6273 7355 6331 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 8294 7392 8300 7404
rect 6871 7364 8300 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 9214 7392 9220 7404
rect 8864 7364 9220 7392
rect 8864 7333 8892 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10560 7364 10609 7392
rect 10560 7352 10566 7364
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 12158 7352 12164 7404
rect 12216 7392 12222 7404
rect 14277 7395 14335 7401
rect 12216 7364 13814 7392
rect 12216 7352 12222 7364
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3200 7296 3433 7324
rect 3200 7284 3206 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4525 7327 4583 7333
rect 4525 7324 4537 7327
rect 4019 7296 4537 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4525 7293 4537 7296
rect 4571 7324 4583 7327
rect 5077 7327 5135 7333
rect 5077 7324 5089 7327
rect 4571 7296 5089 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 5077 7293 5089 7296
rect 5123 7293 5135 7327
rect 8113 7327 8171 7333
rect 8113 7324 8125 7327
rect 5077 7287 5135 7293
rect 6012 7296 8125 7324
rect 2474 7259 2532 7265
rect 2474 7256 2486 7259
rect 2240 7228 2486 7256
rect 2240 7200 2268 7228
rect 2474 7225 2486 7228
rect 2520 7225 2532 7259
rect 2474 7219 2532 7225
rect 5350 7216 5356 7268
rect 5408 7256 5414 7268
rect 5902 7256 5908 7268
rect 5408 7228 5453 7256
rect 5863 7228 5908 7256
rect 5408 7216 5414 7228
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 2133 7191 2191 7197
rect 2133 7188 2145 7191
rect 1811 7160 2145 7188
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 2133 7157 2145 7160
rect 2179 7188 2191 7191
rect 2222 7188 2228 7200
rect 2179 7160 2228 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 6012 7188 6040 7296
rect 8113 7293 8125 7296
rect 8159 7324 8171 7327
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8159 7296 8861 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 9030 7324 9036 7336
rect 8991 7296 9036 7324
rect 8849 7287 8907 7293
rect 9030 7284 9036 7296
rect 9088 7324 9094 7336
rect 11606 7324 11612 7336
rect 9088 7296 11612 7324
rect 9088 7284 9094 7296
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 12360 7296 12541 7324
rect 6641 7259 6699 7265
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 7187 7259 7245 7265
rect 7187 7256 7199 7259
rect 6687 7228 7199 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 7187 7225 7199 7228
rect 7233 7256 7245 7259
rect 7282 7256 7288 7268
rect 7233 7228 7288 7256
rect 7233 7225 7245 7228
rect 7187 7219 7245 7225
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 8478 7256 8484 7268
rect 8391 7228 8484 7256
rect 8478 7216 8484 7228
rect 8536 7256 8542 7268
rect 9122 7256 9128 7268
rect 8536 7228 9128 7256
rect 8536 7216 8542 7228
rect 9122 7216 9128 7228
rect 9180 7216 9186 7268
rect 10505 7259 10563 7265
rect 10505 7225 10517 7259
rect 10551 7256 10563 7259
rect 10959 7259 11017 7265
rect 10959 7256 10971 7259
rect 10551 7228 10971 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 10959 7225 10971 7228
rect 11005 7256 11017 7259
rect 11005 7228 11192 7256
rect 11005 7225 11017 7228
rect 10959 7219 11017 7225
rect 11164 7200 11192 7228
rect 4028 7160 6040 7188
rect 4028 7148 4034 7160
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 8168 7160 8677 7188
rect 8168 7148 8174 7160
rect 8665 7157 8677 7160
rect 8711 7157 8723 7191
rect 8665 7151 8723 7157
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11204 7160 11805 7188
rect 11204 7148 11210 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 11793 7151 11851 7157
rect 12158 7148 12164 7160
rect 12216 7188 12222 7200
rect 12360 7188 12388 7296
rect 12529 7293 12541 7296
rect 12575 7293 12587 7327
rect 13786 7324 13814 7364
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 14323 7364 14964 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 13786 7296 14657 7324
rect 12529 7287 12587 7293
rect 14645 7293 14657 7296
rect 14691 7324 14703 7327
rect 14734 7324 14740 7336
rect 14691 7296 14740 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 14936 7333 14964 7364
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15856 7324 15884 7432
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 20530 7420 20536 7472
rect 20588 7460 20594 7472
rect 22373 7463 22431 7469
rect 22373 7460 22385 7463
rect 20588 7432 22385 7460
rect 20588 7420 20594 7432
rect 22373 7429 22385 7432
rect 22419 7460 22431 7463
rect 22738 7460 22744 7472
rect 22419 7432 22744 7460
rect 22419 7429 22431 7432
rect 22373 7423 22431 7429
rect 22738 7420 22744 7432
rect 22796 7420 22802 7472
rect 27154 7420 27160 7472
rect 27212 7460 27218 7472
rect 27939 7463 27997 7469
rect 27939 7460 27951 7463
rect 27212 7432 27951 7460
rect 27212 7420 27218 7432
rect 27939 7429 27951 7432
rect 27985 7429 27997 7463
rect 27939 7423 27997 7429
rect 28902 7420 28908 7472
rect 28960 7460 28966 7472
rect 30653 7463 30711 7469
rect 30653 7460 30665 7463
rect 28960 7432 30665 7460
rect 28960 7420 28966 7432
rect 30653 7429 30665 7432
rect 30699 7429 30711 7463
rect 30653 7423 30711 7429
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7392 16083 7395
rect 16482 7392 16488 7404
rect 16071 7364 16488 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16666 7392 16672 7404
rect 16627 7364 16672 7392
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7392 18107 7395
rect 18138 7392 18144 7404
rect 18095 7364 18144 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 19944 7364 19993 7392
rect 19944 7352 19950 7364
rect 19981 7361 19993 7364
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 22094 7392 22100 7404
rect 21867 7364 22100 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 22094 7352 22100 7364
rect 22152 7352 22158 7404
rect 23750 7392 23756 7404
rect 23711 7364 23756 7392
rect 23750 7352 23756 7364
rect 23808 7352 23814 7404
rect 24118 7392 24124 7404
rect 24079 7364 24124 7392
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 25590 7352 25596 7404
rect 25648 7392 25654 7404
rect 26050 7392 26056 7404
rect 25648 7364 26056 7392
rect 25648 7352 25654 7364
rect 26050 7352 26056 7364
rect 26108 7352 26114 7404
rect 26326 7352 26332 7404
rect 26384 7392 26390 7404
rect 26786 7392 26792 7404
rect 26384 7364 26792 7392
rect 26384 7352 26390 7364
rect 26786 7352 26792 7364
rect 26844 7392 26850 7404
rect 27249 7395 27307 7401
rect 27249 7392 27261 7395
rect 26844 7364 27261 7392
rect 26844 7352 26850 7364
rect 27249 7361 27261 7364
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 29178 7352 29184 7404
rect 29236 7392 29242 7404
rect 29365 7395 29423 7401
rect 29365 7392 29377 7395
rect 29236 7364 29377 7392
rect 29236 7352 29242 7364
rect 29365 7361 29377 7364
rect 29411 7361 29423 7395
rect 29365 7355 29423 7361
rect 14967 7296 15884 7324
rect 25317 7327 25375 7333
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 25317 7293 25329 7327
rect 25363 7324 25375 7327
rect 25406 7324 25412 7336
rect 25363 7296 25412 7324
rect 25363 7293 25375 7296
rect 25317 7287 25375 7293
rect 25406 7284 25412 7296
rect 25464 7324 25470 7336
rect 27868 7327 27926 7333
rect 25464 7296 26878 7324
rect 25464 7284 25470 7296
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7256 15163 7259
rect 16022 7256 16028 7268
rect 15151 7228 16028 7256
rect 15151 7225 15163 7228
rect 15105 7219 15163 7225
rect 16022 7216 16028 7228
rect 16080 7216 16086 7268
rect 16114 7216 16120 7268
rect 16172 7256 16178 7268
rect 17862 7256 17868 7268
rect 16172 7228 16217 7256
rect 17775 7228 17868 7256
rect 16172 7216 16178 7228
rect 17862 7216 17868 7228
rect 17920 7256 17926 7268
rect 18411 7259 18469 7265
rect 18411 7256 18423 7259
rect 17920 7228 18423 7256
rect 17920 7216 17926 7228
rect 18411 7225 18423 7228
rect 18457 7256 18469 7259
rect 19242 7256 19248 7268
rect 18457 7228 19248 7256
rect 18457 7225 18469 7228
rect 18411 7219 18469 7225
rect 19242 7216 19248 7228
rect 19300 7256 19306 7268
rect 20302 7259 20360 7265
rect 19300 7216 19334 7256
rect 20302 7225 20314 7259
rect 20348 7225 20360 7259
rect 20302 7219 20360 7225
rect 12894 7188 12900 7200
rect 12216 7160 12388 7188
rect 12855 7160 12900 7188
rect 12216 7148 12222 7160
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16132 7188 16160 7216
rect 19306 7200 19334 7216
rect 17126 7188 17132 7200
rect 15887 7160 16160 7188
rect 17087 7160 17132 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 19306 7160 19340 7200
rect 19334 7148 19340 7160
rect 19392 7188 19398 7200
rect 19797 7191 19855 7197
rect 19797 7188 19809 7191
rect 19392 7160 19809 7188
rect 19392 7148 19398 7160
rect 19797 7157 19809 7160
rect 19843 7188 19855 7191
rect 20317 7188 20345 7219
rect 21910 7216 21916 7268
rect 21968 7256 21974 7268
rect 22830 7256 22836 7268
rect 21968 7228 22013 7256
rect 22743 7228 22836 7256
rect 21968 7216 21974 7228
rect 22830 7216 22836 7228
rect 22888 7256 22894 7268
rect 23750 7256 23756 7268
rect 22888 7228 23756 7256
rect 22888 7216 22894 7228
rect 23750 7216 23756 7228
rect 23808 7216 23814 7268
rect 23845 7259 23903 7265
rect 23845 7225 23857 7259
rect 23891 7225 23903 7259
rect 26326 7256 26332 7268
rect 23845 7219 23903 7225
rect 25884 7228 26332 7256
rect 22554 7188 22560 7200
rect 19843 7160 22560 7188
rect 19843 7157 19855 7160
rect 19797 7151 19855 7157
rect 22554 7148 22560 7160
rect 22612 7148 22618 7200
rect 23198 7148 23204 7200
rect 23256 7188 23262 7200
rect 23385 7191 23443 7197
rect 23385 7188 23397 7191
rect 23256 7160 23397 7188
rect 23256 7148 23262 7160
rect 23385 7157 23397 7160
rect 23431 7188 23443 7191
rect 23860 7188 23888 7219
rect 25884 7200 25912 7228
rect 26326 7216 26332 7228
rect 26384 7265 26390 7268
rect 26384 7259 26432 7265
rect 26384 7225 26386 7259
rect 26420 7225 26432 7259
rect 26850 7256 26878 7296
rect 27868 7293 27880 7327
rect 27914 7324 27926 7327
rect 28258 7324 28264 7336
rect 27914 7296 28264 7324
rect 27914 7293 27926 7296
rect 27868 7287 27926 7293
rect 28258 7284 28264 7296
rect 28316 7284 28322 7336
rect 30668 7324 30696 7423
rect 34606 7420 34612 7472
rect 34664 7460 34670 7472
rect 35989 7463 36047 7469
rect 35989 7460 36001 7463
rect 34664 7432 36001 7460
rect 34664 7420 34670 7432
rect 35989 7429 36001 7432
rect 36035 7429 36047 7463
rect 35989 7423 36047 7429
rect 31386 7392 31392 7404
rect 31347 7364 31392 7392
rect 31386 7352 31392 7364
rect 31444 7352 31450 7404
rect 33321 7395 33379 7401
rect 33321 7361 33333 7395
rect 33367 7392 33379 7395
rect 33502 7392 33508 7404
rect 33367 7364 33508 7392
rect 33367 7361 33379 7364
rect 33321 7355 33379 7361
rect 33502 7352 33508 7364
rect 33560 7352 33566 7404
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7392 35035 7395
rect 35894 7392 35900 7404
rect 35023 7364 35900 7392
rect 35023 7361 35035 7364
rect 34977 7355 35035 7361
rect 35894 7352 35900 7364
rect 35952 7352 35958 7404
rect 30837 7327 30895 7333
rect 30837 7324 30849 7327
rect 30668 7296 30849 7324
rect 30837 7293 30849 7296
rect 30883 7293 30895 7327
rect 31294 7324 31300 7336
rect 31255 7296 31300 7324
rect 30837 7287 30895 7293
rect 31294 7284 31300 7296
rect 31352 7284 31358 7336
rect 28442 7256 28448 7268
rect 26850 7228 28448 7256
rect 26384 7219 26432 7225
rect 26384 7216 26390 7219
rect 28442 7216 28448 7228
rect 28500 7216 28506 7268
rect 29454 7216 29460 7268
rect 29512 7256 29518 7268
rect 30006 7256 30012 7268
rect 29512 7228 29557 7256
rect 29967 7228 30012 7256
rect 29512 7216 29518 7228
rect 30006 7216 30012 7228
rect 30064 7216 30070 7268
rect 33042 7216 33048 7268
rect 33100 7256 33106 7268
rect 33413 7259 33471 7265
rect 33100 7228 33180 7256
rect 33100 7216 33106 7228
rect 25866 7188 25872 7200
rect 23431 7160 23888 7188
rect 25827 7160 25872 7188
rect 23431 7157 23443 7160
rect 23385 7151 23443 7157
rect 25866 7148 25872 7160
rect 25924 7148 25930 7200
rect 29089 7191 29147 7197
rect 29089 7157 29101 7191
rect 29135 7188 29147 7191
rect 29472 7188 29500 7216
rect 30282 7188 30288 7200
rect 29135 7160 29500 7188
rect 30243 7160 30288 7188
rect 29135 7157 29147 7160
rect 29089 7151 29147 7157
rect 30282 7148 30288 7160
rect 30340 7188 30346 7200
rect 30466 7188 30472 7200
rect 30340 7160 30472 7188
rect 30340 7148 30346 7160
rect 30466 7148 30472 7160
rect 30524 7148 30530 7200
rect 32217 7191 32275 7197
rect 32217 7157 32229 7191
rect 32263 7188 32275 7191
rect 32490 7188 32496 7200
rect 32263 7160 32496 7188
rect 32263 7157 32275 7160
rect 32217 7151 32275 7157
rect 32490 7148 32496 7160
rect 32548 7148 32554 7200
rect 33152 7188 33180 7228
rect 33413 7225 33425 7259
rect 33459 7225 33471 7259
rect 33413 7219 33471 7225
rect 33965 7259 34023 7265
rect 33965 7225 33977 7259
rect 34011 7256 34023 7259
rect 34974 7256 34980 7268
rect 34011 7228 34980 7256
rect 34011 7225 34023 7228
rect 33965 7219 34023 7225
rect 33428 7188 33456 7219
rect 34974 7216 34980 7228
rect 35032 7216 35038 7268
rect 35069 7259 35127 7265
rect 35069 7225 35081 7259
rect 35115 7225 35127 7259
rect 35618 7256 35624 7268
rect 35579 7228 35624 7256
rect 35069 7219 35127 7225
rect 34698 7188 34704 7200
rect 33152 7160 33456 7188
rect 34659 7160 34704 7188
rect 34698 7148 34704 7160
rect 34756 7148 34762 7200
rect 34790 7148 34796 7200
rect 34848 7188 34854 7200
rect 35084 7188 35112 7219
rect 35618 7216 35624 7228
rect 35676 7216 35682 7268
rect 36004 7256 36032 7423
rect 36354 7352 36360 7404
rect 36412 7392 36418 7404
rect 36541 7395 36599 7401
rect 36541 7392 36553 7395
rect 36412 7364 36553 7392
rect 36412 7352 36418 7364
rect 36541 7361 36553 7364
rect 36587 7361 36599 7395
rect 36814 7392 36820 7404
rect 36775 7364 36820 7392
rect 36541 7355 36599 7361
rect 36814 7352 36820 7364
rect 36872 7352 36878 7404
rect 36633 7259 36691 7265
rect 36633 7256 36645 7259
rect 36004 7228 36645 7256
rect 36633 7225 36645 7228
rect 36679 7225 36691 7259
rect 36633 7219 36691 7225
rect 34848 7160 35112 7188
rect 34848 7148 34854 7160
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 1854 6984 1860 6996
rect 1719 6956 1860 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 1854 6944 1860 6956
rect 1912 6944 1918 6996
rect 2130 6984 2136 6996
rect 2091 6956 2136 6984
rect 2130 6944 2136 6956
rect 2188 6944 2194 6996
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2280 6956 2589 6984
rect 2280 6944 2286 6956
rect 2561 6925 2589 6956
rect 2866 6944 2872 6996
rect 2924 6984 2930 6996
rect 3145 6987 3203 6993
rect 3145 6984 3157 6987
rect 2924 6956 3157 6984
rect 2924 6944 2930 6956
rect 3145 6953 3157 6956
rect 3191 6953 3203 6987
rect 4338 6984 4344 6996
rect 4299 6956 4344 6984
rect 3145 6947 3203 6953
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 5629 6987 5687 6993
rect 5629 6984 5641 6987
rect 5408 6956 5641 6984
rect 5408 6944 5414 6956
rect 5629 6953 5641 6956
rect 5675 6953 5687 6987
rect 5994 6984 6000 6996
rect 5955 6956 6000 6984
rect 5629 6947 5687 6953
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 8294 6984 8300 6996
rect 7699 6956 8300 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 10597 6987 10655 6993
rect 10597 6984 10609 6987
rect 10560 6956 10609 6984
rect 10560 6944 10566 6956
rect 10597 6953 10609 6956
rect 10643 6953 10655 6987
rect 11974 6984 11980 6996
rect 11935 6956 11980 6984
rect 10597 6947 10655 6953
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 14461 6987 14519 6993
rect 14461 6953 14473 6987
rect 14507 6984 14519 6987
rect 14734 6984 14740 6996
rect 14507 6956 14740 6984
rect 14507 6953 14519 6956
rect 14461 6947 14519 6953
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 15010 6944 15016 6996
rect 15068 6984 15074 6996
rect 15749 6987 15807 6993
rect 15749 6984 15761 6987
rect 15068 6956 15761 6984
rect 15068 6944 15074 6956
rect 15749 6953 15761 6956
rect 15795 6953 15807 6987
rect 15749 6947 15807 6953
rect 16301 6987 16359 6993
rect 16301 6953 16313 6987
rect 16347 6984 16359 6987
rect 16390 6984 16396 6996
rect 16347 6956 16396 6984
rect 16347 6953 16359 6956
rect 16301 6947 16359 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18601 6987 18659 6993
rect 18601 6953 18613 6987
rect 18647 6984 18659 6987
rect 18690 6984 18696 6996
rect 18647 6956 18696 6984
rect 18647 6953 18659 6956
rect 18601 6947 18659 6953
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 19886 6944 19892 6996
rect 19944 6984 19950 6996
rect 19981 6987 20039 6993
rect 19981 6984 19993 6987
rect 19944 6956 19993 6984
rect 19944 6944 19950 6956
rect 19981 6953 19993 6956
rect 20027 6953 20039 6987
rect 19981 6947 20039 6953
rect 22554 6944 22560 6996
rect 22612 6984 22618 6996
rect 22649 6987 22707 6993
rect 22649 6984 22661 6987
rect 22612 6956 22661 6984
rect 22612 6944 22618 6956
rect 22649 6953 22661 6956
rect 22695 6953 22707 6987
rect 23198 6984 23204 6996
rect 23159 6956 23204 6984
rect 22649 6947 22707 6953
rect 23198 6944 23204 6956
rect 23256 6944 23262 6996
rect 23750 6944 23756 6996
rect 23808 6984 23814 6996
rect 24949 6987 25007 6993
rect 24949 6984 24961 6987
rect 23808 6956 24961 6984
rect 23808 6944 23814 6956
rect 24949 6953 24961 6956
rect 24995 6953 25007 6987
rect 26050 6984 26056 6996
rect 26011 6956 26056 6984
rect 24949 6947 25007 6953
rect 26050 6944 26056 6956
rect 26108 6944 26114 6996
rect 26927 6987 26985 6993
rect 26927 6953 26939 6987
rect 26973 6984 26985 6987
rect 27522 6984 27528 6996
rect 26973 6956 27528 6984
rect 26973 6953 26985 6956
rect 26927 6947 26985 6953
rect 27522 6944 27528 6956
rect 27580 6944 27586 6996
rect 27709 6987 27767 6993
rect 27709 6953 27721 6987
rect 27755 6984 27767 6987
rect 28534 6984 28540 6996
rect 27755 6956 28540 6984
rect 27755 6953 27767 6956
rect 27709 6947 27767 6953
rect 28534 6944 28540 6956
rect 28592 6944 28598 6996
rect 28626 6944 28632 6996
rect 28684 6984 28690 6996
rect 28721 6987 28779 6993
rect 28721 6984 28733 6987
rect 28684 6956 28733 6984
rect 28684 6944 28690 6956
rect 28721 6953 28733 6956
rect 28767 6953 28779 6987
rect 28721 6947 28779 6953
rect 29178 6944 29184 6996
rect 29236 6984 29242 6996
rect 29273 6987 29331 6993
rect 29273 6984 29285 6987
rect 29236 6956 29285 6984
rect 29236 6944 29242 6956
rect 29273 6953 29285 6956
rect 29319 6953 29331 6987
rect 29273 6947 29331 6953
rect 29454 6944 29460 6996
rect 29512 6984 29518 6996
rect 30469 6987 30527 6993
rect 30469 6984 30481 6987
rect 29512 6956 30481 6984
rect 29512 6944 29518 6956
rect 30469 6953 30481 6956
rect 30515 6953 30527 6987
rect 30469 6947 30527 6953
rect 30650 6944 30656 6996
rect 30708 6984 30714 6996
rect 31113 6987 31171 6993
rect 31113 6984 31125 6987
rect 30708 6956 31125 6984
rect 30708 6944 30714 6956
rect 31113 6953 31125 6956
rect 31159 6984 31171 6987
rect 31570 6984 31576 6996
rect 31159 6956 31576 6984
rect 31159 6953 31171 6956
rect 31113 6947 31171 6953
rect 31570 6944 31576 6956
rect 31628 6944 31634 6996
rect 34146 6984 34152 6996
rect 34107 6956 34152 6984
rect 34146 6944 34152 6956
rect 34204 6944 34210 6996
rect 34698 6944 34704 6996
rect 34756 6984 34762 6996
rect 36449 6987 36507 6993
rect 36449 6984 36461 6987
rect 34756 6956 36461 6984
rect 34756 6944 34762 6956
rect 36449 6953 36461 6956
rect 36495 6953 36507 6987
rect 36449 6947 36507 6953
rect 2546 6919 2604 6925
rect 2546 6885 2558 6919
rect 2592 6885 2604 6919
rect 2546 6879 2604 6885
rect 3050 6876 3056 6928
rect 3108 6916 3114 6928
rect 3421 6919 3479 6925
rect 3421 6916 3433 6919
rect 3108 6888 3433 6916
rect 3108 6876 3114 6888
rect 3421 6885 3433 6888
rect 3467 6885 3479 6919
rect 3421 6879 3479 6885
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 4801 6919 4859 6925
rect 4801 6916 4813 6919
rect 4764 6888 4813 6916
rect 4764 6876 4770 6888
rect 4801 6885 4813 6888
rect 4847 6885 4859 6919
rect 6362 6916 6368 6928
rect 6323 6888 6368 6916
rect 4801 6879 4859 6885
rect 6362 6876 6368 6888
rect 6420 6876 6426 6928
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 7837 6919 7895 6925
rect 7837 6916 7849 6919
rect 7524 6888 7849 6916
rect 7524 6876 7530 6888
rect 7837 6885 7849 6888
rect 7883 6885 7895 6919
rect 7837 6879 7895 6885
rect 7929 6919 7987 6925
rect 7929 6885 7941 6919
rect 7975 6916 7987 6919
rect 8018 6916 8024 6928
rect 7975 6888 8024 6916
rect 7975 6885 7987 6888
rect 7929 6879 7987 6885
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 9815 6919 9873 6925
rect 9815 6916 9827 6919
rect 8536 6888 9827 6916
rect 8536 6876 8542 6888
rect 9815 6885 9827 6888
rect 9861 6885 9873 6919
rect 9815 6879 9873 6885
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 11378 6919 11436 6925
rect 11378 6916 11390 6919
rect 11204 6888 11390 6916
rect 11204 6876 11210 6888
rect 11378 6885 11390 6888
rect 11424 6885 11436 6919
rect 11378 6879 11436 6885
rect 12894 6876 12900 6928
rect 12952 6916 12958 6928
rect 12989 6919 13047 6925
rect 12989 6916 13001 6919
rect 12952 6888 13001 6916
rect 12952 6876 12958 6888
rect 12989 6885 13001 6888
rect 13035 6885 13047 6919
rect 13538 6916 13544 6928
rect 13499 6888 13544 6916
rect 12989 6879 13047 6885
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 16847 6919 16905 6925
rect 16847 6885 16859 6919
rect 16893 6916 16905 6919
rect 16942 6916 16948 6928
rect 16893 6888 16948 6916
rect 16893 6885 16905 6888
rect 16847 6879 16905 6885
rect 16942 6876 16948 6888
rect 17000 6916 17006 6928
rect 17862 6916 17868 6928
rect 17000 6888 17868 6916
rect 17000 6876 17006 6888
rect 17862 6876 17868 6888
rect 17920 6876 17926 6928
rect 18874 6916 18880 6928
rect 18835 6888 18880 6916
rect 18874 6876 18880 6888
rect 18932 6876 18938 6928
rect 18966 6876 18972 6928
rect 19024 6916 19030 6928
rect 20349 6919 20407 6925
rect 20349 6916 20361 6919
rect 19024 6888 20361 6916
rect 19024 6876 19030 6888
rect 20349 6885 20361 6888
rect 20395 6885 20407 6919
rect 20349 6879 20407 6885
rect 21453 6919 21511 6925
rect 21453 6885 21465 6919
rect 21499 6916 21511 6919
rect 22462 6916 22468 6928
rect 21499 6888 22468 6916
rect 21499 6885 21511 6888
rect 21453 6879 21511 6885
rect 22462 6876 22468 6888
rect 22520 6876 22526 6928
rect 24282 6919 24340 6925
rect 24282 6885 24294 6919
rect 24328 6916 24340 6919
rect 24394 6916 24400 6928
rect 24328 6888 24400 6916
rect 24328 6885 24340 6888
rect 24282 6879 24340 6885
rect 24394 6876 24400 6888
rect 24452 6876 24458 6928
rect 28163 6919 28221 6925
rect 28163 6885 28175 6919
rect 28209 6916 28221 6919
rect 28810 6916 28816 6928
rect 28209 6888 28816 6916
rect 28209 6885 28221 6888
rect 28163 6879 28221 6885
rect 28810 6876 28816 6888
rect 28868 6916 28874 6928
rect 29911 6919 29969 6925
rect 29911 6916 29923 6919
rect 28868 6888 29923 6916
rect 28868 6876 28874 6888
rect 29911 6885 29923 6888
rect 29957 6885 29969 6919
rect 35434 6916 35440 6928
rect 35395 6888 35440 6916
rect 29911 6879 29969 6885
rect 35434 6876 35440 6888
rect 35492 6876 35498 6928
rect 35891 6919 35949 6925
rect 35891 6885 35903 6919
rect 35937 6916 35949 6919
rect 35986 6916 35992 6928
rect 35937 6888 35992 6916
rect 35937 6885 35949 6888
rect 35891 6879 35949 6885
rect 35986 6876 35992 6888
rect 36044 6876 36050 6928
rect 36354 6876 36360 6928
rect 36412 6916 36418 6928
rect 36725 6919 36783 6925
rect 36725 6916 36737 6919
rect 36412 6888 36737 6916
rect 36412 6876 36418 6888
rect 36725 6885 36737 6888
rect 36771 6885 36783 6919
rect 36725 6879 36783 6885
rect 2038 6808 2044 6860
rect 2096 6848 2102 6860
rect 2225 6851 2283 6857
rect 2225 6848 2237 6851
rect 2096 6820 2237 6848
rect 2096 6808 2102 6820
rect 2225 6817 2237 6820
rect 2271 6817 2283 6851
rect 2225 6811 2283 6817
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 5902 6848 5908 6860
rect 5399 6820 5908 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9712 6851 9770 6857
rect 9712 6848 9724 6851
rect 9640 6820 9724 6848
rect 9640 6808 9646 6820
rect 9712 6817 9724 6820
rect 9758 6817 9770 6851
rect 11054 6848 11060 6860
rect 11015 6820 11060 6848
rect 9712 6811 9770 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 15286 6848 15292 6860
rect 15199 6820 15292 6848
rect 15286 6808 15292 6820
rect 15344 6848 15350 6860
rect 15470 6848 15476 6860
rect 15344 6820 15476 6848
rect 15344 6808 15350 6820
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 16485 6851 16543 6857
rect 16485 6817 16497 6851
rect 16531 6848 16543 6851
rect 16574 6848 16580 6860
rect 16531 6820 16580 6848
rect 16531 6817 16543 6820
rect 16485 6811 16543 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 20254 6808 20260 6860
rect 20312 6848 20318 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20312 6820 20913 6848
rect 20312 6808 20318 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 21085 6851 21143 6857
rect 21085 6817 21097 6851
rect 21131 6817 21143 6851
rect 21085 6811 21143 6817
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5442 6780 5448 6792
rect 4755 6752 5448 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 6270 6780 6276 6792
rect 6231 6752 6276 6780
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 6564 6712 6592 6740
rect 8128 6712 8156 6743
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12492 6752 12909 6780
rect 12492 6740 12498 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 13354 6780 13360 6792
rect 12897 6743 12955 6749
rect 13004 6752 13360 6780
rect 8202 6712 8208 6724
rect 6564 6684 8208 6712
rect 8202 6672 8208 6684
rect 8260 6712 8266 6724
rect 9125 6715 9183 6721
rect 9125 6712 9137 6715
rect 8260 6684 9137 6712
rect 8260 6672 8266 6684
rect 9125 6681 9137 6684
rect 9171 6681 9183 6715
rect 10226 6712 10232 6724
rect 10139 6684 10232 6712
rect 9125 6675 9183 6681
rect 10226 6672 10232 6684
rect 10284 6712 10290 6724
rect 13004 6712 13032 6752
rect 13354 6740 13360 6752
rect 13412 6780 13418 6792
rect 15378 6780 15384 6792
rect 13412 6752 15384 6780
rect 13412 6740 13418 6752
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 18782 6780 18788 6792
rect 18743 6752 18788 6780
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 21100 6780 21128 6811
rect 22738 6808 22744 6860
rect 22796 6848 22802 6860
rect 23477 6851 23535 6857
rect 23477 6848 23489 6851
rect 22796 6820 23489 6848
rect 22796 6808 22802 6820
rect 23477 6817 23489 6820
rect 23523 6817 23535 6851
rect 23477 6811 23535 6817
rect 26602 6808 26608 6860
rect 26660 6848 26666 6860
rect 26824 6851 26882 6857
rect 26824 6848 26836 6851
rect 26660 6820 26836 6848
rect 26660 6808 26666 6820
rect 26824 6817 26836 6820
rect 26870 6817 26882 6851
rect 32122 6848 32128 6860
rect 32083 6820 32128 6848
rect 26824 6811 26882 6817
rect 32122 6808 32128 6820
rect 32180 6808 32186 6860
rect 32674 6848 32680 6860
rect 32635 6820 32680 6848
rect 32674 6808 32680 6820
rect 32732 6808 32738 6860
rect 34606 6808 34612 6860
rect 34664 6848 34670 6860
rect 34701 6851 34759 6857
rect 34701 6848 34713 6851
rect 34664 6820 34713 6848
rect 34664 6808 34670 6820
rect 34701 6817 34713 6820
rect 34747 6817 34759 6851
rect 34701 6811 34759 6817
rect 20772 6752 21128 6780
rect 22281 6783 22339 6789
rect 20772 6740 20778 6752
rect 22281 6749 22293 6783
rect 22327 6780 22339 6783
rect 22370 6780 22376 6792
rect 22327 6752 22376 6780
rect 22327 6749 22339 6752
rect 22281 6743 22339 6749
rect 22370 6740 22376 6752
rect 22428 6740 22434 6792
rect 24029 6783 24087 6789
rect 24029 6780 24041 6783
rect 23860 6752 24041 6780
rect 10284 6684 13032 6712
rect 10284 6672 10290 6684
rect 13630 6672 13636 6724
rect 13688 6712 13694 6724
rect 15473 6715 15531 6721
rect 15473 6712 15485 6715
rect 13688 6684 15485 6712
rect 13688 6672 13694 6684
rect 15473 6681 15485 6684
rect 15519 6681 15531 6715
rect 15473 6675 15531 6681
rect 23860 6656 23888 6752
rect 24029 6749 24041 6752
rect 24075 6749 24087 6783
rect 27798 6780 27804 6792
rect 27759 6752 27804 6780
rect 24029 6743 24087 6749
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 29546 6780 29552 6792
rect 29507 6752 29552 6780
rect 29546 6740 29552 6752
rect 29604 6740 29610 6792
rect 30837 6783 30895 6789
rect 30837 6749 30849 6783
rect 30883 6780 30895 6783
rect 31294 6780 31300 6792
rect 30883 6752 31300 6780
rect 30883 6749 30895 6752
rect 30837 6743 30895 6749
rect 31294 6740 31300 6752
rect 31352 6780 31358 6792
rect 31573 6783 31631 6789
rect 31573 6780 31585 6783
rect 31352 6752 31585 6780
rect 31352 6740 31358 6752
rect 31573 6749 31585 6752
rect 31619 6780 31631 6783
rect 32692 6780 32720 6808
rect 31619 6752 32720 6780
rect 32861 6783 32919 6789
rect 31619 6749 31631 6752
rect 31573 6743 31631 6749
rect 32861 6749 32873 6783
rect 32907 6780 32919 6783
rect 33778 6780 33784 6792
rect 32907 6752 33784 6780
rect 32907 6749 32919 6752
rect 32861 6743 32919 6749
rect 33778 6740 33784 6752
rect 33836 6740 33842 6792
rect 35250 6740 35256 6792
rect 35308 6780 35314 6792
rect 35529 6783 35587 6789
rect 35529 6780 35541 6783
rect 35308 6752 35541 6780
rect 35308 6740 35314 6752
rect 35529 6749 35541 6752
rect 35575 6749 35587 6783
rect 35529 6743 35587 6749
rect 106 6604 112 6656
rect 164 6644 170 6656
rect 3510 6644 3516 6656
rect 164 6616 3516 6644
rect 164 6604 170 6616
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 7282 6644 7288 6656
rect 7243 6616 7288 6644
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 8849 6647 8907 6653
rect 8849 6613 8861 6647
rect 8895 6644 8907 6647
rect 9030 6644 9036 6656
rect 8895 6616 9036 6644
rect 8895 6613 8907 6616
rect 8849 6607 8907 6613
rect 9030 6604 9036 6616
rect 9088 6644 9094 6656
rect 9490 6644 9496 6656
rect 9088 6616 9496 6644
rect 9088 6604 9094 6616
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 17126 6604 17132 6656
rect 17184 6644 17190 6656
rect 17405 6647 17463 6653
rect 17405 6644 17417 6647
rect 17184 6616 17417 6644
rect 17184 6604 17190 6616
rect 17405 6613 17417 6616
rect 17451 6644 17463 6647
rect 17862 6644 17868 6656
rect 17451 6616 17868 6644
rect 17451 6613 17463 6616
rect 17405 6607 17463 6613
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 20162 6604 20168 6656
rect 20220 6644 20226 6656
rect 21913 6647 21971 6653
rect 21913 6644 21925 6647
rect 20220 6616 21925 6644
rect 20220 6604 20226 6616
rect 21913 6613 21925 6616
rect 21959 6644 21971 6647
rect 22278 6644 22284 6656
rect 21959 6616 22284 6644
rect 21959 6613 21971 6616
rect 21913 6607 21971 6613
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 23842 6644 23848 6656
rect 23803 6616 23848 6644
rect 23842 6604 23848 6616
rect 23900 6604 23906 6656
rect 27341 6647 27399 6653
rect 27341 6613 27353 6647
rect 27387 6644 27399 6647
rect 27522 6644 27528 6656
rect 27387 6616 27528 6644
rect 27387 6613 27399 6616
rect 27341 6607 27399 6613
rect 27522 6604 27528 6616
rect 27580 6604 27586 6656
rect 33318 6644 33324 6656
rect 33279 6616 33324 6644
rect 33318 6604 33324 6616
rect 33376 6604 33382 6656
rect 34790 6604 34796 6656
rect 34848 6644 34854 6656
rect 34977 6647 35035 6653
rect 34977 6644 34989 6647
rect 34848 6616 34989 6644
rect 34848 6604 34854 6616
rect 34977 6613 34989 6616
rect 35023 6613 35035 6647
rect 34977 6607 35035 6613
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 3605 6443 3663 6449
rect 3605 6440 3617 6443
rect 2096 6412 3617 6440
rect 2096 6400 2102 6412
rect 3605 6409 3617 6412
rect 3651 6409 3663 6443
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 3605 6403 3663 6409
rect 4126 6412 4353 6440
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2130 6304 2136 6316
rect 2087 6276 2136 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 3856 6239 3914 6245
rect 3856 6205 3868 6239
rect 3902 6236 3914 6239
rect 4126 6236 4154 6412
rect 4341 6409 4353 6412
rect 4387 6440 4399 6443
rect 4890 6440 4896 6452
rect 4387 6412 4896 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6328 6412 6561 6440
rect 6328 6400 6334 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 9950 6440 9956 6452
rect 6549 6403 6607 6409
rect 7300 6412 9956 6440
rect 4614 6332 4620 6384
rect 4672 6372 4678 6384
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 4672 6344 6193 6372
rect 4672 6332 4678 6344
rect 6181 6341 6193 6344
rect 6227 6372 6239 6375
rect 6362 6372 6368 6384
rect 6227 6344 6368 6372
rect 6227 6341 6239 6344
rect 6181 6335 6239 6341
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 5258 6304 5264 6316
rect 5219 6276 5264 6304
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6546 6304 6552 6316
rect 5951 6276 6552 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 3902 6208 4154 6236
rect 3902 6205 3914 6208
rect 3856 6199 3914 6205
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 7300 6245 7328 6412
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10781 6443 10839 6449
rect 10781 6409 10793 6443
rect 10827 6440 10839 6443
rect 11054 6440 11060 6452
rect 10827 6412 11060 6440
rect 10827 6409 10839 6412
rect 10781 6403 10839 6409
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 12952 6412 13461 6440
rect 12952 6400 12958 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 15749 6443 15807 6449
rect 15749 6409 15761 6443
rect 15795 6440 15807 6443
rect 16574 6440 16580 6452
rect 15795 6412 16580 6440
rect 15795 6409 15807 6412
rect 15749 6403 15807 6409
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 17129 6443 17187 6449
rect 17129 6409 17141 6443
rect 17175 6440 17187 6443
rect 18509 6443 18567 6449
rect 18509 6440 18521 6443
rect 17175 6412 18521 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 18509 6409 18521 6412
rect 18555 6440 18567 6443
rect 18874 6440 18880 6452
rect 18555 6412 18880 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19794 6440 19800 6452
rect 19755 6412 19800 6440
rect 19794 6400 19800 6412
rect 19852 6440 19858 6452
rect 19852 6412 20392 6440
rect 19852 6400 19858 6412
rect 11517 6375 11575 6381
rect 11517 6341 11529 6375
rect 11563 6372 11575 6375
rect 13906 6372 13912 6384
rect 11563 6344 13912 6372
rect 11563 6341 11575 6344
rect 11517 6335 11575 6341
rect 8202 6304 8208 6316
rect 8163 6276 8208 6304
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 11532 6304 11560 6335
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 17497 6375 17555 6381
rect 17497 6341 17509 6375
rect 17543 6372 17555 6375
rect 18782 6372 18788 6384
rect 17543 6344 18788 6372
rect 17543 6341 17555 6344
rect 17497 6335 17555 6341
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 12526 6304 12532 6316
rect 9968 6276 11560 6304
rect 12487 6276 12532 6304
rect 6860 6239 6918 6245
rect 6860 6236 6872 6239
rect 6052 6208 6872 6236
rect 6052 6196 6058 6208
rect 6860 6205 6872 6208
rect 6906 6236 6918 6239
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6906 6208 7297 6236
rect 6906 6205 6918 6208
rect 6860 6199 6918 6205
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 9214 6236 9220 6248
rect 9127 6208 9220 6236
rect 7285 6199 7343 6205
rect 9214 6196 9220 6208
rect 9272 6236 9278 6248
rect 9968 6245 9996 6276
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 13538 6304 13544 6316
rect 13219 6276 13544 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6304 16267 6307
rect 16390 6304 16396 6316
rect 16255 6276 16396 6304
rect 16255 6273 16267 6276
rect 16209 6267 16267 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 20364 6313 20392 6412
rect 24394 6400 24400 6452
rect 24452 6440 24458 6452
rect 24765 6443 24823 6449
rect 24765 6440 24777 6443
rect 24452 6412 24777 6440
rect 24452 6400 24458 6412
rect 24765 6409 24777 6412
rect 24811 6440 24823 6443
rect 24949 6443 25007 6449
rect 24949 6440 24961 6443
rect 24811 6412 24961 6440
rect 24811 6409 24823 6412
rect 24765 6403 24823 6409
rect 24949 6409 24961 6412
rect 24995 6440 25007 6443
rect 25041 6443 25099 6449
rect 25041 6440 25053 6443
rect 24995 6412 25053 6440
rect 24995 6409 25007 6412
rect 24949 6403 25007 6409
rect 25041 6409 25053 6412
rect 25087 6409 25099 6443
rect 25041 6403 25099 6409
rect 26878 6400 26884 6452
rect 26936 6440 26942 6452
rect 28905 6443 28963 6449
rect 28905 6440 28917 6443
rect 26936 6412 28917 6440
rect 26936 6400 26942 6412
rect 28905 6409 28917 6412
rect 28951 6440 28963 6443
rect 28997 6443 29055 6449
rect 28997 6440 29009 6443
rect 28951 6412 29009 6440
rect 28951 6409 28963 6412
rect 28905 6403 28963 6409
rect 28997 6409 29009 6412
rect 29043 6440 29055 6443
rect 32306 6440 32312 6452
rect 29043 6412 32312 6440
rect 29043 6409 29055 6412
rect 28997 6403 29055 6409
rect 32306 6400 32312 6412
rect 32364 6400 32370 6452
rect 32585 6443 32643 6449
rect 32585 6409 32597 6443
rect 32631 6440 32643 6443
rect 32674 6440 32680 6452
rect 32631 6412 32680 6440
rect 32631 6409 32643 6412
rect 32585 6403 32643 6409
rect 32674 6400 32680 6412
rect 32732 6400 32738 6452
rect 34146 6400 34152 6452
rect 34204 6440 34210 6452
rect 34333 6443 34391 6449
rect 34333 6440 34345 6443
rect 34204 6412 34345 6440
rect 34204 6400 34210 6412
rect 34333 6409 34345 6412
rect 34379 6440 34391 6443
rect 35986 6440 35992 6452
rect 34379 6412 35992 6440
rect 34379 6409 34391 6412
rect 34333 6403 34391 6409
rect 35986 6400 35992 6412
rect 36044 6400 36050 6452
rect 24670 6332 24676 6384
rect 24728 6372 24734 6384
rect 30929 6375 30987 6381
rect 30929 6372 30941 6375
rect 24728 6344 30941 6372
rect 24728 6332 24734 6344
rect 30929 6341 30941 6344
rect 30975 6372 30987 6375
rect 32122 6372 32128 6384
rect 30975 6344 32128 6372
rect 30975 6341 30987 6344
rect 30929 6335 30987 6341
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6273 20407 6307
rect 22370 6304 22376 6316
rect 22331 6276 22376 6304
rect 20349 6267 20407 6273
rect 22370 6264 22376 6276
rect 22428 6264 22434 6316
rect 24854 6264 24860 6316
rect 24912 6304 24918 6316
rect 25222 6304 25228 6316
rect 24912 6276 25228 6304
rect 24912 6264 24918 6276
rect 25222 6264 25228 6276
rect 25280 6264 25286 6316
rect 26602 6264 26608 6316
rect 26660 6304 26666 6316
rect 26789 6307 26847 6313
rect 26789 6304 26801 6307
rect 26660 6276 26801 6304
rect 26660 6264 26666 6276
rect 26789 6273 26801 6276
rect 26835 6273 26847 6307
rect 26789 6267 26847 6273
rect 27065 6307 27123 6313
rect 27065 6273 27077 6307
rect 27111 6304 27123 6307
rect 27522 6304 27528 6316
rect 27111 6276 27528 6304
rect 27111 6273 27123 6276
rect 27065 6267 27123 6273
rect 27522 6264 27528 6276
rect 27580 6264 27586 6316
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9272 6208 9965 6236
rect 9272 6196 9278 6208
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 10226 6236 10232 6248
rect 10187 6208 10232 6236
rect 9953 6199 10011 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6236 11391 6239
rect 11379 6208 11928 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 1949 6171 2007 6177
rect 1949 6137 1961 6171
rect 1995 6168 2007 6171
rect 2222 6168 2228 6180
rect 1995 6140 2228 6168
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 2222 6128 2228 6140
rect 2280 6168 2286 6180
rect 2403 6171 2461 6177
rect 2403 6168 2415 6171
rect 2280 6140 2415 6168
rect 2280 6128 2286 6140
rect 2403 6137 2415 6140
rect 2449 6168 2461 6171
rect 3329 6171 3387 6177
rect 3329 6168 3341 6171
rect 2449 6140 3341 6168
rect 2449 6137 2461 6140
rect 2403 6131 2461 6137
rect 3329 6137 3341 6140
rect 3375 6168 3387 6171
rect 4154 6168 4160 6180
rect 3375 6140 4160 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 5350 6128 5356 6180
rect 5408 6168 5414 6180
rect 5408 6140 5453 6168
rect 5408 6128 5414 6140
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 6963 6171 7021 6177
rect 6963 6168 6975 6171
rect 5592 6140 6975 6168
rect 5592 6128 5598 6140
rect 6963 6137 6975 6140
rect 7009 6137 7021 6171
rect 7745 6171 7803 6177
rect 7745 6168 7757 6171
rect 6963 6131 7021 6137
rect 7110 6140 7757 6168
rect 2958 6100 2964 6112
rect 2919 6072 2964 6100
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 3927 6103 3985 6109
rect 3927 6100 3939 6103
rect 3844 6072 3939 6100
rect 3844 6060 3850 6072
rect 3927 6069 3939 6072
rect 3973 6069 3985 6103
rect 4614 6100 4620 6112
rect 4575 6072 4620 6100
rect 3927 6063 3985 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5368 6100 5396 6128
rect 5123 6072 5396 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 7110 6100 7138 6140
rect 7745 6137 7757 6140
rect 7791 6168 7803 6171
rect 8018 6168 8024 6180
rect 7791 6140 8024 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 8018 6128 8024 6140
rect 8076 6128 8082 6180
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8849 6171 8907 6177
rect 8352 6140 8397 6168
rect 8352 6128 8358 6140
rect 8849 6137 8861 6171
rect 8895 6168 8907 6171
rect 10502 6168 10508 6180
rect 8895 6140 10508 6168
rect 8895 6137 8907 6140
rect 8849 6131 8907 6137
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 11900 6112 11928 6208
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13412 6208 13921 6236
rect 13412 6196 13418 6208
rect 13909 6205 13921 6208
rect 13955 6236 13967 6239
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13955 6208 14105 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 21729 6239 21787 6245
rect 21729 6205 21741 6239
rect 21775 6236 21787 6239
rect 22094 6236 22100 6248
rect 21775 6208 22100 6236
rect 21775 6205 21787 6208
rect 21729 6199 21787 6205
rect 22094 6196 22100 6208
rect 22152 6196 22158 6248
rect 22278 6236 22284 6248
rect 22239 6208 22284 6236
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23492 6208 23673 6236
rect 12621 6171 12679 6177
rect 12621 6137 12633 6171
rect 12667 6137 12679 6171
rect 13998 6168 14004 6180
rect 13959 6140 14004 6168
rect 12621 6131 12679 6137
rect 9582 6100 9588 6112
rect 6328 6072 7138 6100
rect 9543 6072 9588 6100
rect 6328 6060 6334 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12158 6100 12164 6112
rect 12119 6072 12164 6100
rect 12158 6060 12164 6072
rect 12216 6100 12222 6112
rect 12636 6100 12664 6131
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 16117 6171 16175 6177
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 16206 6168 16212 6180
rect 16163 6140 16212 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 16206 6128 16212 6140
rect 16264 6168 16270 6180
rect 16571 6171 16629 6177
rect 16571 6168 16583 6171
rect 16264 6140 16583 6168
rect 16264 6128 16270 6140
rect 16571 6137 16583 6140
rect 16617 6168 16629 6171
rect 16942 6168 16948 6180
rect 16617 6140 16948 6168
rect 16617 6137 16629 6140
rect 16571 6131 16629 6137
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 17862 6168 17868 6180
rect 17775 6140 17868 6168
rect 17862 6128 17868 6140
rect 17920 6168 17926 6180
rect 18782 6168 18788 6180
rect 17920 6140 18644 6168
rect 18743 6140 18788 6168
rect 17920 6128 17926 6140
rect 12216 6072 12664 6100
rect 15381 6103 15439 6109
rect 12216 6060 12222 6072
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 15470 6100 15476 6112
rect 15427 6072 15476 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 18616 6100 18644 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 18877 6171 18935 6177
rect 18877 6137 18889 6171
rect 18923 6137 18935 6171
rect 19426 6168 19432 6180
rect 19339 6140 19432 6168
rect 18877 6131 18935 6137
rect 18892 6100 18920 6131
rect 19426 6128 19432 6140
rect 19484 6168 19490 6180
rect 19484 6140 20392 6168
rect 19484 6128 19490 6140
rect 18616 6072 18920 6100
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 19576 6072 20085 6100
rect 19576 6060 19582 6072
rect 20073 6069 20085 6072
rect 20119 6100 20131 6103
rect 20254 6100 20260 6112
rect 20119 6072 20260 6100
rect 20119 6069 20131 6072
rect 20073 6063 20131 6069
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 20364 6100 20392 6140
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 20990 6168 20996 6180
rect 20496 6140 20541 6168
rect 20640 6140 20996 6168
rect 20496 6128 20502 6140
rect 20640 6100 20668 6140
rect 20990 6128 20996 6140
rect 21048 6128 21054 6180
rect 23492 6112 23520 6208
rect 23661 6205 23673 6208
rect 23707 6205 23719 6239
rect 23661 6199 23719 6205
rect 23750 6196 23756 6248
rect 23808 6236 23814 6248
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23808 6208 24225 6236
rect 23808 6196 23814 6208
rect 24213 6205 24225 6208
rect 24259 6236 24271 6239
rect 24762 6236 24768 6248
rect 24259 6208 24768 6236
rect 24259 6205 24271 6208
rect 24213 6199 24271 6205
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 28905 6239 28963 6245
rect 28905 6205 28917 6239
rect 28951 6236 28963 6239
rect 29273 6239 29331 6245
rect 29273 6236 29285 6239
rect 28951 6208 29285 6236
rect 28951 6205 28963 6208
rect 28905 6199 28963 6205
rect 29273 6205 29285 6208
rect 29319 6205 29331 6239
rect 29730 6236 29736 6248
rect 29691 6208 29736 6236
rect 29273 6199 29331 6205
rect 29730 6196 29736 6208
rect 29788 6196 29794 6248
rect 30944 6236 30972 6335
rect 32122 6332 32128 6344
rect 32180 6332 32186 6384
rect 33873 6375 33931 6381
rect 33873 6341 33885 6375
rect 33919 6372 33931 6375
rect 35066 6372 35072 6384
rect 33919 6344 35072 6372
rect 33919 6341 33931 6344
rect 33873 6335 33931 6341
rect 35066 6332 35072 6344
rect 35124 6372 35130 6384
rect 35124 6344 35572 6372
rect 35124 6332 35130 6344
rect 33318 6304 33324 6316
rect 33231 6276 33324 6304
rect 33318 6264 33324 6276
rect 33376 6304 33382 6316
rect 33686 6304 33692 6316
rect 33376 6276 33692 6304
rect 33376 6264 33382 6276
rect 33686 6264 33692 6276
rect 33744 6264 33750 6316
rect 34977 6307 35035 6313
rect 34977 6273 34989 6307
rect 35023 6304 35035 6307
rect 35434 6304 35440 6316
rect 35023 6276 35440 6304
rect 35023 6273 35035 6276
rect 34977 6267 35035 6273
rect 35434 6264 35440 6276
rect 35492 6264 35498 6316
rect 35544 6304 35572 6344
rect 36817 6307 36875 6313
rect 36817 6304 36829 6307
rect 35544 6276 36829 6304
rect 36817 6273 36829 6276
rect 36863 6273 36875 6307
rect 36817 6267 36875 6273
rect 31113 6239 31171 6245
rect 31113 6236 31125 6239
rect 30944 6208 31125 6236
rect 31113 6205 31125 6208
rect 31159 6205 31171 6239
rect 31113 6199 31171 6205
rect 31202 6196 31208 6248
rect 31260 6236 31266 6248
rect 31570 6236 31576 6248
rect 31260 6208 31576 6236
rect 31260 6196 31266 6208
rect 31570 6196 31576 6208
rect 31628 6196 31634 6248
rect 24397 6171 24455 6177
rect 24397 6137 24409 6171
rect 24443 6168 24455 6171
rect 25406 6168 25412 6180
rect 24443 6140 25412 6168
rect 24443 6137 24455 6140
rect 24397 6131 24455 6137
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 26513 6171 26571 6177
rect 25884 6140 26280 6168
rect 25884 6112 25912 6140
rect 20364 6072 20668 6100
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21269 6103 21327 6109
rect 21269 6100 21281 6103
rect 20772 6072 21281 6100
rect 20772 6060 20778 6072
rect 21269 6069 21281 6072
rect 21315 6069 21327 6103
rect 21269 6063 21327 6069
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 22738 6100 22744 6112
rect 22612 6072 22744 6100
rect 22612 6060 22618 6072
rect 22738 6060 22744 6072
rect 22796 6100 22802 6112
rect 22833 6103 22891 6109
rect 22833 6100 22845 6103
rect 22796 6072 22845 6100
rect 22796 6060 22802 6072
rect 22833 6069 22845 6072
rect 22879 6069 22891 6103
rect 23474 6100 23480 6112
rect 23435 6072 23480 6100
rect 22833 6063 22891 6069
rect 23474 6060 23480 6072
rect 23532 6060 23538 6112
rect 24949 6103 25007 6109
rect 24949 6069 24961 6103
rect 24995 6100 25007 6103
rect 25593 6103 25651 6109
rect 25593 6100 25605 6103
rect 24995 6072 25605 6100
rect 24995 6069 25007 6072
rect 24949 6063 25007 6069
rect 25593 6069 25605 6072
rect 25639 6100 25651 6103
rect 25866 6100 25872 6112
rect 25639 6072 25872 6100
rect 25639 6069 25651 6072
rect 25593 6063 25651 6069
rect 25866 6060 25872 6072
rect 25924 6060 25930 6112
rect 26142 6100 26148 6112
rect 26103 6072 26148 6100
rect 26142 6060 26148 6072
rect 26200 6060 26206 6112
rect 26252 6100 26280 6140
rect 26513 6137 26525 6171
rect 26559 6168 26571 6171
rect 26878 6168 26884 6180
rect 26559 6140 26884 6168
rect 26559 6137 26571 6140
rect 26513 6131 26571 6137
rect 26878 6128 26884 6140
rect 26936 6168 26942 6180
rect 27157 6171 27215 6177
rect 27157 6168 27169 6171
rect 26936 6140 27169 6168
rect 26936 6128 26942 6140
rect 27157 6137 27169 6140
rect 27203 6137 27215 6171
rect 27157 6131 27215 6137
rect 27246 6128 27252 6180
rect 27304 6168 27310 6180
rect 27709 6171 27767 6177
rect 27709 6168 27721 6171
rect 27304 6140 27721 6168
rect 27304 6128 27310 6140
rect 27709 6137 27721 6140
rect 27755 6137 27767 6171
rect 27709 6131 27767 6137
rect 27798 6128 27804 6180
rect 27856 6168 27862 6180
rect 28445 6171 28503 6177
rect 28445 6168 28457 6171
rect 27856 6140 28457 6168
rect 27856 6128 27862 6140
rect 28445 6137 28457 6140
rect 28491 6168 28503 6171
rect 31846 6168 31852 6180
rect 28491 6140 29408 6168
rect 31807 6140 31852 6168
rect 28491 6137 28503 6140
rect 28445 6131 28503 6137
rect 27985 6103 28043 6109
rect 27985 6100 27997 6103
rect 26252 6072 27997 6100
rect 27985 6069 27997 6072
rect 28031 6100 28043 6103
rect 28810 6100 28816 6112
rect 28031 6072 28816 6100
rect 28031 6069 28043 6072
rect 27985 6063 28043 6069
rect 28810 6060 28816 6072
rect 28868 6060 28874 6112
rect 29380 6109 29408 6140
rect 31846 6128 31852 6140
rect 31904 6128 31910 6180
rect 33413 6171 33471 6177
rect 33413 6137 33425 6171
rect 33459 6137 33471 6171
rect 34609 6171 34667 6177
rect 34609 6168 34621 6171
rect 33413 6131 33471 6137
rect 34072 6140 34621 6168
rect 29365 6103 29423 6109
rect 29365 6069 29377 6103
rect 29411 6069 29423 6103
rect 30374 6100 30380 6112
rect 30335 6072 30380 6100
rect 29365 6063 29423 6069
rect 30374 6060 30380 6072
rect 30432 6060 30438 6112
rect 33042 6100 33048 6112
rect 33003 6072 33048 6100
rect 33042 6060 33048 6072
rect 33100 6100 33106 6112
rect 33428 6100 33456 6131
rect 34072 6100 34100 6140
rect 34609 6137 34621 6140
rect 34655 6137 34667 6171
rect 34609 6131 34667 6137
rect 35069 6171 35127 6177
rect 35069 6137 35081 6171
rect 35115 6137 35127 6171
rect 35069 6131 35127 6137
rect 35621 6171 35679 6177
rect 35621 6137 35633 6171
rect 35667 6168 35679 6171
rect 35986 6168 35992 6180
rect 35667 6140 35992 6168
rect 35667 6137 35679 6140
rect 35621 6131 35679 6137
rect 33100 6072 34100 6100
rect 34624 6100 34652 6131
rect 35084 6100 35112 6131
rect 35986 6128 35992 6140
rect 36044 6128 36050 6180
rect 36538 6168 36544 6180
rect 36499 6140 36544 6168
rect 36538 6128 36544 6140
rect 36596 6128 36602 6180
rect 36633 6171 36691 6177
rect 36633 6137 36645 6171
rect 36679 6137 36691 6171
rect 36633 6131 36691 6137
rect 34624 6072 35112 6100
rect 33100 6060 33106 6072
rect 35894 6060 35900 6112
rect 35952 6100 35958 6112
rect 36265 6103 36323 6109
rect 36265 6100 36277 6103
rect 35952 6072 36277 6100
rect 35952 6060 35958 6072
rect 36265 6069 36277 6072
rect 36311 6100 36323 6103
rect 36648 6100 36676 6131
rect 36311 6072 36676 6100
rect 36311 6069 36323 6072
rect 36265 6063 36323 6069
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 3234 5896 3240 5908
rect 2740 5868 3240 5896
rect 2740 5856 2746 5868
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 4985 5899 5043 5905
rect 4985 5865 4997 5899
rect 5031 5896 5043 5899
rect 5350 5896 5356 5908
rect 5031 5868 5356 5896
rect 5031 5865 5043 5868
rect 4985 5859 5043 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 7466 5896 7472 5908
rect 7427 5868 7472 5896
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8352 5868 8861 5896
rect 8352 5856 8358 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12492 5868 12817 5896
rect 12492 5856 12498 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 13538 5856 13544 5908
rect 13596 5896 13602 5908
rect 14642 5896 14648 5908
rect 13596 5868 14228 5896
rect 14603 5868 14648 5896
rect 13596 5856 13602 5868
rect 1857 5831 1915 5837
rect 1857 5797 1869 5831
rect 1903 5828 1915 5831
rect 2222 5828 2228 5840
rect 1903 5800 2228 5828
rect 1903 5797 1915 5800
rect 1857 5791 1915 5797
rect 2222 5788 2228 5800
rect 2280 5837 2286 5840
rect 2280 5831 2328 5837
rect 2280 5797 2282 5831
rect 2316 5797 2328 5831
rect 2280 5791 2328 5797
rect 2280 5788 2286 5791
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 4427 5831 4485 5837
rect 4427 5828 4439 5831
rect 4212 5800 4439 5828
rect 4212 5788 4218 5800
rect 4427 5797 4439 5800
rect 4473 5828 4485 5831
rect 5077 5831 5135 5837
rect 5077 5828 5089 5831
rect 4473 5800 5089 5828
rect 4473 5797 4485 5800
rect 4427 5791 4485 5797
rect 5077 5797 5089 5800
rect 5123 5797 5135 5831
rect 5077 5791 5135 5797
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5629 5831 5687 5837
rect 5629 5828 5641 5831
rect 5316 5800 5641 5828
rect 5316 5788 5322 5800
rect 5629 5797 5641 5800
rect 5675 5797 5687 5831
rect 6270 5828 6276 5840
rect 6231 5800 6276 5828
rect 5629 5791 5687 5797
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 8036 5828 8064 5856
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 7340 5800 8064 5828
rect 9600 5800 9873 5828
rect 7340 5788 7346 5800
rect 1946 5760 1952 5772
rect 1907 5732 1952 5760
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 4614 5760 4620 5772
rect 2915 5732 4620 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 5350 5760 5356 5772
rect 5311 5732 5356 5760
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7248 5732 7665 5760
rect 7248 5720 7254 5732
rect 7653 5729 7665 5732
rect 7699 5760 7711 5763
rect 8110 5760 8116 5772
rect 7699 5732 8116 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 8573 5763 8631 5769
rect 8573 5729 8585 5763
rect 8619 5760 8631 5763
rect 9600 5760 9628 5800
rect 9861 5797 9873 5800
rect 9907 5828 9919 5831
rect 10410 5828 10416 5840
rect 9907 5800 10416 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11879 5831 11937 5837
rect 11879 5828 11891 5831
rect 11204 5800 11891 5828
rect 11204 5788 11210 5800
rect 11879 5797 11891 5800
rect 11925 5828 11937 5831
rect 11974 5828 11980 5840
rect 11925 5800 11980 5828
rect 11925 5797 11937 5800
rect 11879 5791 11937 5797
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 13354 5828 13360 5840
rect 12452 5800 13360 5828
rect 12452 5772 12480 5800
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 13449 5831 13507 5837
rect 13449 5797 13461 5831
rect 13495 5828 13507 5831
rect 13998 5828 14004 5840
rect 13495 5800 14004 5828
rect 13495 5797 13507 5800
rect 13449 5791 13507 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 14200 5828 14228 5868
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 16206 5896 16212 5908
rect 16167 5868 16212 5896
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 16298 5856 16304 5908
rect 16356 5896 16362 5908
rect 16850 5896 16856 5908
rect 16356 5868 16856 5896
rect 16356 5856 16362 5868
rect 16850 5856 16856 5868
rect 16908 5896 16914 5908
rect 17589 5899 17647 5905
rect 17589 5896 17601 5899
rect 16908 5868 17601 5896
rect 16908 5856 16914 5868
rect 17589 5865 17601 5868
rect 17635 5865 17647 5899
rect 22189 5899 22247 5905
rect 22189 5896 22201 5899
rect 17589 5859 17647 5865
rect 18202 5868 22201 5896
rect 15013 5831 15071 5837
rect 15013 5828 15025 5831
rect 14200 5800 15025 5828
rect 15013 5797 15025 5800
rect 15059 5797 15071 5831
rect 16224 5828 16252 5856
rect 16714 5831 16772 5837
rect 16714 5828 16726 5831
rect 16224 5800 16726 5828
rect 15013 5791 15071 5797
rect 16714 5797 16726 5800
rect 16760 5797 16772 5831
rect 16714 5791 16772 5797
rect 17494 5788 17500 5840
rect 17552 5828 17558 5840
rect 18202 5828 18230 5868
rect 22189 5865 22201 5868
rect 22235 5865 22247 5899
rect 22370 5896 22376 5908
rect 22331 5868 22376 5896
rect 22189 5859 22247 5865
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 23474 5896 23480 5908
rect 22756 5868 23480 5896
rect 18785 5831 18843 5837
rect 18785 5828 18797 5831
rect 17552 5800 18230 5828
rect 18432 5800 18797 5828
rect 17552 5788 17558 5800
rect 12434 5760 12440 5772
rect 8619 5732 9628 5760
rect 12347 5732 12440 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 15378 5760 15384 5772
rect 15339 5732 15384 5760
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 18432 5769 18460 5800
rect 18785 5797 18797 5800
rect 18831 5828 18843 5831
rect 20257 5831 20315 5837
rect 20257 5828 20269 5831
rect 18831 5800 20269 5828
rect 18831 5797 18843 5800
rect 18785 5791 18843 5797
rect 20257 5797 20269 5800
rect 20303 5828 20315 5831
rect 20438 5828 20444 5840
rect 20303 5800 20444 5828
rect 20303 5797 20315 5800
rect 20257 5791 20315 5797
rect 20438 5788 20444 5800
rect 20496 5788 20502 5840
rect 20530 5788 20536 5840
rect 20588 5828 20594 5840
rect 21085 5831 21143 5837
rect 21085 5828 21097 5831
rect 20588 5800 21097 5828
rect 20588 5788 20594 5800
rect 21085 5797 21097 5800
rect 21131 5797 21143 5831
rect 21634 5828 21640 5840
rect 21547 5800 21640 5828
rect 21085 5791 21143 5797
rect 21634 5788 21640 5800
rect 21692 5828 21698 5840
rect 22646 5828 22652 5840
rect 21692 5800 22652 5828
rect 21692 5788 21698 5800
rect 22646 5788 22652 5800
rect 22704 5788 22710 5840
rect 22756 5769 22784 5868
rect 23474 5856 23480 5868
rect 23532 5856 23538 5908
rect 23750 5896 23756 5908
rect 23711 5868 23756 5896
rect 23750 5856 23756 5868
rect 23808 5856 23814 5908
rect 24394 5896 24400 5908
rect 24355 5868 24400 5896
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 25222 5896 25228 5908
rect 25183 5868 25228 5896
rect 25222 5856 25228 5868
rect 25280 5856 25286 5908
rect 25406 5856 25412 5908
rect 25464 5896 25470 5908
rect 29546 5896 29552 5908
rect 25464 5868 29552 5896
rect 25464 5856 25470 5868
rect 29546 5856 29552 5868
rect 29604 5896 29610 5908
rect 29641 5899 29699 5905
rect 29641 5896 29653 5899
rect 29604 5868 29653 5896
rect 29604 5856 29610 5868
rect 29641 5865 29653 5868
rect 29687 5865 29699 5899
rect 29641 5859 29699 5865
rect 31205 5899 31263 5905
rect 31205 5865 31217 5899
rect 31251 5896 31263 5899
rect 33042 5896 33048 5908
rect 31251 5868 33048 5896
rect 31251 5865 31263 5868
rect 31205 5859 31263 5865
rect 33042 5856 33048 5868
rect 33100 5856 33106 5908
rect 33778 5896 33784 5908
rect 33739 5868 33784 5896
rect 33778 5856 33784 5868
rect 33836 5856 33842 5908
rect 34146 5856 34152 5908
rect 34204 5896 34210 5908
rect 34241 5899 34299 5905
rect 34241 5896 34253 5899
rect 34204 5868 34253 5896
rect 34204 5856 34210 5868
rect 34241 5865 34253 5868
rect 34287 5865 34299 5899
rect 34790 5896 34796 5908
rect 34751 5868 34796 5896
rect 34241 5859 34299 5865
rect 34790 5856 34796 5868
rect 34848 5856 34854 5908
rect 36538 5856 36544 5908
rect 36596 5896 36602 5908
rect 36633 5899 36691 5905
rect 36633 5896 36645 5899
rect 36596 5868 36645 5896
rect 36596 5856 36602 5868
rect 36633 5865 36645 5868
rect 36679 5865 36691 5899
rect 36633 5859 36691 5865
rect 23201 5831 23259 5837
rect 23201 5797 23213 5831
rect 23247 5828 23259 5831
rect 23842 5828 23848 5840
rect 23247 5800 23848 5828
rect 23247 5797 23259 5800
rect 23201 5791 23259 5797
rect 23842 5788 23848 5800
rect 23900 5788 23906 5840
rect 26694 5828 26700 5840
rect 26655 5800 26700 5828
rect 26694 5788 26700 5800
rect 26752 5788 26758 5840
rect 28258 5828 28264 5840
rect 28219 5800 28264 5828
rect 28258 5788 28264 5800
rect 28316 5788 28322 5840
rect 30374 5788 30380 5840
rect 30432 5828 30438 5840
rect 32490 5837 32496 5840
rect 30647 5831 30705 5837
rect 30647 5828 30659 5831
rect 30432 5800 30659 5828
rect 30432 5788 30438 5800
rect 30647 5797 30659 5800
rect 30693 5828 30705 5831
rect 32487 5828 32496 5837
rect 30693 5800 32496 5828
rect 30693 5797 30705 5800
rect 30647 5791 30705 5797
rect 32487 5791 32496 5800
rect 32490 5788 32496 5791
rect 32548 5788 32554 5840
rect 33134 5788 33140 5840
rect 33192 5828 33198 5840
rect 35805 5831 35863 5837
rect 35805 5828 35817 5831
rect 33192 5800 35817 5828
rect 33192 5788 33198 5800
rect 35805 5797 35817 5800
rect 35851 5828 35863 5831
rect 35894 5828 35900 5840
rect 35851 5800 35900 5828
rect 35851 5797 35863 5800
rect 35805 5791 35863 5797
rect 35894 5788 35900 5800
rect 35952 5788 35958 5840
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 16080 5732 16405 5760
rect 16080 5720 16086 5732
rect 16393 5729 16405 5732
rect 16439 5729 16451 5763
rect 16393 5723 16451 5729
rect 17313 5763 17371 5769
rect 17313 5729 17325 5763
rect 17359 5760 17371 5763
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 17359 5732 18429 5760
rect 17359 5729 17371 5732
rect 17313 5723 17371 5729
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5760 22247 5763
rect 22741 5763 22799 5769
rect 22741 5760 22753 5763
rect 22235 5732 22753 5760
rect 22235 5729 22247 5732
rect 22189 5723 22247 5729
rect 22741 5729 22753 5732
rect 22787 5729 22799 5763
rect 22741 5723 22799 5729
rect 22925 5763 22983 5769
rect 22925 5729 22937 5763
rect 22971 5729 22983 5763
rect 22925 5723 22983 5729
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 2832 5664 4077 5692
rect 2832 5652 2838 5664
rect 4065 5661 4077 5664
rect 4111 5692 4123 5695
rect 5442 5692 5448 5704
rect 4111 5664 5448 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6362 5692 6368 5704
rect 6227 5664 6368 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 6503 5664 9413 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 9401 5661 9413 5664
rect 9447 5692 9459 5695
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9447 5664 9781 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10502 5692 10508 5704
rect 10459 5664 10508 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 5902 5584 5908 5636
rect 5960 5624 5966 5636
rect 6472 5624 6500 5655
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11348 5664 11529 5692
rect 5960 5596 6500 5624
rect 5960 5584 5966 5596
rect 11348 5568 11376 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 12308 5664 13369 5692
rect 12308 5652 12314 5664
rect 13357 5661 13369 5664
rect 13403 5692 13415 5695
rect 13538 5692 13544 5704
rect 13403 5664 13544 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 16408 5692 16436 5723
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 16408 5664 17969 5692
rect 17957 5661 17969 5664
rect 18003 5661 18015 5695
rect 18690 5692 18696 5704
rect 18651 5664 18696 5692
rect 17957 5655 18015 5661
rect 18690 5652 18696 5664
rect 18748 5652 18754 5704
rect 19058 5692 19064 5704
rect 19019 5664 19064 5692
rect 19058 5652 19064 5664
rect 19116 5652 19122 5704
rect 20990 5692 20996 5704
rect 20903 5664 20996 5692
rect 20990 5652 20996 5664
rect 21048 5692 21054 5704
rect 21910 5692 21916 5704
rect 21048 5664 21916 5692
rect 21048 5652 21054 5664
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 22278 5652 22284 5704
rect 22336 5692 22342 5704
rect 22940 5692 22968 5723
rect 32858 5720 32864 5772
rect 32916 5760 32922 5772
rect 32916 5732 33916 5760
rect 32916 5720 32922 5732
rect 33888 5704 33916 5732
rect 24026 5692 24032 5704
rect 22336 5664 22968 5692
rect 23987 5664 24032 5692
rect 22336 5652 22342 5664
rect 24026 5652 24032 5664
rect 24084 5652 24090 5704
rect 25958 5652 25964 5704
rect 26016 5692 26022 5704
rect 26605 5695 26663 5701
rect 26605 5692 26617 5695
rect 26016 5664 26617 5692
rect 26016 5652 26022 5664
rect 26605 5661 26617 5664
rect 26651 5661 26663 5695
rect 27246 5692 27252 5704
rect 27207 5664 27252 5692
rect 26605 5655 26663 5661
rect 27246 5652 27252 5664
rect 27304 5652 27310 5704
rect 28166 5692 28172 5704
rect 28127 5664 28172 5692
rect 28166 5652 28172 5664
rect 28224 5692 28230 5704
rect 28350 5692 28356 5704
rect 28224 5664 28356 5692
rect 28224 5652 28230 5664
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 28445 5695 28503 5701
rect 28445 5661 28457 5695
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 30285 5695 30343 5701
rect 30285 5661 30297 5695
rect 30331 5692 30343 5695
rect 30466 5692 30472 5704
rect 30331 5664 30472 5692
rect 30331 5661 30343 5664
rect 30285 5655 30343 5661
rect 12526 5584 12532 5636
rect 12584 5624 12590 5636
rect 13722 5624 13728 5636
rect 12584 5596 13728 5624
rect 12584 5584 12590 5596
rect 13722 5584 13728 5596
rect 13780 5624 13786 5636
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 13780 5596 13921 5624
rect 13780 5584 13786 5596
rect 13909 5593 13921 5596
rect 13955 5593 13967 5627
rect 13909 5587 13967 5593
rect 15565 5627 15623 5633
rect 15565 5593 15577 5627
rect 15611 5624 15623 5627
rect 21818 5624 21824 5636
rect 15611 5596 21824 5624
rect 15611 5593 15623 5596
rect 15565 5587 15623 5593
rect 21818 5584 21824 5596
rect 21876 5624 21882 5636
rect 22094 5624 22100 5636
rect 21876 5596 22100 5624
rect 21876 5584 21882 5596
rect 22094 5584 22100 5596
rect 22152 5584 22158 5636
rect 5077 5559 5135 5565
rect 5077 5525 5089 5559
rect 5123 5556 5135 5559
rect 7282 5556 7288 5568
rect 5123 5528 7288 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 10962 5556 10968 5568
rect 10923 5528 10968 5556
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11330 5556 11336 5568
rect 11291 5528 11336 5556
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 13596 5528 14289 5556
rect 13596 5516 13602 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 15838 5556 15844 5568
rect 15799 5528 15844 5556
rect 14277 5519 14335 5525
rect 15838 5516 15844 5528
rect 15896 5516 15902 5568
rect 19610 5556 19616 5568
rect 19571 5528 19616 5556
rect 19610 5516 19616 5528
rect 19668 5516 19674 5568
rect 20622 5556 20628 5568
rect 20583 5528 20628 5556
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 21450 5516 21456 5568
rect 21508 5556 21514 5568
rect 21913 5559 21971 5565
rect 21913 5556 21925 5559
rect 21508 5528 21925 5556
rect 21508 5516 21514 5528
rect 21913 5525 21925 5528
rect 21959 5525 21971 5559
rect 24946 5556 24952 5568
rect 24907 5528 24952 5556
rect 21913 5519 21971 5525
rect 24946 5516 24952 5528
rect 25004 5516 25010 5568
rect 26050 5516 26056 5568
rect 26108 5556 26114 5568
rect 27062 5556 27068 5568
rect 26108 5528 27068 5556
rect 26108 5516 26114 5528
rect 27062 5516 27068 5528
rect 27120 5516 27126 5568
rect 28166 5516 28172 5568
rect 28224 5556 28230 5568
rect 28460 5556 28488 5655
rect 30466 5652 30472 5664
rect 30524 5652 30530 5704
rect 31570 5652 31576 5704
rect 31628 5692 31634 5704
rect 32125 5695 32183 5701
rect 32125 5692 32137 5695
rect 31628 5664 32137 5692
rect 31628 5652 31634 5664
rect 32125 5661 32137 5664
rect 32171 5661 32183 5695
rect 32125 5655 32183 5661
rect 32398 5652 32404 5704
rect 32456 5692 32462 5704
rect 32456 5664 33824 5692
rect 32456 5652 32462 5664
rect 33796 5624 33824 5664
rect 33870 5652 33876 5704
rect 33928 5692 33934 5704
rect 35713 5695 35771 5701
rect 35713 5692 35725 5695
rect 33928 5664 33973 5692
rect 35084 5664 35725 5692
rect 33928 5652 33934 5664
rect 35084 5633 35112 5664
rect 35713 5661 35725 5664
rect 35759 5661 35771 5695
rect 35986 5692 35992 5704
rect 35947 5664 35992 5692
rect 35713 5655 35771 5661
rect 35986 5652 35992 5664
rect 36044 5652 36050 5704
rect 35069 5627 35127 5633
rect 35069 5624 35081 5627
rect 33796 5596 35081 5624
rect 35069 5593 35081 5596
rect 35115 5593 35127 5627
rect 35069 5587 35127 5593
rect 28224 5528 28488 5556
rect 28224 5516 28230 5528
rect 28626 5516 28632 5568
rect 28684 5556 28690 5568
rect 29273 5559 29331 5565
rect 29273 5556 29285 5559
rect 28684 5528 29285 5556
rect 28684 5516 28690 5528
rect 29273 5525 29285 5528
rect 29319 5556 29331 5559
rect 29730 5556 29736 5568
rect 29319 5528 29736 5556
rect 29319 5525 29331 5528
rect 29273 5519 29331 5525
rect 29730 5516 29736 5528
rect 29788 5516 29794 5568
rect 33042 5556 33048 5568
rect 33003 5528 33048 5556
rect 33042 5516 33048 5528
rect 33100 5516 33106 5568
rect 35250 5516 35256 5568
rect 35308 5556 35314 5568
rect 35437 5559 35495 5565
rect 35437 5556 35449 5559
rect 35308 5528 35449 5556
rect 35308 5516 35314 5528
rect 35437 5525 35449 5528
rect 35483 5525 35495 5559
rect 35437 5519 35495 5525
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1486 5312 1492 5364
rect 1544 5352 1550 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1544 5324 1593 5352
rect 1544 5312 1550 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 5442 5352 5448 5364
rect 3016 5324 4154 5352
rect 5403 5324 5448 5352
rect 3016 5312 3022 5324
rect 4126 5284 4154 5324
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 6454 5352 6460 5364
rect 6415 5324 6460 5352
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 7190 5352 7196 5364
rect 7151 5324 7196 5352
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8573 5355 8631 5361
rect 8573 5352 8585 5355
rect 8352 5324 8585 5352
rect 8352 5312 8358 5324
rect 8573 5321 8585 5324
rect 8619 5321 8631 5355
rect 8573 5315 8631 5321
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9766 5352 9772 5364
rect 8987 5324 9772 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 6089 5287 6147 5293
rect 6089 5284 6101 5287
rect 4126 5256 6101 5284
rect 6089 5253 6101 5256
rect 6135 5284 6147 5287
rect 6270 5284 6276 5296
rect 6135 5256 6276 5284
rect 6135 5253 6147 5256
rect 6089 5247 6147 5253
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 3844 5188 4537 5216
rect 3844 5176 3850 5188
rect 4525 5185 4537 5188
rect 4571 5185 4583 5219
rect 4890 5216 4896 5228
rect 4851 5188 4896 5216
rect 4525 5179 4583 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 8956 5216 8984 5315
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10410 5352 10416 5364
rect 10371 5324 10416 5352
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 12618 5352 12624 5364
rect 12531 5324 12624 5352
rect 12618 5312 12624 5324
rect 12676 5352 12682 5364
rect 13078 5352 13084 5364
rect 12676 5324 13084 5352
rect 12676 5312 12682 5324
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 15286 5352 15292 5364
rect 13188 5324 15292 5352
rect 11609 5287 11667 5293
rect 11609 5253 11621 5287
rect 11655 5284 11667 5287
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 11655 5256 11897 5284
rect 11655 5253 11667 5256
rect 11609 5247 11667 5253
rect 11885 5253 11897 5256
rect 11931 5284 11943 5287
rect 13188 5284 13216 5324
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 16206 5312 16212 5364
rect 16264 5352 16270 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 16264 5324 16405 5352
rect 16264 5312 16270 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 16393 5315 16451 5321
rect 17037 5355 17095 5361
rect 17037 5321 17049 5355
rect 17083 5352 17095 5355
rect 17494 5352 17500 5364
rect 17083 5324 17500 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 22005 5355 22063 5361
rect 22005 5352 22017 5355
rect 18748 5324 22017 5352
rect 18748 5312 18754 5324
rect 22005 5321 22017 5324
rect 22051 5321 22063 5355
rect 22005 5315 22063 5321
rect 22738 5312 22744 5364
rect 22796 5352 22802 5364
rect 23293 5355 23351 5361
rect 23293 5352 23305 5355
rect 22796 5324 23305 5352
rect 22796 5312 22802 5324
rect 23293 5321 23305 5324
rect 23339 5352 23351 5355
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 23339 5324 23397 5352
rect 23339 5321 23351 5324
rect 23293 5315 23351 5321
rect 23385 5321 23397 5324
rect 23431 5321 23443 5355
rect 23385 5315 23443 5321
rect 24946 5312 24952 5364
rect 25004 5352 25010 5364
rect 26329 5355 26387 5361
rect 26329 5352 26341 5355
rect 25004 5324 26341 5352
rect 25004 5312 25010 5324
rect 26329 5321 26341 5324
rect 26375 5352 26387 5355
rect 26694 5352 26700 5364
rect 26375 5324 26700 5352
rect 26375 5321 26387 5324
rect 26329 5315 26387 5321
rect 26694 5312 26700 5324
rect 26752 5352 26758 5364
rect 28077 5355 28135 5361
rect 28077 5352 28089 5355
rect 26752 5324 28089 5352
rect 26752 5312 26758 5324
rect 28077 5321 28089 5324
rect 28123 5352 28135 5355
rect 28258 5352 28264 5364
rect 28123 5324 28264 5352
rect 28123 5321 28135 5324
rect 28077 5315 28135 5321
rect 28258 5312 28264 5324
rect 28316 5312 28322 5364
rect 28350 5312 28356 5364
rect 28408 5352 28414 5364
rect 28445 5355 28503 5361
rect 28445 5352 28457 5355
rect 28408 5324 28457 5352
rect 28408 5312 28414 5324
rect 28445 5321 28457 5324
rect 28491 5321 28503 5355
rect 31018 5352 31024 5364
rect 30931 5324 31024 5352
rect 28445 5315 28503 5321
rect 31018 5312 31024 5324
rect 31076 5352 31082 5364
rect 31294 5352 31300 5364
rect 31076 5324 31300 5352
rect 31076 5312 31082 5324
rect 31294 5312 31300 5324
rect 31352 5312 31358 5364
rect 33870 5312 33876 5364
rect 33928 5352 33934 5364
rect 34241 5355 34299 5361
rect 34241 5352 34253 5355
rect 33928 5324 34253 5352
rect 33928 5312 33934 5324
rect 34241 5321 34253 5324
rect 34287 5321 34299 5355
rect 35894 5352 35900 5364
rect 35855 5324 35900 5352
rect 34241 5315 34299 5321
rect 35894 5312 35900 5324
rect 35952 5312 35958 5364
rect 11931 5256 13216 5284
rect 13449 5287 13507 5293
rect 11931 5253 11943 5256
rect 11885 5247 11943 5253
rect 13449 5253 13461 5287
rect 13495 5284 13507 5287
rect 16224 5284 16252 5312
rect 13495 5256 16252 5284
rect 13495 5253 13507 5256
rect 13449 5247 13507 5253
rect 7699 5188 8984 5216
rect 9309 5219 9367 5225
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 9355 5188 9674 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1949 5151 2007 5157
rect 1949 5148 1961 5151
rect 1443 5120 1961 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 1949 5117 1961 5120
rect 1995 5148 2007 5151
rect 2590 5148 2596 5160
rect 1995 5120 2596 5148
rect 1995 5117 2007 5120
rect 1949 5111 2007 5117
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 2866 5148 2872 5160
rect 2731 5120 2872 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 3970 5148 3976 5160
rect 3651 5120 3976 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 3970 5108 3976 5120
rect 4028 5148 4034 5160
rect 4028 5120 4384 5148
rect 4028 5108 4034 5120
rect 2498 5080 2504 5092
rect 2411 5052 2504 5080
rect 2498 5040 2504 5052
rect 2556 5080 2562 5092
rect 3047 5083 3105 5089
rect 3047 5080 3059 5083
rect 2556 5052 3059 5080
rect 2556 5040 2562 5052
rect 3047 5049 3059 5052
rect 3093 5080 3105 5083
rect 4154 5080 4160 5092
rect 3093 5052 4160 5080
rect 3093 5049 3105 5052
rect 3047 5043 3105 5049
rect 4154 5040 4160 5052
rect 4212 5080 4218 5092
rect 4212 5052 4257 5080
rect 4212 5040 4218 5052
rect 4356 5012 4384 5120
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 9324 5148 9352 5179
rect 6788 5120 9352 5148
rect 6788 5108 6794 5120
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9493 5151 9551 5157
rect 9493 5148 9505 5151
rect 9456 5120 9505 5148
rect 9456 5108 9462 5120
rect 9493 5117 9505 5120
rect 9539 5117 9551 5151
rect 9646 5148 9674 5188
rect 10594 5176 10600 5228
rect 10652 5176 10658 5228
rect 11974 5176 11980 5228
rect 12032 5216 12038 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 12032 5188 12265 5216
rect 12032 5176 12038 5188
rect 12253 5185 12265 5188
rect 12299 5216 12311 5219
rect 13464 5216 13492 5247
rect 12299 5188 13492 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9646 5120 9965 5148
rect 9493 5111 9551 5117
rect 9953 5117 9965 5120
rect 9999 5148 10011 5151
rect 10612 5148 10640 5176
rect 9999 5120 10640 5148
rect 10873 5151 10931 5157
rect 9999 5117 10011 5120
rect 9953 5111 10011 5117
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 11146 5148 11152 5160
rect 10919 5120 11152 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 11514 5148 11520 5160
rect 11475 5120 11520 5148
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 12066 5148 12072 5160
rect 11979 5120 12072 5148
rect 12066 5108 12072 5120
rect 12124 5148 12130 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12124 5120 12449 5148
rect 12124 5108 12130 5120
rect 12437 5117 12449 5120
rect 12483 5148 12495 5151
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12483 5120 12909 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 13538 5148 13544 5160
rect 13499 5120 13544 5148
rect 12897 5111 12955 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 4617 5083 4675 5089
rect 4617 5049 4629 5083
rect 4663 5049 4675 5083
rect 4617 5043 4675 5049
rect 7561 5083 7619 5089
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 8015 5083 8073 5089
rect 8015 5080 8027 5083
rect 7607 5052 8027 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 8015 5049 8027 5052
rect 8061 5080 8073 5083
rect 8110 5080 8116 5092
rect 8061 5052 8116 5080
rect 8061 5049 8073 5052
rect 8015 5043 8073 5049
rect 4632 5012 4660 5043
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 13924 5089 13952 5256
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 21450 5284 21456 5296
rect 19116 5256 21456 5284
rect 19116 5244 19122 5256
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15378 5216 15384 5228
rect 14875 5188 15384 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 19242 5216 19248 5228
rect 19155 5188 19248 5216
rect 19242 5176 19248 5188
rect 19300 5216 19306 5228
rect 19610 5216 19616 5228
rect 19300 5188 19616 5216
rect 19300 5176 19306 5188
rect 19610 5176 19616 5188
rect 19668 5176 19674 5228
rect 21100 5225 21128 5256
rect 21450 5244 21456 5256
rect 21508 5244 21514 5296
rect 21634 5284 21640 5296
rect 21595 5256 21640 5284
rect 21634 5244 21640 5256
rect 21692 5244 21698 5296
rect 24581 5287 24639 5293
rect 24581 5253 24593 5287
rect 24627 5284 24639 5287
rect 26878 5284 26884 5296
rect 24627 5256 26884 5284
rect 24627 5253 24639 5256
rect 24581 5247 24639 5253
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 33229 5287 33287 5293
rect 33229 5253 33241 5287
rect 33275 5284 33287 5287
rect 34698 5284 34704 5296
rect 33275 5256 34704 5284
rect 33275 5253 33287 5256
rect 33229 5247 33287 5253
rect 34698 5244 34704 5256
rect 34756 5284 34762 5296
rect 36265 5287 36323 5293
rect 36265 5284 36277 5287
rect 34756 5256 36277 5284
rect 34756 5244 34762 5256
rect 36265 5253 36277 5256
rect 36311 5284 36323 5287
rect 36630 5284 36636 5296
rect 36311 5256 36636 5284
rect 36311 5253 36323 5256
rect 36265 5247 36323 5253
rect 36630 5244 36636 5256
rect 36688 5244 36694 5296
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 23109 5219 23167 5225
rect 23109 5185 23121 5219
rect 23155 5216 23167 5219
rect 23474 5216 23480 5228
rect 23155 5188 23480 5216
rect 23155 5185 23167 5188
rect 23109 5179 23167 5185
rect 23474 5176 23480 5188
rect 23532 5216 23538 5228
rect 24854 5216 24860 5228
rect 23532 5188 24860 5216
rect 23532 5176 23538 5188
rect 24854 5176 24860 5188
rect 24912 5176 24918 5228
rect 26050 5216 26056 5228
rect 26011 5188 26056 5216
rect 26050 5176 26056 5188
rect 26108 5176 26114 5228
rect 26142 5176 26148 5228
rect 26200 5216 26206 5228
rect 26697 5219 26755 5225
rect 26697 5216 26709 5219
rect 26200 5188 26709 5216
rect 26200 5176 26206 5188
rect 26697 5185 26709 5188
rect 26743 5216 26755 5219
rect 26973 5219 27031 5225
rect 26743 5188 26832 5216
rect 26743 5185 26755 5188
rect 26697 5179 26755 5185
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5117 14519 5151
rect 15194 5148 15200 5160
rect 15155 5120 15200 5148
rect 14461 5111 14519 5117
rect 10965 5083 11023 5089
rect 10965 5049 10977 5083
rect 11011 5080 11023 5083
rect 11609 5083 11667 5089
rect 11609 5080 11621 5083
rect 11011 5052 11621 5080
rect 11011 5049 11023 5052
rect 10965 5043 11023 5049
rect 11609 5049 11621 5052
rect 11655 5049 11667 5083
rect 11609 5043 11667 5049
rect 13903 5083 13961 5089
rect 13903 5049 13915 5083
rect 13949 5049 13961 5083
rect 14476 5080 14504 5111
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 18046 5108 18052 5120
rect 18104 5148 18110 5160
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 18104 5120 18521 5148
rect 18104 5108 18110 5120
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 24302 5148 24308 5160
rect 23707 5120 24308 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 24302 5108 24308 5120
rect 24360 5108 24366 5160
rect 15473 5083 15531 5089
rect 14476 5052 15332 5080
rect 13903 5043 13961 5049
rect 9490 5012 9496 5024
rect 4356 4984 4660 5012
rect 9451 4984 9496 5012
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 12069 5015 12127 5021
rect 12069 5012 12081 5015
rect 10836 4984 12081 5012
rect 10836 4972 10842 4984
rect 12069 4981 12081 4984
rect 12115 4981 12127 5015
rect 15304 5012 15332 5052
rect 15473 5049 15485 5083
rect 15519 5080 15531 5083
rect 15838 5080 15844 5092
rect 15519 5052 15844 5080
rect 15519 5049 15531 5052
rect 15473 5043 15531 5049
rect 15488 5012 15516 5043
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 19153 5083 19211 5089
rect 19153 5049 19165 5083
rect 19199 5080 19211 5083
rect 19334 5080 19340 5092
rect 19199 5052 19340 5080
rect 19199 5049 19211 5052
rect 19153 5043 19211 5049
rect 19334 5040 19340 5052
rect 19392 5080 19398 5092
rect 19607 5083 19665 5089
rect 19607 5080 19619 5083
rect 19392 5052 19619 5080
rect 19392 5040 19398 5052
rect 19607 5049 19619 5052
rect 19653 5080 19665 5083
rect 19702 5080 19708 5092
rect 19653 5052 19708 5080
rect 19653 5049 19665 5052
rect 19607 5043 19665 5049
rect 19702 5040 19708 5052
rect 19760 5040 19766 5092
rect 21177 5083 21235 5089
rect 20456 5052 21036 5080
rect 15304 4984 15516 5012
rect 12069 4975 12127 4981
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 17000 4984 17325 5012
rect 17000 4972 17006 4984
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 17678 5012 17684 5024
rect 17639 4984 17684 5012
rect 17313 4975 17371 4981
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 20456 5021 20484 5052
rect 20165 5015 20223 5021
rect 20165 4981 20177 5015
rect 20211 5012 20223 5015
rect 20441 5015 20499 5021
rect 20441 5012 20453 5015
rect 20211 4984 20453 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 20441 4981 20453 4984
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 20530 4972 20536 5024
rect 20588 5012 20594 5024
rect 20809 5015 20867 5021
rect 20809 5012 20821 5015
rect 20588 4984 20821 5012
rect 20588 4972 20594 4984
rect 20809 4981 20821 4984
rect 20855 4981 20867 5015
rect 21008 5012 21036 5052
rect 21177 5049 21189 5083
rect 21223 5049 21235 5083
rect 21177 5043 21235 5049
rect 23293 5083 23351 5089
rect 23293 5049 23305 5083
rect 23339 5080 23351 5083
rect 23982 5083 24040 5089
rect 23982 5080 23994 5083
rect 23339 5052 23994 5080
rect 23339 5049 23351 5052
rect 23293 5043 23351 5049
rect 23982 5049 23994 5052
rect 24028 5080 24040 5083
rect 24394 5080 24400 5092
rect 24028 5052 24400 5080
rect 24028 5049 24040 5052
rect 23982 5043 24040 5049
rect 21192 5012 21220 5043
rect 24394 5040 24400 5052
rect 24452 5080 24458 5092
rect 24857 5083 24915 5089
rect 24857 5080 24869 5083
rect 24452 5052 24869 5080
rect 24452 5040 24458 5052
rect 24857 5049 24869 5052
rect 24903 5049 24915 5083
rect 24857 5043 24915 5049
rect 21008 4984 21220 5012
rect 20809 4975 20867 4981
rect 22278 4972 22284 5024
rect 22336 5012 22342 5024
rect 22373 5015 22431 5021
rect 22373 5012 22385 5015
rect 22336 4984 22385 5012
rect 22336 4972 22342 4984
rect 22373 4981 22385 4984
rect 22419 4981 22431 5015
rect 22554 5012 22560 5024
rect 22515 4984 22560 5012
rect 22373 4975 22431 4981
rect 22554 4972 22560 4984
rect 22612 4972 22618 5024
rect 25406 5012 25412 5024
rect 25367 4984 25412 5012
rect 25406 4972 25412 4984
rect 25464 4972 25470 5024
rect 26804 5012 26832 5188
rect 26973 5185 26985 5219
rect 27019 5216 27031 5219
rect 27062 5216 27068 5228
rect 27019 5188 27068 5216
rect 27019 5185 27031 5188
rect 26973 5179 27031 5185
rect 27062 5176 27068 5188
rect 27120 5176 27126 5228
rect 27246 5216 27252 5228
rect 27207 5188 27252 5216
rect 27246 5176 27252 5188
rect 27304 5176 27310 5228
rect 28166 5176 28172 5228
rect 28224 5216 28230 5228
rect 29641 5219 29699 5225
rect 29641 5216 29653 5219
rect 28224 5188 29653 5216
rect 28224 5176 28230 5188
rect 29641 5185 29653 5188
rect 29687 5185 29699 5219
rect 29641 5179 29699 5185
rect 31846 5176 31852 5228
rect 31904 5216 31910 5228
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 31904 5188 32321 5216
rect 31904 5176 31910 5188
rect 32309 5185 32321 5188
rect 32355 5216 32367 5219
rect 32950 5216 32956 5228
rect 32355 5188 32956 5216
rect 32355 5185 32367 5188
rect 32309 5179 32367 5185
rect 32950 5176 32956 5188
rect 33008 5176 33014 5228
rect 33965 5219 34023 5225
rect 33965 5185 33977 5219
rect 34011 5216 34023 5219
rect 34146 5216 34152 5228
rect 34011 5188 34152 5216
rect 34011 5185 34023 5188
rect 33965 5179 34023 5185
rect 30834 5148 30840 5160
rect 30795 5120 30840 5148
rect 30834 5108 30840 5120
rect 30892 5148 30898 5160
rect 31297 5151 31355 5157
rect 31297 5148 31309 5151
rect 30892 5120 31309 5148
rect 30892 5108 30898 5120
rect 31297 5117 31309 5120
rect 31343 5117 31355 5151
rect 31297 5111 31355 5117
rect 31570 5108 31576 5160
rect 31628 5148 31634 5160
rect 33505 5151 33563 5157
rect 33505 5148 33517 5151
rect 31628 5120 33517 5148
rect 31628 5108 31634 5120
rect 33505 5117 33517 5120
rect 33551 5117 33563 5151
rect 33505 5111 33563 5117
rect 27065 5083 27123 5089
rect 27065 5049 27077 5083
rect 27111 5080 27123 5083
rect 28997 5083 29055 5089
rect 28997 5080 29009 5083
rect 27111 5052 29009 5080
rect 27111 5049 27123 5052
rect 27065 5043 27123 5049
rect 28997 5049 29009 5052
rect 29043 5049 29055 5083
rect 28997 5043 29055 5049
rect 27080 5012 27108 5043
rect 26804 4984 27108 5012
rect 29012 5012 29040 5043
rect 29086 5040 29092 5092
rect 29144 5080 29150 5092
rect 29365 5083 29423 5089
rect 29365 5080 29377 5083
rect 29144 5052 29377 5080
rect 29144 5040 29150 5052
rect 29365 5049 29377 5052
rect 29411 5049 29423 5083
rect 29365 5043 29423 5049
rect 29457 5083 29515 5089
rect 29457 5049 29469 5083
rect 29503 5049 29515 5083
rect 29457 5043 29515 5049
rect 29472 5012 29500 5043
rect 30190 5040 30196 5092
rect 30248 5080 30254 5092
rect 30377 5083 30435 5089
rect 30377 5080 30389 5083
rect 30248 5052 30389 5080
rect 30248 5040 30254 5052
rect 30377 5049 30389 5052
rect 30423 5080 30435 5083
rect 31849 5083 31907 5089
rect 31849 5080 31861 5083
rect 30423 5052 31861 5080
rect 30423 5049 30435 5052
rect 30377 5043 30435 5049
rect 31849 5049 31861 5052
rect 31895 5080 31907 5083
rect 32217 5083 32275 5089
rect 32217 5080 32229 5083
rect 31895 5052 32229 5080
rect 31895 5049 31907 5052
rect 31849 5043 31907 5049
rect 32217 5049 32229 5052
rect 32263 5080 32275 5083
rect 32490 5080 32496 5092
rect 32263 5052 32496 5080
rect 32263 5049 32275 5052
rect 32217 5043 32275 5049
rect 32490 5040 32496 5052
rect 32548 5080 32554 5092
rect 32671 5083 32729 5089
rect 32671 5080 32683 5083
rect 32548 5052 32683 5080
rect 32548 5040 32554 5052
rect 32671 5049 32683 5052
rect 32717 5080 32729 5083
rect 33980 5080 34008 5179
rect 34146 5176 34152 5188
rect 34204 5176 34210 5228
rect 34977 5219 35035 5225
rect 34977 5185 34989 5219
rect 35023 5216 35035 5219
rect 35066 5216 35072 5228
rect 35023 5188 35072 5216
rect 35023 5185 35035 5188
rect 34977 5179 35035 5185
rect 35066 5176 35072 5188
rect 35124 5176 35130 5228
rect 35342 5216 35348 5228
rect 35303 5188 35348 5216
rect 35342 5176 35348 5188
rect 35400 5176 35406 5228
rect 35986 5176 35992 5228
rect 36044 5216 36050 5228
rect 36817 5219 36875 5225
rect 36817 5216 36829 5219
rect 36044 5188 36829 5216
rect 36044 5176 36050 5188
rect 36817 5185 36829 5188
rect 36863 5185 36875 5219
rect 36817 5179 36875 5185
rect 32717 5052 34008 5080
rect 32717 5049 32729 5052
rect 32671 5043 32729 5049
rect 35066 5040 35072 5092
rect 35124 5080 35130 5092
rect 35124 5052 35169 5080
rect 35124 5040 35130 5052
rect 36170 5040 36176 5092
rect 36228 5080 36234 5092
rect 36541 5083 36599 5089
rect 36541 5080 36553 5083
rect 36228 5052 36553 5080
rect 36228 5040 36234 5052
rect 36541 5049 36553 5052
rect 36587 5049 36599 5083
rect 36541 5043 36599 5049
rect 36630 5040 36636 5092
rect 36688 5080 36694 5092
rect 36688 5052 36733 5080
rect 36688 5040 36694 5052
rect 29012 4984 29500 5012
rect 30466 4972 30472 5024
rect 30524 5012 30530 5024
rect 30653 5015 30711 5021
rect 30653 5012 30665 5015
rect 30524 4984 30665 5012
rect 30524 4972 30530 4984
rect 30653 4981 30665 4984
rect 30699 4981 30711 5015
rect 30653 4975 30711 4981
rect 34701 5015 34759 5021
rect 34701 4981 34713 5015
rect 34747 5012 34759 5015
rect 35084 5012 35112 5040
rect 34747 4984 35112 5012
rect 34747 4981 34759 4984
rect 34701 4975 34759 4981
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 1946 4808 1952 4820
rect 1719 4780 1952 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6086 4808 6092 4820
rect 5859 4780 6092 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 8110 4808 8116 4820
rect 7791 4780 8116 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8110 4768 8116 4780
rect 8168 4808 8174 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 8168 4780 8217 4808
rect 8168 4768 8174 4780
rect 8205 4777 8217 4780
rect 8251 4808 8263 4811
rect 12158 4808 12164 4820
rect 8251 4780 11646 4808
rect 12119 4780 12164 4808
rect 8251 4777 8263 4780
rect 8205 4771 8263 4777
rect 2127 4743 2185 4749
rect 2127 4709 2139 4743
rect 2173 4740 2185 4743
rect 2498 4740 2504 4752
rect 2173 4712 2504 4740
rect 2173 4709 2185 4712
rect 2127 4703 2185 4709
rect 2498 4700 2504 4712
rect 2556 4700 2562 4752
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 4249 4743 4307 4749
rect 4249 4740 4261 4743
rect 4028 4712 4261 4740
rect 4028 4700 4034 4712
rect 4249 4709 4261 4712
rect 4295 4740 4307 4743
rect 5077 4743 5135 4749
rect 5077 4740 5089 4743
rect 4295 4712 5089 4740
rect 4295 4709 4307 4712
rect 4249 4703 4307 4709
rect 5077 4709 5089 4712
rect 5123 4709 5135 4743
rect 9214 4740 9220 4752
rect 5077 4703 5135 4709
rect 8772 4712 9220 4740
rect 6546 4672 6552 4684
rect 6507 4644 6552 4672
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 8478 4672 8484 4684
rect 6840 4644 8484 4672
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 3142 4604 3148 4616
rect 1811 4576 3148 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4604 3571 4607
rect 4157 4607 4215 4613
rect 4157 4604 4169 4607
rect 3559 4576 4169 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 4157 4573 4169 4576
rect 4203 4604 4215 4607
rect 6840 4604 6868 4644
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 8772 4681 8800 4712
rect 9214 4700 9220 4712
rect 9272 4740 9278 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9272 4712 9873 4740
rect 9272 4700 9278 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 9861 4703 9919 4709
rect 10134 4700 10140 4752
rect 10192 4740 10198 4752
rect 10413 4743 10471 4749
rect 10413 4740 10425 4743
rect 10192 4712 10425 4740
rect 10192 4700 10198 4712
rect 10413 4709 10425 4712
rect 10459 4740 10471 4743
rect 10962 4740 10968 4752
rect 10459 4712 10968 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11618 4749 11646 4780
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 13078 4808 13084 4820
rect 12943 4780 13084 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 13078 4768 13084 4780
rect 13136 4808 13142 4820
rect 13446 4808 13452 4820
rect 13136 4780 13452 4808
rect 13136 4768 13142 4780
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 14240 4780 14381 4808
rect 14240 4768 14246 4780
rect 14369 4777 14381 4780
rect 14415 4777 14427 4811
rect 14369 4771 14427 4777
rect 16942 4768 16948 4820
rect 17000 4808 17006 4820
rect 18049 4811 18107 4817
rect 18049 4808 18061 4811
rect 17000 4780 18061 4808
rect 17000 4768 17006 4780
rect 18049 4777 18061 4780
rect 18095 4808 18107 4811
rect 18138 4808 18144 4820
rect 18095 4780 18144 4808
rect 18095 4777 18107 4780
rect 18049 4771 18107 4777
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4808 19671 4811
rect 20530 4808 20536 4820
rect 19659 4780 20536 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 21910 4808 21916 4820
rect 21871 4780 21916 4808
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 24302 4808 24308 4820
rect 24263 4780 24308 4808
rect 24302 4768 24308 4780
rect 24360 4808 24366 4820
rect 24949 4811 25007 4817
rect 24949 4808 24961 4811
rect 24360 4780 24961 4808
rect 24360 4768 24366 4780
rect 24949 4777 24961 4780
rect 24995 4777 25007 4811
rect 24949 4771 25007 4777
rect 25958 4768 25964 4820
rect 26016 4808 26022 4820
rect 26237 4811 26295 4817
rect 26237 4808 26249 4811
rect 26016 4780 26249 4808
rect 26016 4768 26022 4780
rect 26237 4777 26249 4780
rect 26283 4777 26295 4811
rect 26237 4771 26295 4777
rect 29086 4768 29092 4820
rect 29144 4808 29150 4820
rect 29273 4811 29331 4817
rect 29273 4808 29285 4811
rect 29144 4780 29285 4808
rect 29144 4768 29150 4780
rect 29273 4777 29285 4780
rect 29319 4777 29331 4811
rect 32582 4808 32588 4820
rect 32543 4780 32588 4808
rect 29273 4771 29331 4777
rect 32582 4768 32588 4780
rect 32640 4768 32646 4820
rect 32950 4808 32956 4820
rect 32911 4780 32956 4808
rect 32950 4768 32956 4780
rect 33008 4768 33014 4820
rect 34974 4808 34980 4820
rect 34935 4780 34980 4808
rect 34974 4768 34980 4780
rect 35032 4768 35038 4820
rect 35066 4768 35072 4820
rect 35124 4808 35130 4820
rect 36081 4811 36139 4817
rect 36081 4808 36093 4811
rect 35124 4780 36093 4808
rect 35124 4768 35130 4780
rect 36081 4777 36093 4780
rect 36127 4777 36139 4811
rect 36081 4771 36139 4777
rect 36170 4768 36176 4820
rect 36228 4808 36234 4820
rect 36449 4811 36507 4817
rect 36449 4808 36461 4811
rect 36228 4780 36461 4808
rect 36228 4768 36234 4780
rect 36449 4777 36461 4780
rect 36495 4777 36507 4811
rect 36449 4771 36507 4777
rect 11603 4743 11661 4749
rect 11603 4709 11615 4743
rect 11649 4740 11661 4743
rect 11974 4740 11980 4752
rect 11649 4712 11980 4740
rect 11649 4709 11661 4712
rect 11603 4703 11661 4709
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 12452 4740 12480 4768
rect 13173 4743 13231 4749
rect 13173 4740 13185 4743
rect 12452 4712 13185 4740
rect 13173 4709 13185 4712
rect 13219 4709 13231 4743
rect 13722 4740 13728 4752
rect 13683 4712 13728 4740
rect 13173 4703 13231 4709
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 16853 4743 16911 4749
rect 16853 4740 16865 4743
rect 15948 4712 16865 4740
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4641 8815 4675
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 8757 4635 8815 4641
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 15580 4644 15853 4672
rect 4203 4576 6868 4604
rect 7009 4607 7067 4613
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 7055 4576 7297 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7285 4573 7297 4576
rect 7331 4604 7343 4607
rect 7466 4604 7472 4616
rect 7331 4576 7472 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8018 4604 8024 4616
rect 7883 4576 8024 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8018 4564 8024 4576
rect 8076 4604 8082 4616
rect 9490 4604 9496 4616
rect 8076 4576 9496 4604
rect 8076 4564 8082 4576
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9766 4604 9772 4616
rect 9727 4576 9772 4604
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11112 4576 11253 4604
rect 11112 4564 11118 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 14642 4604 14648 4616
rect 13127 4576 14648 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 15102 4564 15108 4616
rect 15160 4604 15166 4616
rect 15580 4604 15608 4644
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 15841 4635 15899 4641
rect 15160 4576 15608 4604
rect 15657 4607 15715 4613
rect 15160 4564 15166 4576
rect 15657 4573 15669 4607
rect 15703 4604 15715 4607
rect 15948 4604 15976 4712
rect 16853 4709 16865 4712
rect 16899 4740 16911 4743
rect 17494 4740 17500 4752
rect 16899 4712 17500 4740
rect 16899 4709 16911 4712
rect 16853 4703 16911 4709
rect 17494 4700 17500 4712
rect 17552 4740 17558 4752
rect 17678 4740 17684 4752
rect 17552 4712 17684 4740
rect 17552 4700 17558 4712
rect 17678 4700 17684 4712
rect 17736 4700 17742 4752
rect 19055 4743 19113 4749
rect 19055 4709 19067 4743
rect 19101 4740 19113 4743
rect 19702 4740 19708 4752
rect 19101 4712 19708 4740
rect 19101 4709 19113 4712
rect 19055 4703 19113 4709
rect 19702 4700 19708 4712
rect 19760 4700 19766 4752
rect 20717 4743 20775 4749
rect 20717 4709 20729 4743
rect 20763 4740 20775 4743
rect 20806 4740 20812 4752
rect 20763 4712 20812 4740
rect 20763 4709 20775 4712
rect 20717 4703 20775 4709
rect 20806 4700 20812 4712
rect 20864 4740 20870 4752
rect 21085 4743 21143 4749
rect 21085 4740 21097 4743
rect 20864 4712 21097 4740
rect 20864 4700 20870 4712
rect 21085 4709 21097 4712
rect 21131 4709 21143 4743
rect 21634 4740 21640 4752
rect 21595 4712 21640 4740
rect 21085 4703 21143 4709
rect 21634 4700 21640 4712
rect 21692 4700 21698 4752
rect 24026 4740 24032 4752
rect 23987 4712 24032 4740
rect 24026 4700 24032 4712
rect 24084 4740 24090 4752
rect 24673 4743 24731 4749
rect 24673 4740 24685 4743
rect 24084 4712 24685 4740
rect 24084 4700 24090 4712
rect 24673 4709 24685 4712
rect 24719 4709 24731 4743
rect 26694 4740 26700 4752
rect 26655 4712 26700 4740
rect 24673 4703 24731 4709
rect 26694 4700 26700 4712
rect 26752 4700 26758 4752
rect 28258 4740 28264 4752
rect 28219 4712 28264 4740
rect 28258 4700 28264 4712
rect 28316 4700 28322 4752
rect 33775 4743 33833 4749
rect 33775 4709 33787 4743
rect 33821 4740 33833 4743
rect 34146 4740 34152 4752
rect 33821 4712 34152 4740
rect 33821 4709 33833 4712
rect 33775 4703 33833 4709
rect 34146 4700 34152 4712
rect 34204 4740 34210 4752
rect 34882 4740 34888 4752
rect 34204 4712 34888 4740
rect 34204 4700 34210 4712
rect 34882 4700 34888 4712
rect 34940 4700 34946 4752
rect 34992 4740 35020 4768
rect 34992 4712 35388 4740
rect 18506 4632 18512 4684
rect 18564 4672 18570 4684
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 18564 4644 18705 4672
rect 18564 4632 18570 4644
rect 18693 4641 18705 4644
rect 18739 4672 18751 4675
rect 20257 4675 20315 4681
rect 20257 4672 20269 4675
rect 18739 4644 20269 4672
rect 18739 4641 18751 4644
rect 18693 4635 18751 4641
rect 20257 4641 20269 4644
rect 20303 4641 20315 4675
rect 23382 4672 23388 4684
rect 23343 4644 23388 4672
rect 20257 4635 20315 4641
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 23658 4632 23664 4684
rect 23716 4672 23722 4684
rect 23753 4675 23811 4681
rect 23753 4672 23765 4675
rect 23716 4644 23765 4672
rect 23716 4632 23722 4644
rect 23753 4641 23765 4644
rect 23799 4641 23811 4675
rect 23753 4635 23811 4641
rect 15703 4576 15976 4604
rect 16393 4607 16451 4613
rect 15703 4573 15715 4576
rect 15657 4567 15715 4573
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16666 4604 16672 4616
rect 16439 4576 16672 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16666 4564 16672 4576
rect 16724 4604 16730 4616
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 16724 4576 17233 4604
rect 16724 4564 16730 4576
rect 17221 4573 17233 4576
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4604 21051 4607
rect 21266 4604 21272 4616
rect 21039 4576 21272 4604
rect 21039 4573 21051 4576
rect 20993 4567 21051 4573
rect 21266 4564 21272 4576
rect 21324 4604 21330 4616
rect 22554 4604 22560 4616
rect 21324 4576 22560 4604
rect 21324 4564 21330 4576
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 23768 4604 23796 4635
rect 24762 4632 24768 4684
rect 24820 4672 24826 4684
rect 24857 4675 24915 4681
rect 24857 4672 24869 4675
rect 24820 4644 24869 4672
rect 24820 4632 24826 4644
rect 24857 4641 24869 4644
rect 24903 4641 24915 4675
rect 25317 4675 25375 4681
rect 25317 4672 25329 4675
rect 24857 4635 24915 4641
rect 25148 4644 25329 4672
rect 25148 4616 25176 4644
rect 25317 4641 25329 4644
rect 25363 4641 25375 4675
rect 25317 4635 25375 4641
rect 30374 4632 30380 4684
rect 30432 4672 30438 4684
rect 30469 4675 30527 4681
rect 30469 4672 30481 4675
rect 30432 4644 30481 4672
rect 30432 4632 30438 4644
rect 30469 4641 30481 4644
rect 30515 4641 30527 4675
rect 31018 4672 31024 4684
rect 30979 4644 31024 4672
rect 30469 4635 30527 4641
rect 31018 4632 31024 4644
rect 31076 4632 31082 4684
rect 31205 4675 31263 4681
rect 31205 4641 31217 4675
rect 31251 4672 31263 4675
rect 35250 4672 35256 4684
rect 31251 4644 35256 4672
rect 31251 4641 31263 4644
rect 31205 4635 31263 4641
rect 35250 4632 35256 4644
rect 35308 4632 35314 4684
rect 35360 4672 35388 4712
rect 35434 4700 35440 4752
rect 35492 4740 35498 4752
rect 35492 4712 35537 4740
rect 35492 4700 35498 4712
rect 35802 4672 35808 4684
rect 35360 4644 35808 4672
rect 35802 4632 35808 4644
rect 35860 4632 35866 4684
rect 25130 4604 25136 4616
rect 23768 4576 25136 4604
rect 25130 4564 25136 4576
rect 25188 4564 25194 4616
rect 25958 4564 25964 4616
rect 26016 4604 26022 4616
rect 26605 4607 26663 4613
rect 26605 4604 26617 4607
rect 26016 4576 26617 4604
rect 26016 4564 26022 4576
rect 26605 4573 26617 4576
rect 26651 4604 26663 4607
rect 27246 4604 27252 4616
rect 26651 4576 27252 4604
rect 26651 4573 26663 4576
rect 26605 4567 26663 4573
rect 27246 4564 27252 4576
rect 27304 4564 27310 4616
rect 28166 4604 28172 4616
rect 28127 4576 28172 4604
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 28445 4607 28503 4613
rect 28445 4573 28457 4607
rect 28491 4573 28503 4607
rect 32122 4604 32128 4616
rect 32083 4576 32128 4604
rect 28445 4567 28503 4573
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 3053 4539 3111 4545
rect 3053 4536 3065 4539
rect 2924 4508 3065 4536
rect 2924 4496 2930 4508
rect 3053 4505 3065 4508
rect 3099 4536 3111 4539
rect 4246 4536 4252 4548
rect 3099 4508 4252 4536
rect 3099 4505 3111 4508
rect 3053 4499 3111 4505
rect 4246 4496 4252 4508
rect 4304 4496 4310 4548
rect 4706 4536 4712 4548
rect 4619 4508 4712 4536
rect 4706 4496 4712 4508
rect 4764 4536 4770 4548
rect 4764 4508 9076 4536
rect 4764 4496 4770 4508
rect 9048 4480 9076 4508
rect 11146 4496 11152 4548
rect 11204 4536 11210 4548
rect 17954 4536 17960 4548
rect 11204 4508 17960 4536
rect 11204 4496 11210 4508
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 23014 4496 23020 4548
rect 23072 4536 23078 4548
rect 23290 4536 23296 4548
rect 23072 4508 23296 4536
rect 23072 4496 23078 4508
rect 23290 4496 23296 4508
rect 23348 4496 23354 4548
rect 27154 4536 27160 4548
rect 27115 4508 27160 4536
rect 27154 4496 27160 4508
rect 27212 4536 27218 4548
rect 28460 4536 28488 4567
rect 32122 4564 32128 4576
rect 32180 4564 32186 4616
rect 33413 4607 33471 4613
rect 33413 4573 33425 4607
rect 33459 4604 33471 4607
rect 33962 4604 33968 4616
rect 33459 4576 33968 4604
rect 33459 4573 33471 4576
rect 33413 4567 33471 4573
rect 33962 4564 33968 4576
rect 34020 4564 34026 4616
rect 35158 4604 35164 4616
rect 35119 4576 35164 4604
rect 35158 4564 35164 4576
rect 35216 4564 35222 4616
rect 28810 4536 28816 4548
rect 27212 4508 28816 4536
rect 27212 4496 27218 4508
rect 28810 4496 28816 4508
rect 28868 4496 28874 4548
rect 2685 4471 2743 4477
rect 2685 4437 2697 4471
rect 2731 4468 2743 4471
rect 2774 4468 2780 4480
rect 2731 4440 2780 4468
rect 2731 4437 2743 4440
rect 2685 4431 2743 4437
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 9030 4468 9036 4480
rect 8991 4440 9036 4468
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 9398 4468 9404 4480
rect 9359 4440 9404 4468
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4468 10931 4471
rect 10962 4468 10968 4480
rect 10919 4440 10968 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 13814 4468 13820 4480
rect 13044 4440 13820 4468
rect 13044 4428 13050 4440
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 15105 4471 15163 4477
rect 15105 4437 15117 4471
rect 15151 4468 15163 4471
rect 15194 4468 15200 4480
rect 15151 4440 15200 4468
rect 15151 4437 15163 4440
rect 15105 4431 15163 4437
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 16482 4428 16488 4480
rect 16540 4468 16546 4480
rect 16669 4471 16727 4477
rect 16669 4468 16681 4471
rect 16540 4440 16681 4468
rect 16540 4428 16546 4440
rect 16669 4437 16681 4440
rect 16715 4468 16727 4471
rect 16942 4468 16948 4480
rect 16715 4440 16948 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16942 4428 16948 4440
rect 17000 4477 17006 4480
rect 17000 4471 17049 4477
rect 17000 4437 17003 4471
rect 17037 4437 17049 4471
rect 17126 4468 17132 4480
rect 17087 4440 17132 4468
rect 17000 4431 17049 4437
rect 17000 4428 17006 4431
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 17310 4468 17316 4480
rect 17271 4440 17316 4468
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 18322 4428 18328 4480
rect 18380 4468 18386 4480
rect 18417 4471 18475 4477
rect 18417 4468 18429 4471
rect 18380 4440 18429 4468
rect 18380 4428 18386 4440
rect 18417 4437 18429 4440
rect 18463 4437 18475 4471
rect 18417 4431 18475 4437
rect 19150 4428 19156 4480
rect 19208 4468 19214 4480
rect 19889 4471 19947 4477
rect 19889 4468 19901 4471
rect 19208 4440 19901 4468
rect 19208 4428 19214 4440
rect 19889 4437 19901 4440
rect 19935 4437 19947 4471
rect 31478 4468 31484 4480
rect 31439 4440 31484 4468
rect 19889 4431 19947 4437
rect 31478 4428 31484 4440
rect 31536 4428 31542 4480
rect 34333 4471 34391 4477
rect 34333 4437 34345 4471
rect 34379 4468 34391 4471
rect 34606 4468 34612 4480
rect 34379 4440 34612 4468
rect 34379 4437 34391 4440
rect 34333 4431 34391 4437
rect 34606 4428 34612 4440
rect 34664 4428 34670 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 2498 4264 2504 4276
rect 2459 4236 2504 4264
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 4706 4264 4712 4276
rect 3252 4236 4712 4264
rect 2133 4199 2191 4205
rect 2133 4196 2145 4199
rect 2043 4168 2145 4196
rect 2133 4165 2145 4168
rect 2179 4196 2191 4199
rect 2314 4196 2320 4208
rect 2179 4168 2320 4196
rect 2179 4165 2191 4168
rect 2133 4159 2191 4165
rect 1486 4060 1492 4072
rect 1447 4032 1492 4060
rect 1486 4020 1492 4032
rect 1544 4060 1550 4072
rect 2148 4060 2176 4159
rect 2314 4156 2320 4168
rect 2372 4156 2378 4208
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 3252 4205 3280 4236
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 5537 4267 5595 4273
rect 5537 4233 5549 4267
rect 5583 4264 5595 4267
rect 6365 4267 6423 4273
rect 5583 4236 6316 4264
rect 5583 4233 5595 4236
rect 5537 4227 5595 4233
rect 3237 4199 3295 4205
rect 3237 4196 3249 4199
rect 2924 4168 3249 4196
rect 2924 4156 2930 4168
rect 3237 4165 3249 4168
rect 3283 4165 3295 4199
rect 3970 4196 3976 4208
rect 3931 4168 3976 4196
rect 3237 4159 3295 4165
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 5626 4156 5632 4208
rect 5684 4196 5690 4208
rect 5810 4196 5816 4208
rect 5684 4168 5816 4196
rect 5684 4156 5690 4168
rect 5810 4156 5816 4168
rect 5868 4196 5874 4208
rect 5905 4199 5963 4205
rect 5905 4196 5917 4199
rect 5868 4168 5917 4196
rect 5868 4156 5874 4168
rect 5905 4165 5917 4168
rect 5951 4165 5963 4199
rect 6288 4196 6316 4236
rect 6365 4233 6377 4267
rect 6411 4264 6423 4267
rect 6730 4264 6736 4276
rect 6411 4236 6736 4264
rect 6411 4233 6423 4236
rect 6365 4227 6423 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 6822 4224 6828 4276
rect 6880 4264 6886 4276
rect 7009 4267 7067 4273
rect 7009 4264 7021 4267
rect 6880 4236 7021 4264
rect 6880 4224 6886 4236
rect 7009 4233 7021 4236
rect 7055 4233 7067 4267
rect 9214 4264 9220 4276
rect 9175 4236 9220 4264
rect 7009 4227 7067 4233
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 11514 4224 11520 4276
rect 11572 4264 11578 4276
rect 15746 4264 15752 4276
rect 11572 4236 15752 4264
rect 11572 4224 11578 4236
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 16577 4267 16635 4273
rect 16577 4264 16589 4267
rect 16172 4236 16589 4264
rect 16172 4224 16178 4236
rect 16577 4233 16589 4236
rect 16623 4264 16635 4267
rect 17126 4264 17132 4276
rect 16623 4236 17132 4264
rect 16623 4233 16635 4236
rect 16577 4227 16635 4233
rect 17126 4224 17132 4236
rect 17184 4264 17190 4276
rect 17313 4267 17371 4273
rect 17313 4264 17325 4267
rect 17184 4236 17325 4264
rect 17184 4224 17190 4236
rect 17313 4233 17325 4236
rect 17359 4233 17371 4267
rect 17313 4227 17371 4233
rect 18138 4224 18144 4276
rect 18196 4273 18202 4276
rect 18196 4267 18245 4273
rect 18196 4233 18199 4267
rect 18233 4233 18245 4267
rect 18196 4227 18245 4233
rect 19153 4267 19211 4273
rect 19153 4233 19165 4267
rect 19199 4264 19211 4267
rect 19702 4264 19708 4276
rect 19199 4236 19708 4264
rect 19199 4233 19211 4236
rect 19153 4227 19211 4233
rect 18196 4224 18202 4227
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 21266 4264 21272 4276
rect 21227 4236 21272 4264
rect 20901 4227 20959 4233
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 23017 4267 23075 4273
rect 23017 4233 23029 4267
rect 23063 4264 23075 4267
rect 23382 4264 23388 4276
rect 23063 4236 23388 4264
rect 23063 4233 23075 4236
rect 23017 4227 23075 4233
rect 23382 4224 23388 4236
rect 23440 4264 23446 4276
rect 23658 4264 23664 4276
rect 23440 4236 23664 4264
rect 23440 4224 23446 4236
rect 23658 4224 23664 4236
rect 23716 4224 23722 4276
rect 24394 4224 24400 4276
rect 24452 4264 24458 4276
rect 24765 4267 24823 4273
rect 24765 4264 24777 4267
rect 24452 4236 24777 4264
rect 24452 4224 24458 4236
rect 24765 4233 24777 4236
rect 24811 4233 24823 4267
rect 24765 4227 24823 4233
rect 25869 4267 25927 4273
rect 25869 4233 25881 4267
rect 25915 4264 25927 4267
rect 26234 4264 26240 4276
rect 25915 4236 26240 4264
rect 25915 4233 25927 4236
rect 25869 4227 25927 4233
rect 6546 4196 6552 4208
rect 6288 4168 6552 4196
rect 5905 4159 5963 4165
rect 6546 4156 6552 4168
rect 6604 4196 6610 4208
rect 9858 4196 9864 4208
rect 6604 4168 9864 4196
rect 6604 4156 6610 4168
rect 9858 4156 9864 4168
rect 9916 4196 9922 4208
rect 10226 4196 10232 4208
rect 9916 4168 10232 4196
rect 9916 4156 9922 4168
rect 10226 4156 10232 4168
rect 10284 4156 10290 4208
rect 11330 4196 11336 4208
rect 11291 4168 11336 4196
rect 11330 4156 11336 4168
rect 11388 4156 11394 4208
rect 11885 4199 11943 4205
rect 11885 4165 11897 4199
rect 11931 4196 11943 4199
rect 11974 4196 11980 4208
rect 11931 4168 11980 4196
rect 11931 4165 11943 4168
rect 11885 4159 11943 4165
rect 11974 4156 11980 4168
rect 12032 4156 12038 4208
rect 12710 4196 12716 4208
rect 12671 4168 12716 4196
rect 12710 4156 12716 4168
rect 12768 4196 12774 4208
rect 13814 4196 13820 4208
rect 12768 4168 13820 4196
rect 12768 4156 12774 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 16482 4205 16488 4208
rect 16466 4199 16488 4205
rect 16466 4165 16478 4199
rect 16466 4159 16488 4165
rect 16482 4156 16488 4159
rect 16540 4156 16546 4208
rect 17862 4156 17868 4208
rect 17920 4196 17926 4208
rect 18322 4196 18328 4208
rect 17920 4168 18328 4196
rect 17920 4156 17926 4168
rect 18322 4156 18328 4168
rect 18380 4196 18386 4208
rect 18380 4168 18644 4196
rect 18380 4156 18386 4168
rect 2682 4128 2688 4140
rect 2643 4100 2688 4128
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 3936 4100 4261 4128
rect 3936 4088 3942 4100
rect 4249 4097 4261 4100
rect 4295 4128 4307 4131
rect 5442 4128 5448 4140
rect 4295 4100 5448 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7524 4100 7849 4128
rect 7524 4088 7530 4100
rect 7837 4097 7849 4100
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 16298 4128 16304 4140
rect 13136 4100 16304 4128
rect 13136 4088 13142 4100
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 16666 4088 16672 4100
rect 16724 4128 16730 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 16724 4100 17785 4128
rect 16724 4088 16730 4100
rect 17773 4097 17785 4100
rect 17819 4128 17831 4131
rect 18417 4131 18475 4137
rect 18417 4128 18429 4131
rect 17819 4100 18429 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 18417 4097 18429 4100
rect 18463 4097 18475 4131
rect 18417 4091 18475 4097
rect 1544 4032 2176 4060
rect 5721 4063 5779 4069
rect 1544 4020 1550 4032
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6086 4060 6092 4072
rect 5767 4032 6092 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 6871 4032 7389 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7377 4029 7389 4032
rect 7423 4060 7435 4063
rect 9674 4060 9680 4072
rect 7423 4032 9680 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 9999 4032 10701 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10689 4029 10701 4032
rect 10735 4060 10747 4063
rect 10962 4060 10968 4072
rect 10735 4032 10968 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 11425 4063 11483 4069
rect 11425 4029 11437 4063
rect 11471 4029 11483 4063
rect 11425 4023 11483 4029
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4060 13231 4063
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 13219 4032 13553 4060
rect 13219 4029 13231 4032
rect 13173 4023 13231 4029
rect 13541 4029 13553 4032
rect 13587 4060 13599 4063
rect 13630 4060 13636 4072
rect 13587 4032 13636 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 2774 3992 2780 4004
rect 2735 3964 2780 3992
rect 2774 3952 2780 3964
rect 2832 3992 2838 4004
rect 3605 3995 3663 4001
rect 3605 3992 3617 3995
rect 2832 3964 3617 3992
rect 2832 3952 2838 3964
rect 3605 3961 3617 3964
rect 3651 3992 3663 3995
rect 4341 3995 4399 4001
rect 3651 3964 4154 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 1719 3927 1777 3933
rect 1719 3893 1731 3927
rect 1765 3924 1777 3927
rect 2222 3924 2228 3936
rect 1765 3896 2228 3924
rect 1765 3893 1777 3896
rect 1719 3887 1777 3893
rect 2222 3884 2228 3896
rect 2280 3884 2286 3936
rect 4126 3924 4154 3964
rect 4341 3961 4353 3995
rect 4387 3961 4399 3995
rect 4890 3992 4896 4004
rect 4803 3964 4896 3992
rect 4341 3955 4399 3961
rect 4356 3924 4384 3955
rect 4890 3952 4896 3964
rect 4948 3992 4954 4004
rect 7745 3995 7803 4001
rect 4948 3964 5764 3992
rect 4948 3952 4954 3964
rect 5258 3924 5264 3936
rect 4126 3896 4384 3924
rect 5219 3896 5264 3924
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 5736 3924 5764 3964
rect 7745 3961 7757 3995
rect 7791 3992 7803 3995
rect 7926 3992 7932 4004
rect 7791 3964 7932 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 7926 3952 7932 3964
rect 7984 3992 7990 4004
rect 8110 3992 8116 4004
rect 7984 3964 8116 3992
rect 7984 3952 7990 3964
rect 8110 3952 8116 3964
rect 8168 4001 8174 4004
rect 8168 3995 8216 4001
rect 8168 3961 8170 3995
rect 8204 3961 8216 3995
rect 8168 3955 8216 3961
rect 9585 3995 9643 4001
rect 9585 3961 9597 3995
rect 9631 3992 9643 3995
rect 11054 3992 11060 4004
rect 9631 3964 11060 3992
rect 9631 3961 9643 3964
rect 9585 3955 9643 3961
rect 8168 3952 8174 3955
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 8294 3924 8300 3936
rect 5736 3896 8300 3924
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8754 3924 8760 3936
rect 8715 3896 8760 3924
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 10321 3927 10379 3933
rect 10321 3893 10333 3927
rect 10367 3924 10379 3927
rect 10502 3924 10508 3936
rect 10367 3896 10508 3924
rect 10367 3893 10379 3896
rect 10321 3887 10379 3893
rect 10502 3884 10508 3896
rect 10560 3924 10566 3936
rect 11256 3924 11284 4023
rect 11440 3992 11468 4023
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 13906 4069 13912 4072
rect 13863 4063 13912 4069
rect 13863 4029 13875 4063
rect 13909 4029 13912 4063
rect 13863 4023 13912 4029
rect 13906 4020 13912 4023
rect 13964 4060 13970 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13964 4032 14289 4060
rect 13964 4020 13970 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 15102 4060 15108 4072
rect 15063 4032 15108 4060
rect 14277 4023 14335 4029
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 15252 4032 15485 4060
rect 15252 4020 15258 4032
rect 15473 4029 15485 4032
rect 15519 4060 15531 4063
rect 15654 4060 15660 4072
rect 15519 4032 15660 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 15654 4020 15660 4032
rect 15712 4060 15718 4072
rect 17037 4063 17095 4069
rect 15712 4032 16344 4060
rect 15712 4020 15718 4032
rect 11790 3992 11796 4004
rect 11440 3964 11796 3992
rect 11790 3952 11796 3964
rect 11848 3992 11854 4004
rect 14642 3992 14648 4004
rect 11848 3964 14648 3992
rect 11848 3952 11854 3964
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 14829 3995 14887 4001
rect 14829 3961 14841 3995
rect 14875 3992 14887 3995
rect 14918 3992 14924 4004
rect 14875 3964 14924 3992
rect 14875 3961 14887 3964
rect 14829 3955 14887 3961
rect 14918 3952 14924 3964
rect 14976 3992 14982 4004
rect 15286 3992 15292 4004
rect 14976 3964 15292 3992
rect 14976 3952 14982 3964
rect 15286 3952 15292 3964
rect 15344 3992 15350 4004
rect 16316 4001 16344 4032
rect 17037 4029 17049 4063
rect 17083 4060 17095 4063
rect 18138 4060 18144 4072
rect 17083 4032 18144 4060
rect 17083 4029 17095 4032
rect 17037 4023 17095 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 18616 4060 18644 4168
rect 21358 4156 21364 4208
rect 21416 4196 21422 4208
rect 21545 4199 21603 4205
rect 21545 4196 21557 4199
rect 21416 4168 21557 4196
rect 21416 4156 21422 4168
rect 21545 4165 21557 4168
rect 21591 4196 21603 4199
rect 22278 4196 22284 4208
rect 21591 4168 22284 4196
rect 21591 4165 21603 4168
rect 21545 4159 21603 4165
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 23198 4156 23204 4208
rect 23256 4196 23262 4208
rect 23293 4199 23351 4205
rect 23293 4196 23305 4199
rect 23256 4168 23305 4196
rect 23256 4156 23262 4168
rect 23293 4165 23305 4168
rect 23339 4165 23351 4199
rect 23293 4159 23351 4165
rect 24489 4199 24547 4205
rect 24489 4165 24501 4199
rect 24535 4196 24547 4199
rect 24670 4196 24676 4208
rect 24535 4168 24676 4196
rect 24535 4165 24547 4168
rect 24489 4159 24547 4165
rect 24670 4156 24676 4168
rect 24728 4156 24734 4208
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4128 18843 4131
rect 21082 4128 21088 4140
rect 18831 4100 21088 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 19429 4063 19487 4069
rect 19429 4060 19441 4063
rect 18616 4032 19441 4060
rect 19429 4029 19441 4032
rect 19475 4029 19487 4063
rect 19429 4023 19487 4029
rect 19886 4020 19892 4072
rect 19944 4060 19950 4072
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19944 4032 19993 4060
rect 19944 4020 19950 4032
rect 19981 4029 19993 4032
rect 20027 4060 20039 4063
rect 20622 4060 20628 4072
rect 20027 4032 20628 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 21726 4060 21732 4072
rect 21687 4032 21732 4060
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 22278 4060 22284 4072
rect 22239 4032 22284 4060
rect 22278 4020 22284 4032
rect 22336 4020 22342 4072
rect 15749 3995 15807 4001
rect 15749 3992 15761 3995
rect 15344 3964 15761 3992
rect 15344 3952 15350 3964
rect 15749 3961 15761 3964
rect 15795 3961 15807 3995
rect 15749 3955 15807 3961
rect 16301 3995 16359 4001
rect 16301 3961 16313 3995
rect 16347 3992 16359 3995
rect 16574 3992 16580 4004
rect 16347 3964 16580 3992
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 17494 3952 17500 4004
rect 17552 3992 17558 4004
rect 18049 3995 18107 4001
rect 18049 3992 18061 3995
rect 17552 3964 18061 3992
rect 17552 3952 17558 3964
rect 18049 3961 18061 3964
rect 18095 3961 18107 3995
rect 20302 3995 20360 4001
rect 20302 3992 20314 3995
rect 18049 3955 18107 3961
rect 19812 3964 20314 3992
rect 10560 3896 11284 3924
rect 12253 3927 12311 3933
rect 10560 3884 10566 3896
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 12986 3924 12992 3936
rect 12299 3896 12992 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13538 3924 13544 3936
rect 13499 3896 13544 3924
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 19702 3884 19708 3936
rect 19760 3924 19766 3936
rect 19812 3933 19840 3964
rect 20302 3961 20314 3964
rect 20348 3961 20360 3995
rect 24780 3992 24808 4227
rect 26234 4224 26240 4236
rect 26292 4264 26298 4276
rect 26694 4264 26700 4276
rect 26292 4236 26700 4264
rect 26292 4224 26298 4236
rect 26694 4224 26700 4236
rect 26752 4224 26758 4276
rect 27617 4267 27675 4273
rect 27617 4233 27629 4267
rect 27663 4264 27675 4267
rect 28169 4267 28227 4273
rect 28169 4264 28181 4267
rect 27663 4236 28181 4264
rect 27663 4233 27675 4236
rect 27617 4227 27675 4233
rect 28169 4233 28181 4236
rect 28215 4264 28227 4267
rect 28258 4264 28264 4276
rect 28215 4236 28264 4264
rect 28215 4233 28227 4236
rect 28169 4227 28227 4233
rect 28258 4224 28264 4236
rect 28316 4224 28322 4276
rect 30929 4267 30987 4273
rect 30929 4233 30941 4267
rect 30975 4264 30987 4267
rect 31018 4264 31024 4276
rect 30975 4236 31024 4264
rect 30975 4233 30987 4236
rect 30929 4227 30987 4233
rect 31018 4224 31024 4236
rect 31076 4264 31082 4276
rect 32401 4267 32459 4273
rect 32401 4264 32413 4267
rect 31076 4236 32413 4264
rect 31076 4224 31082 4236
rect 32401 4233 32413 4236
rect 32447 4233 32459 4267
rect 34606 4264 34612 4276
rect 32401 4227 32459 4233
rect 33152 4236 34514 4264
rect 34567 4236 34612 4264
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 30374 4196 30380 4208
rect 24912 4168 30380 4196
rect 24912 4156 24918 4168
rect 30374 4156 30380 4168
rect 30432 4196 30438 4208
rect 30469 4199 30527 4205
rect 30469 4196 30481 4199
rect 30432 4168 30481 4196
rect 30432 4156 30438 4168
rect 30469 4165 30481 4168
rect 30515 4165 30527 4199
rect 31202 4196 31208 4208
rect 30469 4159 30527 4165
rect 30944 4168 31208 4196
rect 26513 4131 26571 4137
rect 26513 4128 26525 4131
rect 25285 4100 26525 4128
rect 24946 4060 24952 4072
rect 24907 4032 24952 4060
rect 24946 4020 24952 4032
rect 25004 4020 25010 4072
rect 25285 4001 25313 4100
rect 26513 4097 26525 4100
rect 26559 4128 26571 4131
rect 26559 4100 27108 4128
rect 26559 4097 26571 4100
rect 26513 4091 26571 4097
rect 26697 4063 26755 4069
rect 26697 4060 26709 4063
rect 26160 4032 26709 4060
rect 25270 3995 25328 4001
rect 25270 3992 25282 3995
rect 24780 3964 25282 3992
rect 20302 3955 20360 3961
rect 25270 3961 25282 3964
rect 25316 3961 25328 3995
rect 25270 3955 25328 3961
rect 26160 3936 26188 4032
rect 26697 4029 26709 4032
rect 26743 4029 26755 4063
rect 26697 4023 26755 4029
rect 27080 4001 27108 4100
rect 28902 4088 28908 4140
rect 28960 4128 28966 4140
rect 29546 4128 29552 4140
rect 28960 4100 29552 4128
rect 28960 4088 28966 4100
rect 29546 4088 29552 4100
rect 29604 4088 29610 4140
rect 29362 4060 29368 4072
rect 29323 4032 29368 4060
rect 29362 4020 29368 4032
rect 29420 4020 29426 4072
rect 29825 4063 29883 4069
rect 29825 4029 29837 4063
rect 29871 4060 29883 4063
rect 30944 4060 30972 4168
rect 31202 4156 31208 4168
rect 31260 4156 31266 4208
rect 31113 4131 31171 4137
rect 31113 4097 31125 4131
rect 31159 4128 31171 4131
rect 31386 4128 31392 4140
rect 31159 4100 31392 4128
rect 31159 4097 31171 4100
rect 31113 4091 31171 4097
rect 31386 4088 31392 4100
rect 31444 4088 31450 4140
rect 32416 4128 32444 4227
rect 32600 4168 32720 4196
rect 32600 4128 32628 4168
rect 32416 4100 32628 4128
rect 32582 4060 32588 4072
rect 29871 4032 30972 4060
rect 32543 4032 32588 4060
rect 29871 4029 29883 4032
rect 29825 4023 29883 4029
rect 27059 3995 27117 4001
rect 27059 3961 27071 3995
rect 27105 3992 27117 3995
rect 28350 3992 28356 4004
rect 27105 3964 28356 3992
rect 27105 3961 27117 3964
rect 27059 3955 27117 3961
rect 28350 3952 28356 3964
rect 28408 3952 28414 4004
rect 29840 3992 29868 4023
rect 32582 4020 32588 4032
rect 32640 4020 32646 4072
rect 32692 4060 32720 4168
rect 33045 4063 33103 4069
rect 33045 4060 33057 4063
rect 32692 4032 33057 4060
rect 33045 4029 33057 4032
rect 33091 4029 33103 4063
rect 33045 4023 33103 4029
rect 30098 3992 30104 4004
rect 29012 3964 29868 3992
rect 30059 3964 30104 3992
rect 29012 3936 29040 3964
rect 30098 3952 30104 3964
rect 30156 3952 30162 4004
rect 31205 3995 31263 4001
rect 31205 3961 31217 3995
rect 31251 3992 31263 3995
rect 31478 3992 31484 4004
rect 31251 3964 31484 3992
rect 31251 3961 31263 3964
rect 31205 3955 31263 3961
rect 31478 3952 31484 3964
rect 31536 3952 31542 4004
rect 31757 3995 31815 4001
rect 31757 3961 31769 3995
rect 31803 3992 31815 3995
rect 33152 3992 33180 4236
rect 33594 4156 33600 4208
rect 33652 4196 33658 4208
rect 33689 4199 33747 4205
rect 33689 4196 33701 4199
rect 33652 4168 33701 4196
rect 33652 4156 33658 4168
rect 33689 4165 33701 4168
rect 33735 4196 33747 4199
rect 34146 4196 34152 4208
rect 33735 4168 34152 4196
rect 33735 4165 33747 4168
rect 33689 4159 33747 4165
rect 34146 4156 34152 4168
rect 34204 4156 34210 4208
rect 34486 4196 34514 4236
rect 34606 4224 34612 4236
rect 34664 4224 34670 4276
rect 34882 4224 34888 4276
rect 34940 4264 34946 4276
rect 35434 4264 35440 4276
rect 34940 4236 35440 4264
rect 34940 4224 34946 4236
rect 35434 4224 35440 4236
rect 35492 4264 35498 4276
rect 35897 4267 35955 4273
rect 35897 4264 35909 4267
rect 35492 4236 35909 4264
rect 35492 4224 35498 4236
rect 35897 4233 35909 4236
rect 35943 4233 35955 4267
rect 35897 4227 35955 4233
rect 35986 4224 35992 4276
rect 36044 4264 36050 4276
rect 36265 4267 36323 4273
rect 36265 4264 36277 4267
rect 36044 4236 36277 4264
rect 36044 4224 36050 4236
rect 36265 4233 36277 4236
rect 36311 4233 36323 4267
rect 36265 4227 36323 4233
rect 36633 4267 36691 4273
rect 36633 4233 36645 4267
rect 36679 4264 36691 4267
rect 36722 4264 36728 4276
rect 36679 4236 36728 4264
rect 36679 4233 36691 4236
rect 36633 4227 36691 4233
rect 36722 4224 36728 4236
rect 36780 4224 36786 4276
rect 35342 4196 35348 4208
rect 34486 4168 35348 4196
rect 35342 4156 35348 4168
rect 35400 4196 35406 4208
rect 35529 4199 35587 4205
rect 35529 4196 35541 4199
rect 35400 4168 35541 4196
rect 35400 4156 35406 4168
rect 35529 4165 35541 4168
rect 35575 4165 35587 4199
rect 35529 4159 35587 4165
rect 34977 4131 35035 4137
rect 34977 4097 34989 4131
rect 35023 4128 35035 4131
rect 36004 4128 36032 4224
rect 35023 4100 36032 4128
rect 35023 4097 35035 4100
rect 34977 4091 35035 4097
rect 36446 4060 36452 4072
rect 36407 4032 36452 4060
rect 36446 4020 36452 4032
rect 36504 4060 36510 4072
rect 36998 4060 37004 4072
rect 36504 4032 37004 4060
rect 36504 4020 36510 4032
rect 36998 4020 37004 4032
rect 37056 4020 37062 4072
rect 37366 4020 37372 4072
rect 37424 4060 37430 4072
rect 37588 4063 37646 4069
rect 37588 4060 37600 4063
rect 37424 4032 37600 4060
rect 37424 4020 37430 4032
rect 37588 4029 37600 4032
rect 37634 4060 37646 4063
rect 38013 4063 38071 4069
rect 38013 4060 38025 4063
rect 37634 4032 38025 4060
rect 37634 4029 37646 4032
rect 37588 4023 37646 4029
rect 38013 4029 38025 4032
rect 38059 4029 38071 4063
rect 38013 4023 38071 4029
rect 33318 3992 33324 4004
rect 31803 3964 33180 3992
rect 33279 3964 33324 3992
rect 31803 3961 31815 3964
rect 31757 3955 31815 3961
rect 19797 3927 19855 3933
rect 19797 3924 19809 3927
rect 19760 3896 19809 3924
rect 19760 3884 19766 3896
rect 19797 3893 19809 3896
rect 19843 3893 19855 3927
rect 22002 3924 22008 3936
rect 21963 3896 22008 3924
rect 19797 3887 19855 3893
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 23658 3924 23664 3936
rect 23619 3896 23664 3924
rect 23658 3884 23664 3896
rect 23716 3884 23722 3936
rect 26142 3924 26148 3936
rect 26103 3896 26148 3924
rect 26142 3884 26148 3896
rect 26200 3884 26206 3936
rect 27338 3884 27344 3936
rect 27396 3924 27402 3936
rect 28166 3924 28172 3936
rect 27396 3896 28172 3924
rect 27396 3884 27402 3896
rect 28166 3884 28172 3896
rect 28224 3924 28230 3936
rect 28445 3927 28503 3933
rect 28445 3924 28457 3927
rect 28224 3896 28457 3924
rect 28224 3884 28230 3896
rect 28445 3893 28457 3896
rect 28491 3893 28503 3927
rect 28994 3924 29000 3936
rect 28955 3896 29000 3924
rect 28445 3887 28503 3893
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 29086 3884 29092 3936
rect 29144 3924 29150 3936
rect 31772 3924 31800 3955
rect 33318 3952 33324 3964
rect 33376 3952 33382 4004
rect 35069 3995 35127 4001
rect 35069 3961 35081 3995
rect 35115 3961 35127 3995
rect 35069 3955 35127 3961
rect 29144 3896 31800 3924
rect 29144 3884 29150 3896
rect 33134 3884 33140 3936
rect 33192 3924 33198 3936
rect 33962 3924 33968 3936
rect 33192 3896 33968 3924
rect 33192 3884 33198 3896
rect 33962 3884 33968 3896
rect 34020 3884 34026 3936
rect 34606 3884 34612 3936
rect 34664 3924 34670 3936
rect 35084 3924 35112 3955
rect 35434 3952 35440 4004
rect 35492 3992 35498 4004
rect 37691 3995 37749 4001
rect 37691 3992 37703 3995
rect 35492 3964 37703 3992
rect 35492 3952 35498 3964
rect 37691 3961 37703 3964
rect 37737 3961 37749 3995
rect 37691 3955 37749 3961
rect 34664 3896 35112 3924
rect 34664 3884 34670 3896
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 2774 3720 2780 3732
rect 2735 3692 2780 3720
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3142 3720 3148 3732
rect 3103 3692 3148 3720
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4157 3723 4215 3729
rect 4157 3689 4169 3723
rect 4203 3689 4215 3723
rect 4157 3683 4215 3689
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 1943 3655 2001 3661
rect 1943 3652 1955 3655
rect 1728 3624 1955 3652
rect 1728 3612 1734 3624
rect 1943 3621 1955 3624
rect 1989 3652 2001 3655
rect 2498 3652 2504 3664
rect 1989 3624 2504 3652
rect 1989 3621 2001 3624
rect 1943 3615 2001 3621
rect 2498 3612 2504 3624
rect 2556 3612 2562 3664
rect 3160 3652 3188 3680
rect 4172 3652 4200 3683
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 4304 3692 5733 3720
rect 4304 3680 4310 3692
rect 5721 3689 5733 3692
rect 5767 3689 5779 3723
rect 5721 3683 5779 3689
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 6917 3723 6975 3729
rect 6917 3720 6929 3723
rect 6788 3692 6929 3720
rect 6788 3680 6794 3692
rect 6917 3689 6929 3692
rect 6963 3689 6975 3723
rect 6917 3683 6975 3689
rect 7561 3723 7619 3729
rect 7561 3689 7573 3723
rect 7607 3720 7619 3723
rect 8018 3720 8024 3732
rect 7607 3692 8024 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8352 3692 9137 3720
rect 8352 3680 8358 3692
rect 9125 3689 9137 3692
rect 9171 3720 9183 3723
rect 9214 3720 9220 3732
rect 9171 3692 9220 3720
rect 9171 3689 9183 3692
rect 9125 3683 9183 3689
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 9858 3720 9864 3732
rect 9819 3692 9864 3720
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 11054 3720 11060 3732
rect 11015 3692 11060 3720
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 11940 3692 13461 3720
rect 11940 3680 11946 3692
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13449 3683 13507 3689
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 13998 3720 14004 3732
rect 13688 3692 14004 3720
rect 13688 3680 13694 3692
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 14093 3723 14151 3729
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 14277 3723 14335 3729
rect 14277 3720 14289 3723
rect 14139 3692 14289 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14277 3689 14289 3692
rect 14323 3720 14335 3723
rect 18322 3720 18328 3732
rect 14323 3692 18328 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 18322 3680 18328 3692
rect 18380 3680 18386 3732
rect 18966 3720 18972 3732
rect 18927 3692 18972 3720
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 20806 3720 20812 3732
rect 19576 3692 20812 3720
rect 19576 3680 19582 3692
rect 20806 3680 20812 3692
rect 20864 3720 20870 3732
rect 20864 3692 21128 3720
rect 20864 3680 20870 3692
rect 6362 3652 6368 3664
rect 3160 3624 4200 3652
rect 5736 3624 6368 3652
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3752 3556 4077 3584
rect 3752 3544 3758 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4614 3584 4620 3596
rect 4575 3556 4620 3584
rect 4065 3547 4123 3553
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 4080 3516 4108 3547
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5736 3593 5764 3624
rect 6362 3612 6368 3624
rect 6420 3652 6426 3664
rect 6822 3652 6828 3664
rect 6420 3624 6828 3652
rect 6420 3612 6426 3624
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8205 3655 8263 3661
rect 8205 3652 8217 3655
rect 8168 3624 8217 3652
rect 8168 3612 8174 3624
rect 8205 3621 8217 3624
rect 8251 3652 8263 3655
rect 8754 3652 8760 3664
rect 8251 3624 8760 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 12986 3612 12992 3664
rect 13044 3612 13050 3664
rect 13078 3612 13084 3664
rect 13136 3612 13142 3664
rect 13814 3652 13820 3664
rect 13775 3624 13820 3652
rect 13814 3612 13820 3624
rect 13872 3652 13878 3664
rect 16393 3655 16451 3661
rect 13872 3624 15792 3652
rect 13872 3612 13878 3624
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3553 5779 3587
rect 5721 3547 5779 3553
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 6270 3584 6276 3596
rect 6227 3556 6276 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 6270 3544 6276 3556
rect 6328 3584 6334 3596
rect 6730 3584 6736 3596
rect 6328 3556 6736 3584
rect 6328 3544 6334 3556
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9640 3556 9689 3584
rect 9640 3544 9646 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 11054 3584 11060 3596
rect 11015 3556 11060 3584
rect 9677 3547 9735 3553
rect 11054 3544 11060 3556
rect 11112 3544 11118 3596
rect 11606 3584 11612 3596
rect 11567 3556 11612 3584
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11790 3584 11796 3596
rect 11751 3556 11796 3584
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 12802 3584 12808 3596
rect 12763 3556 12808 3584
rect 12802 3544 12808 3556
rect 12860 3584 12866 3596
rect 13004 3584 13032 3612
rect 12860 3556 13032 3584
rect 12860 3544 12866 3556
rect 5810 3516 5816 3528
rect 4080 3488 5816 3516
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 9030 3516 9036 3528
rect 8159 3488 9036 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10870 3516 10876 3528
rect 10551 3488 10876 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 11808 3516 11836 3544
rect 10928 3488 11836 3516
rect 12952 3519 13010 3525
rect 10928 3476 10934 3488
rect 12952 3485 12964 3519
rect 12998 3516 13010 3519
rect 13096 3516 13124 3612
rect 13906 3584 13912 3596
rect 13188 3556 13912 3584
rect 13188 3528 13216 3556
rect 13906 3544 13912 3556
rect 13964 3584 13970 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13964 3556 14105 3584
rect 13964 3544 13970 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 15654 3584 15660 3596
rect 15615 3556 15660 3584
rect 14093 3547 14151 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 15764 3584 15792 3624
rect 16393 3621 16405 3655
rect 16439 3652 16451 3655
rect 18046 3652 18052 3664
rect 16439 3624 18052 3652
rect 16439 3621 16451 3624
rect 16393 3615 16451 3621
rect 18046 3612 18052 3624
rect 18104 3612 18110 3664
rect 18230 3652 18236 3664
rect 18191 3624 18236 3652
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 19886 3652 19892 3664
rect 19847 3624 19892 3652
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 20901 3655 20959 3661
rect 20901 3621 20913 3655
rect 20947 3652 20959 3655
rect 20947 3624 21036 3652
rect 20947 3621 20959 3624
rect 20901 3615 20959 3621
rect 15887 3587 15945 3593
rect 15887 3584 15899 3587
rect 15764 3556 15899 3584
rect 15887 3553 15899 3556
rect 15933 3584 15945 3587
rect 17037 3587 17095 3593
rect 17037 3584 17049 3587
rect 15933 3556 17049 3584
rect 15933 3553 15945 3556
rect 15887 3547 15945 3553
rect 17037 3553 17049 3556
rect 17083 3553 17095 3587
rect 17037 3547 17095 3553
rect 17221 3587 17279 3593
rect 17221 3553 17233 3587
rect 17267 3584 17279 3587
rect 18248 3584 18276 3612
rect 17267 3556 18276 3584
rect 17267 3553 17279 3556
rect 17221 3547 17279 3553
rect 18966 3544 18972 3596
rect 19024 3584 19030 3596
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 19024 3556 19165 3584
rect 19024 3544 19030 3556
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 19610 3584 19616 3596
rect 19571 3556 19616 3584
rect 19153 3547 19211 3553
rect 19610 3544 19616 3556
rect 19668 3544 19674 3596
rect 12998 3488 13124 3516
rect 12998 3485 13010 3488
rect 12952 3479 13010 3485
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13228 3488 13273 3516
rect 13228 3476 13234 3488
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 14700 3488 16037 3516
rect 14700 3476 14706 3488
rect 16025 3485 16037 3488
rect 16071 3516 16083 3519
rect 16666 3516 16672 3528
rect 16071 3488 16672 3516
rect 16071 3485 16083 3488
rect 16025 3479 16083 3485
rect 16666 3476 16672 3488
rect 16724 3516 16730 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16724 3488 16865 3516
rect 16724 3476 16730 3488
rect 16853 3485 16865 3488
rect 16899 3516 16911 3519
rect 17126 3516 17132 3528
rect 16899 3488 17132 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 17126 3476 17132 3488
rect 17184 3516 17190 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17184 3488 17601 3516
rect 17184 3476 17190 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 21008 3516 21036 3624
rect 21100 3593 21128 3692
rect 22002 3680 22008 3732
rect 22060 3720 22066 3732
rect 22189 3723 22247 3729
rect 22189 3720 22201 3723
rect 22060 3692 22201 3720
rect 22060 3680 22066 3692
rect 22189 3689 22201 3692
rect 22235 3720 22247 3723
rect 22738 3720 22744 3732
rect 22235 3692 22416 3720
rect 22699 3692 22744 3720
rect 22235 3689 22247 3692
rect 22189 3683 22247 3689
rect 22388 3593 22416 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 23293 3723 23351 3729
rect 23293 3689 23305 3723
rect 23339 3720 23351 3723
rect 23474 3720 23480 3732
rect 23339 3692 23480 3720
rect 23339 3689 23351 3692
rect 23293 3683 23351 3689
rect 23474 3680 23480 3692
rect 23532 3720 23538 3732
rect 25130 3720 25136 3732
rect 23532 3692 24348 3720
rect 25091 3692 25136 3720
rect 23532 3680 23538 3692
rect 23658 3612 23664 3664
rect 23716 3652 23722 3664
rect 24210 3652 24216 3664
rect 23716 3624 24216 3652
rect 23716 3612 23722 3624
rect 24210 3612 24216 3624
rect 24268 3612 24274 3664
rect 24320 3661 24348 3692
rect 25130 3680 25136 3692
rect 25188 3680 25194 3732
rect 25958 3720 25964 3732
rect 25919 3692 25964 3720
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 26234 3720 26240 3732
rect 26195 3692 26240 3720
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 28074 3720 28080 3732
rect 27987 3692 28080 3720
rect 28074 3680 28080 3692
rect 28132 3720 28138 3732
rect 29086 3720 29092 3732
rect 28132 3692 29092 3720
rect 28132 3680 28138 3692
rect 29086 3680 29092 3692
rect 29144 3680 29150 3732
rect 30098 3720 30104 3732
rect 30059 3692 30104 3720
rect 30098 3680 30104 3692
rect 30156 3720 30162 3732
rect 31113 3723 31171 3729
rect 30156 3692 30236 3720
rect 30156 3680 30162 3692
rect 24305 3655 24363 3661
rect 24305 3621 24317 3655
rect 24351 3621 24363 3655
rect 24305 3615 24363 3621
rect 26050 3612 26056 3664
rect 26108 3652 26114 3664
rect 26789 3655 26847 3661
rect 26789 3652 26801 3655
rect 26108 3624 26801 3652
rect 26108 3612 26114 3624
rect 26789 3621 26801 3624
rect 26835 3652 26847 3655
rect 26878 3652 26884 3664
rect 26835 3624 26884 3652
rect 26835 3621 26847 3624
rect 26789 3615 26847 3621
rect 26878 3612 26884 3624
rect 26936 3612 26942 3664
rect 27338 3652 27344 3664
rect 27299 3624 27344 3652
rect 27338 3612 27344 3624
rect 27396 3612 27402 3664
rect 28350 3612 28356 3664
rect 28408 3652 28414 3664
rect 28490 3655 28548 3661
rect 28490 3652 28502 3655
rect 28408 3624 28502 3652
rect 28408 3612 28414 3624
rect 28490 3621 28502 3624
rect 28536 3621 28548 3655
rect 28490 3615 28548 3621
rect 30208 3593 30236 3692
rect 31113 3689 31125 3723
rect 31159 3720 31171 3723
rect 31478 3720 31484 3732
rect 31159 3692 31484 3720
rect 31159 3689 31171 3692
rect 31113 3683 31171 3689
rect 31478 3680 31484 3692
rect 31536 3680 31542 3732
rect 34609 3723 34667 3729
rect 34609 3689 34621 3723
rect 34655 3720 34667 3723
rect 34655 3692 35664 3720
rect 34655 3689 34667 3692
rect 34609 3683 34667 3689
rect 30514 3655 30572 3661
rect 30514 3652 30526 3655
rect 30300 3624 30526 3652
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3553 21143 3587
rect 21085 3547 21143 3553
rect 22373 3587 22431 3593
rect 22373 3553 22385 3587
rect 22419 3553 22431 3587
rect 22373 3547 22431 3553
rect 30193 3587 30251 3593
rect 30193 3553 30205 3587
rect 30239 3553 30251 3587
rect 30193 3547 30251 3553
rect 21266 3516 21272 3528
rect 18003 3488 20944 3516
rect 21008 3488 21272 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 8665 3451 8723 3457
rect 8665 3417 8677 3451
rect 8711 3448 8723 3451
rect 10134 3448 10140 3460
rect 8711 3420 10140 3448
rect 8711 3417 8723 3420
rect 8665 3411 8723 3417
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 12618 3408 12624 3460
rect 12676 3448 12682 3460
rect 15795 3451 15853 3457
rect 15795 3448 15807 3451
rect 12676 3420 15807 3448
rect 12676 3408 12682 3420
rect 15795 3417 15807 3420
rect 15841 3448 15853 3451
rect 16482 3448 16488 3460
rect 15841 3420 16488 3448
rect 15841 3417 15853 3420
rect 15795 3411 15853 3417
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 17037 3451 17095 3457
rect 17037 3417 17049 3451
rect 17083 3448 17095 3451
rect 17497 3451 17555 3457
rect 17497 3448 17509 3451
rect 17083 3420 17509 3448
rect 17083 3417 17095 3420
rect 17037 3411 17095 3417
rect 17497 3417 17509 3420
rect 17543 3448 17555 3451
rect 17862 3448 17868 3460
rect 17543 3420 17868 3448
rect 17543 3417 17555 3420
rect 17497 3411 17555 3417
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 20165 3451 20223 3457
rect 20165 3448 20177 3451
rect 18064 3420 20177 3448
rect 18064 3392 18092 3420
rect 20165 3417 20177 3420
rect 20211 3448 20223 3451
rect 20533 3451 20591 3457
rect 20533 3448 20545 3451
rect 20211 3420 20545 3448
rect 20211 3417 20223 3420
rect 20165 3411 20223 3417
rect 20533 3417 20545 3420
rect 20579 3417 20591 3451
rect 20916 3448 20944 3488
rect 21266 3476 21272 3488
rect 21324 3476 21330 3528
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 24394 3516 24400 3528
rect 21499 3488 24400 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 24489 3519 24547 3525
rect 24489 3485 24501 3519
rect 24535 3485 24547 3519
rect 24489 3479 24547 3485
rect 23106 3448 23112 3460
rect 20916 3420 23112 3448
rect 20533 3411 20591 3417
rect 23106 3408 23112 3420
rect 23164 3408 23170 3460
rect 24118 3408 24124 3460
rect 24176 3448 24182 3460
rect 24504 3448 24532 3479
rect 26326 3476 26332 3528
rect 26384 3516 26390 3528
rect 26697 3519 26755 3525
rect 26697 3516 26709 3519
rect 26384 3488 26709 3516
rect 26384 3476 26390 3488
rect 26697 3485 26709 3488
rect 26743 3516 26755 3519
rect 26786 3516 26792 3528
rect 26743 3488 26792 3516
rect 26743 3485 26755 3488
rect 26697 3479 26755 3485
rect 26786 3476 26792 3488
rect 26844 3476 26850 3528
rect 28166 3516 28172 3528
rect 28127 3488 28172 3516
rect 28166 3476 28172 3488
rect 28224 3476 28230 3528
rect 25406 3448 25412 3460
rect 24176 3420 25412 3448
rect 24176 3408 24182 3420
rect 25406 3408 25412 3420
rect 25464 3408 25470 3460
rect 29089 3451 29147 3457
rect 29089 3417 29101 3451
rect 29135 3448 29147 3451
rect 29454 3448 29460 3460
rect 29135 3420 29460 3448
rect 29135 3417 29147 3420
rect 29089 3411 29147 3417
rect 29454 3408 29460 3420
rect 29512 3408 29518 3460
rect 30190 3408 30196 3460
rect 30248 3448 30254 3460
rect 30300 3448 30328 3624
rect 30514 3621 30526 3624
rect 30560 3621 30572 3655
rect 30514 3615 30572 3621
rect 31202 3612 31208 3664
rect 31260 3652 31266 3664
rect 31260 3624 32628 3652
rect 31260 3612 31266 3624
rect 30374 3544 30380 3596
rect 30432 3584 30438 3596
rect 31846 3584 31852 3596
rect 30432 3556 31852 3584
rect 30432 3544 30438 3556
rect 31846 3544 31852 3556
rect 31904 3584 31910 3596
rect 32600 3593 32628 3624
rect 33594 3612 33600 3664
rect 33652 3652 33658 3664
rect 35636 3661 35664 3692
rect 34010 3655 34068 3661
rect 34010 3652 34022 3655
rect 33652 3624 34022 3652
rect 33652 3612 33658 3624
rect 34010 3621 34022 3624
rect 34056 3621 34068 3655
rect 34010 3615 34068 3621
rect 35621 3655 35679 3661
rect 35621 3621 35633 3655
rect 35667 3652 35679 3655
rect 36262 3652 36268 3664
rect 35667 3624 36268 3652
rect 35667 3621 35679 3624
rect 35621 3615 35679 3621
rect 36262 3612 36268 3624
rect 36320 3612 36326 3664
rect 32125 3587 32183 3593
rect 32125 3584 32137 3587
rect 31904 3556 32137 3584
rect 31904 3544 31910 3556
rect 32125 3553 32137 3556
rect 32171 3553 32183 3587
rect 32125 3547 32183 3553
rect 32585 3587 32643 3593
rect 32585 3553 32597 3587
rect 32631 3553 32643 3587
rect 32585 3547 32643 3553
rect 33318 3544 33324 3596
rect 33376 3584 33382 3596
rect 33689 3587 33747 3593
rect 33689 3584 33701 3587
rect 33376 3556 33701 3584
rect 33376 3544 33382 3556
rect 33689 3553 33701 3556
rect 33735 3553 33747 3587
rect 33689 3547 33747 3553
rect 32861 3519 32919 3525
rect 32861 3485 32873 3519
rect 32907 3516 32919 3519
rect 35158 3516 35164 3528
rect 32907 3488 35164 3516
rect 32907 3485 32919 3488
rect 32861 3479 32919 3485
rect 35158 3476 35164 3488
rect 35216 3476 35222 3528
rect 35529 3519 35587 3525
rect 35529 3485 35541 3519
rect 35575 3516 35587 3519
rect 35894 3516 35900 3528
rect 35575 3488 35900 3516
rect 35575 3485 35587 3488
rect 35529 3479 35587 3485
rect 35894 3476 35900 3488
rect 35952 3476 35958 3528
rect 30248 3420 30328 3448
rect 30248 3408 30254 3420
rect 35618 3408 35624 3460
rect 35676 3448 35682 3460
rect 36081 3451 36139 3457
rect 36081 3448 36093 3451
rect 35676 3420 36093 3448
rect 35676 3408 35682 3420
rect 36081 3417 36093 3420
rect 36127 3417 36139 3451
rect 36081 3411 36139 3417
rect 2498 3380 2504 3392
rect 2459 3352 2504 3380
rect 2498 3340 2504 3352
rect 2556 3340 2562 3392
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 5261 3383 5319 3389
rect 5261 3380 5273 3383
rect 5132 3352 5273 3380
rect 5132 3340 5138 3352
rect 5261 3349 5273 3352
rect 5307 3380 5319 3383
rect 5442 3380 5448 3392
rect 5307 3352 5448 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 7929 3383 7987 3389
rect 7929 3349 7941 3383
rect 7975 3380 7987 3383
rect 8018 3380 8024 3392
rect 7975 3352 8024 3380
rect 7975 3349 7987 3352
rect 7929 3343 7987 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 12526 3380 12532 3392
rect 12487 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 13081 3383 13139 3389
rect 13081 3349 13093 3383
rect 13127 3380 13139 3383
rect 13814 3380 13820 3392
rect 13127 3352 13820 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 14734 3380 14740 3392
rect 14691 3352 14740 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 15013 3383 15071 3389
rect 15013 3349 15025 3383
rect 15059 3380 15071 3383
rect 15102 3380 15108 3392
rect 15059 3352 15108 3380
rect 15059 3349 15071 3352
rect 15013 3343 15071 3349
rect 15102 3340 15108 3352
rect 15160 3380 15166 3392
rect 15562 3380 15568 3392
rect 15160 3352 15568 3380
rect 15160 3340 15166 3352
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 17359 3383 17417 3389
rect 17359 3380 17371 3383
rect 16356 3352 17371 3380
rect 16356 3340 16362 3352
rect 17359 3349 17371 3352
rect 17405 3380 17417 3383
rect 18046 3380 18052 3392
rect 17405 3352 18052 3380
rect 17405 3349 17417 3352
rect 17359 3343 17417 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18322 3340 18328 3392
rect 18380 3380 18386 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18380 3352 18613 3380
rect 18380 3340 18386 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 21726 3380 21732 3392
rect 21687 3352 21732 3380
rect 18601 3343 18659 3349
rect 21726 3340 21732 3352
rect 21784 3340 21790 3392
rect 24394 3340 24400 3392
rect 24452 3380 24458 3392
rect 24946 3380 24952 3392
rect 24452 3352 24952 3380
rect 24452 3340 24458 3352
rect 24946 3340 24952 3352
rect 25004 3380 25010 3392
rect 25501 3383 25559 3389
rect 25501 3380 25513 3383
rect 25004 3352 25513 3380
rect 25004 3340 25010 3352
rect 25501 3349 25513 3352
rect 25547 3349 25559 3383
rect 25501 3343 25559 3349
rect 27430 3340 27436 3392
rect 27488 3380 27494 3392
rect 29362 3380 29368 3392
rect 27488 3352 29368 3380
rect 27488 3340 27494 3352
rect 29362 3340 29368 3352
rect 29420 3340 29426 3392
rect 31478 3380 31484 3392
rect 31439 3352 31484 3380
rect 31478 3340 31484 3352
rect 31536 3340 31542 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 3694 3176 3700 3188
rect 3655 3148 3700 3176
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 4614 3176 4620 3188
rect 4111 3148 4620 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 4614 3136 4620 3148
rect 4672 3176 4678 3188
rect 6270 3176 6276 3188
rect 4672 3148 6276 3176
rect 4672 3136 4678 3148
rect 6270 3136 6276 3148
rect 6328 3176 6334 3188
rect 8110 3176 8116 3188
rect 6328 3148 6960 3176
rect 8071 3148 8116 3176
rect 6328 3136 6334 3148
rect 3145 3111 3203 3117
rect 3145 3108 3157 3111
rect 2240 3080 3157 3108
rect 1762 3000 1768 3052
rect 1820 3040 1826 3052
rect 2240 3049 2268 3080
rect 3145 3077 3157 3080
rect 3191 3077 3203 3111
rect 3145 3071 3203 3077
rect 3234 3068 3240 3120
rect 3292 3108 3298 3120
rect 4341 3111 4399 3117
rect 4341 3108 4353 3111
rect 3292 3080 4353 3108
rect 3292 3068 3298 3080
rect 4341 3077 4353 3080
rect 4387 3108 4399 3111
rect 4387 3080 6684 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1820 3012 2237 3040
rect 1820 3000 1826 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2225 3003 2283 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 5074 3040 5080 3052
rect 4987 3012 5080 3040
rect 5074 3000 5080 3012
rect 5132 3040 5138 3052
rect 5718 3040 5724 3052
rect 5132 3012 5724 3040
rect 5132 3000 5138 3012
rect 5184 2981 5212 3012
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 5169 2975 5227 2981
rect 4203 2944 4752 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 2317 2907 2375 2913
rect 2317 2873 2329 2907
rect 2363 2904 2375 2907
rect 2498 2904 2504 2916
rect 2363 2876 2504 2904
rect 2363 2873 2375 2876
rect 2317 2867 2375 2873
rect 2038 2836 2044 2848
rect 1951 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2836 2102 2848
rect 2332 2836 2360 2867
rect 2498 2864 2504 2876
rect 2556 2864 2562 2916
rect 4724 2848 4752 2944
rect 5169 2941 5181 2975
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 5442 2972 5448 2984
rect 5316 2944 5361 2972
rect 5403 2944 5448 2972
rect 5316 2932 5322 2944
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 6656 2981 6684 3080
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6687 2944 6837 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6932 2972 6960 3148
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9548 3148 9873 3176
rect 9548 3136 9554 3148
rect 9861 3145 9873 3148
rect 9907 3176 9919 3179
rect 9950 3176 9956 3188
rect 9907 3148 9956 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10502 3176 10508 3188
rect 10463 3148 10508 3176
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12710 3176 12716 3188
rect 12299 3148 12716 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 13449 3179 13507 3185
rect 13449 3176 13461 3179
rect 13228 3148 13461 3176
rect 13228 3136 13234 3148
rect 13449 3145 13461 3148
rect 13495 3145 13507 3179
rect 13449 3139 13507 3145
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 16172 3148 17785 3176
rect 16172 3136 16178 3148
rect 17773 3145 17785 3148
rect 17819 3176 17831 3179
rect 17819 3148 18184 3176
rect 17819 3145 17831 3148
rect 17773 3139 17831 3145
rect 8938 3068 8944 3120
rect 8996 3108 9002 3120
rect 13262 3108 13268 3120
rect 8996 3080 13268 3108
rect 8996 3068 9002 3080
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 13780 3080 14105 3108
rect 13780 3068 13786 3080
rect 14093 3077 14105 3080
rect 14139 3108 14151 3111
rect 15194 3108 15200 3120
rect 14139 3080 15200 3108
rect 14139 3077 14151 3080
rect 14093 3071 14151 3077
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 16482 3068 16488 3120
rect 16540 3108 16546 3120
rect 16577 3111 16635 3117
rect 16577 3108 16589 3111
rect 16540 3080 16589 3108
rect 16540 3068 16546 3080
rect 16577 3077 16589 3080
rect 16623 3077 16635 3111
rect 16577 3071 16635 3077
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 18156 3117 18184 3148
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 20901 3179 20959 3185
rect 20901 3176 20913 3179
rect 20864 3148 20913 3176
rect 20864 3136 20870 3148
rect 20901 3145 20913 3148
rect 20947 3145 20959 3179
rect 21266 3176 21272 3188
rect 21227 3148 21272 3176
rect 20901 3139 20959 3145
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 21818 3176 21824 3188
rect 21779 3148 21824 3176
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 22738 3136 22744 3188
rect 22796 3176 22802 3188
rect 23017 3179 23075 3185
rect 23017 3176 23029 3179
rect 22796 3148 23029 3176
rect 22796 3136 22802 3148
rect 23017 3145 23029 3148
rect 23063 3145 23075 3179
rect 23017 3139 23075 3145
rect 17221 3111 17279 3117
rect 17221 3108 17233 3111
rect 17184 3080 17233 3108
rect 17184 3068 17190 3080
rect 17221 3077 17233 3080
rect 17267 3077 17279 3111
rect 17221 3071 17279 3077
rect 18141 3111 18199 3117
rect 18141 3077 18153 3111
rect 18187 3077 18199 3111
rect 23032 3108 23060 3139
rect 23474 3136 23480 3188
rect 23532 3176 23538 3188
rect 24210 3176 24216 3188
rect 23532 3148 23577 3176
rect 24171 3148 24216 3176
rect 23532 3136 23538 3148
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 26050 3176 26056 3188
rect 26011 3148 26056 3176
rect 26050 3136 26056 3148
rect 26108 3136 26114 3188
rect 28350 3136 28356 3188
rect 28408 3176 28414 3188
rect 28629 3179 28687 3185
rect 28629 3176 28641 3179
rect 28408 3148 28641 3176
rect 28408 3136 28414 3148
rect 28629 3145 28641 3148
rect 28675 3176 28687 3179
rect 30190 3176 30196 3188
rect 28675 3148 30196 3176
rect 28675 3145 28687 3148
rect 28629 3139 28687 3145
rect 30190 3136 30196 3148
rect 30248 3136 30254 3188
rect 30282 3136 30288 3188
rect 30340 3176 30346 3188
rect 30653 3179 30711 3185
rect 30653 3176 30665 3179
rect 30340 3148 30665 3176
rect 30340 3136 30346 3148
rect 30653 3145 30665 3148
rect 30699 3145 30711 3179
rect 31846 3176 31852 3188
rect 31807 3148 31852 3176
rect 30653 3139 30711 3145
rect 24489 3111 24547 3117
rect 24489 3108 24501 3111
rect 23032 3080 24501 3108
rect 18141 3071 18199 3077
rect 24489 3077 24501 3080
rect 24535 3108 24547 3111
rect 24581 3111 24639 3117
rect 24581 3108 24593 3111
rect 24535 3080 24593 3108
rect 24535 3077 24547 3080
rect 24489 3071 24547 3077
rect 24581 3077 24593 3080
rect 24627 3077 24639 3111
rect 27154 3108 27160 3120
rect 27115 3080 27160 3108
rect 24581 3071 24639 3077
rect 27154 3068 27160 3080
rect 27212 3068 27218 3120
rect 30208 3108 30236 3136
rect 30377 3111 30435 3117
rect 30377 3108 30389 3111
rect 30208 3080 30389 3108
rect 30377 3077 30389 3080
rect 30423 3077 30435 3111
rect 30377 3071 30435 3077
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3040 10287 3043
rect 11425 3043 11483 3049
rect 11425 3040 11437 3043
rect 10275 3012 11437 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 11425 3009 11437 3012
rect 11471 3040 11483 3043
rect 11606 3040 11612 3052
rect 11471 3012 11612 3040
rect 11471 3009 11483 3012
rect 11425 3003 11483 3009
rect 11606 3000 11612 3012
rect 11664 3040 11670 3052
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11664 3012 11897 3040
rect 11664 3000 11670 3012
rect 11885 3009 11897 3012
rect 11931 3040 11943 3043
rect 16022 3040 16028 3052
rect 11931 3012 13814 3040
rect 15983 3012 16028 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6932 2944 7297 2972
rect 6825 2935 6883 2941
rect 7285 2941 7297 2944
rect 7331 2972 7343 2975
rect 7926 2972 7932 2984
rect 7331 2944 7932 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8846 2972 8852 2984
rect 8527 2944 8852 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 8846 2932 8852 2944
rect 8904 2972 8910 2984
rect 8941 2975 8999 2981
rect 8941 2972 8953 2975
rect 8904 2944 8953 2972
rect 8904 2932 8910 2944
rect 8941 2941 8953 2944
rect 8987 2941 8999 2975
rect 8941 2935 8999 2941
rect 10502 2932 10508 2984
rect 10560 2972 10566 2984
rect 12452 2981 12480 3012
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 10560 2944 10793 2972
rect 10560 2932 10566 2944
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 12584 2944 12629 2972
rect 12584 2932 12590 2944
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13786 2972 13814 3012
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 16816 3012 18521 3040
rect 16816 3000 16822 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 19610 3000 19616 3052
rect 19668 3040 19674 3052
rect 23753 3043 23811 3049
rect 19668 3012 20116 3040
rect 19668 3000 19674 3012
rect 13998 2972 14004 2984
rect 12768 2944 12861 2972
rect 13786 2944 14004 2972
rect 12768 2932 12774 2944
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14240 2944 14289 2972
rect 14240 2932 14246 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 14792 2944 15577 2972
rect 14792 2932 14798 2944
rect 15565 2941 15577 2944
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 15841 2975 15899 2981
rect 15712 2944 15757 2972
rect 15712 2932 15718 2944
rect 15841 2941 15853 2975
rect 15887 2941 15899 2975
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 15841 2935 15899 2941
rect 5905 2907 5963 2913
rect 5905 2873 5917 2907
rect 5951 2904 5963 2907
rect 9490 2904 9496 2916
rect 5951 2876 9496 2904
rect 5951 2873 5963 2876
rect 5905 2867 5963 2873
rect 9490 2864 9496 2876
rect 9548 2864 9554 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 12728 2904 12756 2932
rect 15381 2907 15439 2913
rect 15381 2904 15393 2907
rect 9732 2876 12664 2904
rect 12728 2876 15393 2904
rect 9732 2864 9738 2876
rect 4706 2836 4712 2848
rect 2096 2808 2360 2836
rect 4667 2808 4712 2836
rect 2096 2796 2102 2808
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 6917 2839 6975 2845
rect 6917 2836 6929 2839
rect 6328 2808 6929 2836
rect 6328 2796 6334 2808
rect 6917 2805 6929 2808
rect 6963 2805 6975 2839
rect 6917 2799 6975 2805
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 8076 2808 8861 2836
rect 8076 2796 8082 2808
rect 8849 2805 8861 2808
rect 8895 2836 8907 2839
rect 9309 2839 9367 2845
rect 9309 2836 9321 2839
rect 8895 2808 9321 2836
rect 8895 2805 8907 2808
rect 8849 2799 8907 2805
rect 9309 2805 9321 2808
rect 9355 2805 9367 2839
rect 12636 2836 12664 2876
rect 15381 2873 15393 2876
rect 15427 2904 15439 2907
rect 15856 2904 15884 2935
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18322 2972 18328 2984
rect 18283 2944 18328 2972
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 20088 2981 20116 3012
rect 23753 3009 23765 3043
rect 23799 3040 23811 3043
rect 26329 3043 26387 3049
rect 26329 3040 26341 3043
rect 23799 3012 26341 3040
rect 23799 3009 23811 3012
rect 23753 3003 23811 3009
rect 26329 3009 26341 3012
rect 26375 3040 26387 3043
rect 26605 3043 26663 3049
rect 26605 3040 26617 3043
rect 26375 3012 26617 3040
rect 26375 3009 26387 3012
rect 26329 3003 26387 3009
rect 26605 3009 26617 3012
rect 26651 3009 26663 3043
rect 30006 3040 30012 3052
rect 29967 3012 30012 3040
rect 26605 3003 26663 3009
rect 30006 3000 30012 3012
rect 30064 3000 30070 3052
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 20073 2975 20131 2981
rect 20073 2941 20085 2975
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 22005 2975 22063 2981
rect 22005 2941 22017 2975
rect 22051 2941 22063 2975
rect 22005 2935 22063 2941
rect 22557 2975 22615 2981
rect 22557 2941 22569 2975
rect 22603 2972 22615 2975
rect 23382 2972 23388 2984
rect 22603 2944 23388 2972
rect 22603 2941 22615 2944
rect 22557 2935 22615 2941
rect 15427 2876 15884 2904
rect 15427 2873 15439 2876
rect 15381 2867 15439 2873
rect 17770 2864 17776 2916
rect 17828 2904 17834 2916
rect 19061 2907 19119 2913
rect 19061 2904 19073 2907
rect 17828 2876 19073 2904
rect 17828 2864 17834 2876
rect 19061 2873 19073 2876
rect 19107 2904 19119 2907
rect 19429 2907 19487 2913
rect 19429 2904 19441 2907
rect 19107 2876 19441 2904
rect 19107 2873 19119 2876
rect 19061 2867 19119 2873
rect 19429 2873 19441 2876
rect 19475 2904 19487 2907
rect 19610 2904 19616 2916
rect 19475 2876 19616 2904
rect 19475 2873 19487 2876
rect 19429 2867 19487 2873
rect 19610 2864 19616 2876
rect 19668 2864 19674 2916
rect 19794 2864 19800 2916
rect 19852 2904 19858 2916
rect 19904 2904 19932 2935
rect 21818 2904 21824 2916
rect 19852 2876 21824 2904
rect 19852 2864 19858 2876
rect 21818 2864 21824 2876
rect 21876 2904 21882 2916
rect 22020 2904 22048 2935
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 24762 2972 24768 2984
rect 24723 2944 24768 2972
rect 24762 2932 24768 2944
rect 24820 2932 24826 2984
rect 28074 2932 28080 2984
rect 28132 2972 28138 2984
rect 28204 2975 28262 2981
rect 28204 2972 28216 2975
rect 28132 2944 28216 2972
rect 28132 2932 28138 2944
rect 28204 2941 28216 2944
rect 28250 2941 28262 2975
rect 30668 2972 30696 3139
rect 31846 3136 31852 3148
rect 31904 3136 31910 3188
rect 32306 3176 32312 3188
rect 32267 3148 32312 3176
rect 32306 3136 32312 3148
rect 32364 3136 32370 3188
rect 33318 3136 33324 3188
rect 33376 3176 33382 3188
rect 34057 3179 34115 3185
rect 34057 3176 34069 3179
rect 33376 3148 34069 3176
rect 33376 3136 33382 3148
rect 34057 3145 34069 3148
rect 34103 3145 34115 3179
rect 34698 3176 34704 3188
rect 34659 3148 34704 3176
rect 34057 3139 34115 3145
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 35894 3176 35900 3188
rect 35855 3148 35900 3176
rect 35894 3136 35900 3148
rect 35952 3136 35958 3188
rect 36262 3176 36268 3188
rect 36223 3148 36268 3176
rect 36262 3136 36268 3148
rect 36320 3136 36326 3188
rect 33594 3068 33600 3120
rect 33652 3108 33658 3120
rect 33689 3111 33747 3117
rect 33689 3108 33701 3111
rect 33652 3080 33701 3108
rect 33652 3068 33658 3080
rect 33689 3077 33701 3080
rect 33735 3077 33747 3111
rect 33689 3071 33747 3077
rect 33778 3068 33784 3120
rect 33836 3108 33842 3120
rect 35713 3111 35771 3117
rect 35713 3108 35725 3111
rect 33836 3080 35725 3108
rect 33836 3068 33842 3080
rect 35713 3077 35725 3080
rect 35759 3077 35771 3111
rect 35713 3071 35771 3077
rect 31570 3040 31576 3052
rect 31531 3012 31576 3040
rect 31570 3000 31576 3012
rect 31628 3000 31634 3052
rect 33134 3000 33140 3052
rect 33192 3040 33198 3052
rect 34974 3040 34980 3052
rect 33192 3012 33237 3040
rect 34887 3012 34980 3040
rect 33192 3000 33198 3012
rect 34974 3000 34980 3012
rect 35032 3040 35038 3052
rect 35434 3040 35440 3052
rect 35032 3012 35440 3040
rect 35032 3000 35038 3012
rect 35434 3000 35440 3012
rect 35492 3000 35498 3052
rect 35621 3043 35679 3049
rect 35621 3009 35633 3043
rect 35667 3040 35679 3043
rect 35802 3040 35808 3052
rect 35667 3012 35808 3040
rect 35667 3009 35679 3012
rect 35621 3003 35679 3009
rect 35802 3000 35808 3012
rect 35860 3000 35866 3052
rect 35912 3040 35940 3136
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 35912 3012 36461 3040
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 30837 2975 30895 2981
rect 30837 2972 30849 2975
rect 30668 2944 30849 2972
rect 28204 2935 28262 2941
rect 30837 2941 30849 2944
rect 30883 2941 30895 2975
rect 30837 2935 30895 2941
rect 31202 2932 31208 2984
rect 31260 2972 31266 2984
rect 31297 2975 31355 2981
rect 31297 2972 31309 2975
rect 31260 2944 31309 2972
rect 31260 2932 31266 2944
rect 31297 2941 31309 2944
rect 31343 2941 31355 2975
rect 31297 2935 31355 2941
rect 32306 2932 32312 2984
rect 32364 2972 32370 2984
rect 32401 2975 32459 2981
rect 32401 2972 32413 2975
rect 32364 2944 32413 2972
rect 32364 2932 32370 2944
rect 32401 2941 32413 2944
rect 32447 2941 32459 2975
rect 32858 2972 32864 2984
rect 32819 2944 32864 2972
rect 32401 2935 32459 2941
rect 32858 2932 32864 2944
rect 32916 2932 32922 2984
rect 36998 2932 37004 2984
rect 37056 2972 37062 2984
rect 37496 2975 37554 2981
rect 37496 2972 37508 2975
rect 37056 2944 37508 2972
rect 37056 2932 37062 2944
rect 37496 2941 37508 2944
rect 37542 2972 37554 2975
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 37542 2944 37933 2972
rect 37542 2941 37554 2944
rect 37496 2935 37554 2941
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 21876 2876 22048 2904
rect 22741 2907 22799 2913
rect 21876 2864 21882 2876
rect 22741 2873 22753 2907
rect 22787 2904 22799 2907
rect 24394 2904 24400 2916
rect 22787 2876 24400 2904
rect 22787 2873 22799 2876
rect 22741 2867 22799 2873
rect 24394 2864 24400 2876
rect 24452 2864 24458 2916
rect 24489 2907 24547 2913
rect 24489 2873 24501 2907
rect 24535 2904 24547 2907
rect 25086 2907 25144 2913
rect 25086 2904 25098 2907
rect 24535 2876 25098 2904
rect 24535 2873 24547 2876
rect 24489 2867 24547 2873
rect 25086 2873 25098 2876
rect 25132 2873 25144 2907
rect 26697 2907 26755 2913
rect 25086 2867 25144 2873
rect 25700 2876 26556 2904
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12636 2808 12909 2836
rect 9309 2799 9367 2805
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 12897 2799 12955 2805
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 13817 2839 13875 2845
rect 13817 2836 13829 2839
rect 13780 2808 13829 2836
rect 13780 2796 13786 2808
rect 13817 2805 13829 2808
rect 13863 2805 13875 2839
rect 13817 2799 13875 2805
rect 14090 2796 14096 2848
rect 14148 2836 14154 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 14148 2808 14473 2836
rect 14148 2796 14154 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 14461 2799 14519 2805
rect 14642 2796 14648 2848
rect 14700 2836 14706 2848
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 14700 2808 15025 2836
rect 14700 2796 14706 2808
rect 15013 2805 15025 2808
rect 15059 2805 15071 2839
rect 15013 2799 15071 2805
rect 15562 2796 15568 2848
rect 15620 2836 15626 2848
rect 18322 2836 18328 2848
rect 15620 2808 18328 2836
rect 15620 2796 15626 2808
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 25700 2845 25728 2876
rect 19705 2839 19763 2845
rect 19705 2836 19717 2839
rect 19576 2808 19717 2836
rect 19576 2796 19582 2808
rect 19705 2805 19717 2808
rect 19751 2805 19763 2839
rect 19705 2799 19763 2805
rect 25685 2839 25743 2845
rect 25685 2805 25697 2839
rect 25731 2805 25743 2839
rect 26528 2836 26556 2876
rect 26697 2873 26709 2907
rect 26743 2904 26755 2907
rect 27525 2907 27583 2913
rect 27525 2904 27537 2907
rect 26743 2876 27537 2904
rect 26743 2873 26755 2876
rect 26697 2867 26755 2873
rect 27525 2873 27537 2876
rect 27571 2873 27583 2907
rect 27525 2867 27583 2873
rect 28307 2907 28365 2913
rect 28307 2873 28319 2907
rect 28353 2904 28365 2907
rect 29086 2904 29092 2916
rect 28353 2876 29092 2904
rect 28353 2873 28365 2876
rect 28307 2867 28365 2873
rect 26712 2836 26740 2867
rect 29086 2864 29092 2876
rect 29144 2864 29150 2916
rect 29365 2907 29423 2913
rect 29365 2873 29377 2907
rect 29411 2873 29423 2907
rect 29365 2867 29423 2873
rect 26528 2808 26740 2836
rect 28077 2839 28135 2845
rect 25685 2799 25743 2805
rect 28077 2805 28089 2839
rect 28123 2836 28135 2839
rect 28166 2836 28172 2848
rect 28123 2808 28172 2836
rect 28123 2805 28135 2808
rect 28077 2799 28135 2805
rect 28166 2796 28172 2808
rect 28224 2796 28230 2848
rect 28997 2839 29055 2845
rect 28997 2805 29009 2839
rect 29043 2836 29055 2839
rect 29380 2836 29408 2867
rect 29454 2864 29460 2916
rect 29512 2904 29518 2916
rect 32122 2904 32128 2916
rect 29512 2876 29557 2904
rect 30208 2876 32128 2904
rect 29512 2864 29518 2876
rect 30208 2836 30236 2876
rect 32122 2864 32128 2876
rect 32180 2864 32186 2916
rect 35069 2907 35127 2913
rect 35069 2873 35081 2907
rect 35115 2873 35127 2907
rect 35069 2867 35127 2873
rect 35713 2907 35771 2913
rect 35713 2873 35725 2907
rect 35759 2904 35771 2907
rect 37599 2907 37657 2913
rect 37599 2904 37611 2907
rect 35759 2876 37611 2904
rect 35759 2873 35771 2876
rect 35713 2867 35771 2873
rect 37599 2873 37611 2876
rect 37645 2873 37657 2907
rect 37599 2867 37657 2873
rect 29043 2808 30236 2836
rect 29043 2805 29055 2808
rect 28997 2799 29055 2805
rect 34698 2796 34704 2848
rect 34756 2836 34762 2848
rect 35084 2836 35112 2867
rect 34756 2808 35112 2836
rect 34756 2796 34762 2808
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 2038 2632 2044 2644
rect 1999 2604 2044 2632
rect 2038 2592 2044 2604
rect 2096 2632 2102 2644
rect 2096 2604 2360 2632
rect 2096 2592 2102 2604
rect 2222 2564 2228 2576
rect 2183 2536 2228 2564
rect 2222 2524 2228 2536
rect 2280 2524 2286 2576
rect 2332 2573 2360 2604
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 4764 2604 5365 2632
rect 4764 2592 4770 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 5353 2595 5411 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 9217 2635 9275 2641
rect 9217 2601 9229 2635
rect 9263 2632 9275 2635
rect 9306 2632 9312 2644
rect 9263 2604 9312 2632
rect 9263 2601 9275 2604
rect 9217 2595 9275 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 12802 2592 12808 2644
rect 12860 2592 12866 2644
rect 13262 2632 13268 2644
rect 13223 2604 13268 2632
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 14056 2604 14105 2632
rect 14056 2592 14062 2604
rect 14093 2601 14105 2604
rect 14139 2632 14151 2635
rect 14734 2632 14740 2644
rect 14139 2604 14740 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17310 2632 17316 2644
rect 16991 2604 17316 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2533 2375 2567
rect 2317 2527 2375 2533
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 4798 2564 4804 2576
rect 2915 2536 4804 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 7944 2564 7972 2592
rect 8846 2564 8852 2576
rect 7944 2536 8616 2564
rect 8807 2536 8852 2564
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 3384 2468 4721 2496
rect 3384 2456 3390 2468
rect 4709 2465 4721 2468
rect 4755 2496 4767 2499
rect 4893 2499 4951 2505
rect 4893 2496 4905 2499
rect 4755 2468 4905 2496
rect 4755 2465 4767 2468
rect 4709 2459 4767 2465
rect 4893 2465 4905 2468
rect 4939 2496 4951 2499
rect 5074 2496 5080 2508
rect 4939 2468 5080 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5442 2496 5448 2508
rect 5215 2468 5448 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6914 2496 6920 2508
rect 6779 2468 6920 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 7699 2468 8401 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8389 2465 8401 2468
rect 8435 2496 8447 2499
rect 8478 2496 8484 2508
rect 8435 2468 8484 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8588 2505 8616 2536
rect 8846 2524 8852 2536
rect 8904 2524 8910 2576
rect 9950 2564 9956 2576
rect 9911 2536 9956 2564
rect 9950 2524 9956 2536
rect 10008 2524 10014 2576
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 11241 2567 11299 2573
rect 11241 2564 11253 2567
rect 11112 2536 11253 2564
rect 11112 2524 11118 2536
rect 11241 2533 11253 2536
rect 11287 2564 11299 2567
rect 12621 2567 12679 2573
rect 12621 2564 12633 2567
rect 11287 2536 12633 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 12621 2533 12633 2536
rect 12667 2564 12679 2567
rect 12820 2564 12848 2592
rect 12667 2536 16988 2564
rect 12667 2533 12679 2536
rect 12621 2527 12679 2533
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2465 8631 2499
rect 8573 2459 8631 2465
rect 11368 2499 11426 2505
rect 11368 2465 11380 2499
rect 11414 2465 11426 2499
rect 12526 2496 12532 2508
rect 11368 2459 11426 2465
rect 11992 2468 12532 2496
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 3145 2431 3203 2437
rect 3145 2428 3157 2431
rect 2280 2400 3157 2428
rect 2280 2388 2286 2400
rect 3145 2397 3157 2400
rect 3191 2397 3203 2431
rect 6270 2428 6276 2440
rect 3145 2391 3203 2397
rect 4126 2400 6276 2428
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 1673 2363 1731 2369
rect 1673 2360 1685 2363
rect 1636 2332 1685 2360
rect 1636 2320 1642 2332
rect 1673 2329 1685 2332
rect 1719 2360 1731 2363
rect 4126 2360 4154 2400
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9364 2400 9873 2428
rect 9364 2388 9370 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 9861 2391 9919 2397
rect 10134 2388 10140 2400
rect 10192 2428 10198 2440
rect 11383 2428 11411 2459
rect 10192 2400 11411 2428
rect 10192 2388 10198 2400
rect 4982 2360 4988 2372
rect 1719 2332 4154 2360
rect 4943 2332 4988 2360
rect 1719 2329 1731 2332
rect 1673 2323 1731 2329
rect 4982 2320 4988 2332
rect 5040 2360 5046 2372
rect 5905 2363 5963 2369
rect 5905 2360 5917 2363
rect 5040 2332 5917 2360
rect 5040 2320 5046 2332
rect 5905 2329 5917 2332
rect 5951 2329 5963 2363
rect 5905 2323 5963 2329
rect 7101 2363 7159 2369
rect 7101 2329 7113 2363
rect 7147 2360 7159 2363
rect 9398 2360 9404 2372
rect 7147 2332 9404 2360
rect 7147 2329 7159 2332
rect 7101 2323 7159 2329
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2292 4491 2295
rect 5442 2292 5448 2304
rect 4479 2264 5448 2292
rect 4479 2261 4491 2264
rect 4433 2255 4491 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5920 2292 5948 2323
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 11992 2360 12020 2468
rect 12526 2456 12532 2468
rect 12584 2496 12590 2508
rect 13722 2496 13728 2508
rect 12584 2468 13728 2496
rect 12584 2456 12590 2468
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13964 2468 14197 2496
rect 13964 2456 13970 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15252 2468 15577 2496
rect 15252 2456 15258 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 16574 2496 16580 2508
rect 16535 2468 16580 2496
rect 15565 2459 15623 2465
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12115 2400 13001 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12989 2397 13001 2400
rect 13035 2428 13047 2431
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 13035 2400 13829 2428
rect 13035 2397 13047 2400
rect 12989 2391 13047 2397
rect 13817 2397 13829 2400
rect 13863 2397 13875 2431
rect 16960 2428 16988 2536
rect 17052 2505 17080 2604
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17586 2632 17592 2644
rect 17547 2604 17592 2632
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 18064 2604 20085 2632
rect 18064 2564 18092 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 21358 2632 21364 2644
rect 21319 2604 21364 2632
rect 20073 2595 20131 2601
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 24762 2632 24768 2644
rect 23835 2604 24768 2632
rect 18322 2564 18328 2576
rect 17144 2536 18092 2564
rect 18283 2536 18328 2564
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 17144 2428 17172 2536
rect 18322 2524 18328 2536
rect 18380 2524 18386 2576
rect 19705 2567 19763 2573
rect 19705 2533 19717 2567
rect 19751 2564 19763 2567
rect 19794 2564 19800 2576
rect 19751 2536 19800 2564
rect 19751 2533 19763 2536
rect 19705 2527 19763 2533
rect 19794 2524 19800 2536
rect 19852 2524 19858 2576
rect 21729 2567 21787 2573
rect 21729 2533 21741 2567
rect 21775 2564 21787 2567
rect 22097 2567 22155 2573
rect 22097 2564 22109 2567
rect 21775 2536 22109 2564
rect 21775 2533 21787 2536
rect 21729 2527 21787 2533
rect 22097 2533 22109 2536
rect 22143 2564 22155 2567
rect 23109 2567 23167 2573
rect 22143 2536 22968 2564
rect 22143 2533 22155 2536
rect 22097 2527 22155 2533
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18049 2499 18107 2505
rect 18049 2496 18061 2499
rect 18012 2468 18061 2496
rect 18012 2456 18018 2468
rect 18049 2465 18061 2468
rect 18095 2496 18107 2499
rect 18417 2499 18475 2505
rect 18417 2496 18429 2499
rect 18095 2468 18429 2496
rect 18095 2465 18107 2468
rect 18049 2459 18107 2465
rect 18417 2465 18429 2468
rect 18463 2465 18475 2499
rect 18417 2459 18475 2465
rect 19150 2456 19156 2508
rect 19208 2496 19214 2508
rect 22940 2505 22968 2536
rect 23109 2533 23121 2567
rect 23155 2564 23167 2567
rect 23835 2564 23863 2604
rect 24762 2592 24768 2604
rect 24820 2632 24826 2644
rect 25041 2635 25099 2641
rect 25041 2632 25053 2635
rect 24820 2604 25053 2632
rect 24820 2592 24826 2604
rect 25041 2601 25053 2604
rect 25087 2601 25099 2635
rect 25406 2632 25412 2644
rect 25367 2604 25412 2632
rect 25041 2595 25099 2601
rect 25406 2592 25412 2604
rect 25464 2592 25470 2644
rect 26326 2632 26332 2644
rect 26287 2604 26332 2632
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 28813 2635 28871 2641
rect 28813 2601 28825 2635
rect 28859 2632 28871 2635
rect 29454 2632 29460 2644
rect 28859 2604 29460 2632
rect 28859 2601 28871 2604
rect 28813 2595 28871 2601
rect 29454 2592 29460 2604
rect 29512 2592 29518 2644
rect 29546 2592 29552 2644
rect 29604 2632 29610 2644
rect 29604 2604 29649 2632
rect 29604 2592 29610 2604
rect 30006 2592 30012 2644
rect 30064 2632 30070 2644
rect 30064 2604 31375 2632
rect 30064 2592 30070 2604
rect 24854 2564 24860 2576
rect 23155 2536 23863 2564
rect 24228 2536 24860 2564
rect 23155 2533 23167 2536
rect 23109 2527 23167 2533
rect 24228 2505 24256 2536
rect 24854 2524 24860 2536
rect 24912 2524 24918 2576
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19208 2468 19901 2496
rect 19208 2456 19214 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 19889 2459 19947 2465
rect 20916 2468 21189 2496
rect 16960 2400 17172 2428
rect 13817 2391 13875 2397
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 20916 2437 20944 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 22373 2499 22431 2505
rect 22373 2496 22385 2499
rect 21177 2459 21235 2465
rect 21744 2468 22385 2496
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 18196 2400 20913 2428
rect 18196 2388 18202 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21744 2372 21772 2468
rect 22373 2465 22385 2468
rect 22419 2465 22431 2499
rect 22373 2459 22431 2465
rect 22925 2499 22983 2505
rect 22925 2465 22937 2499
rect 22971 2496 22983 2499
rect 23845 2499 23903 2505
rect 22971 2468 23428 2496
rect 22971 2465 22983 2468
rect 22925 2459 22983 2465
rect 9646 2332 12020 2360
rect 12437 2363 12495 2369
rect 8202 2292 8208 2304
rect 5920 2264 8208 2292
rect 8202 2252 8208 2264
rect 8260 2292 8266 2304
rect 9646 2292 9674 2332
rect 12437 2329 12449 2363
rect 12483 2360 12495 2363
rect 16114 2360 16120 2372
rect 12483 2332 16120 2360
rect 12483 2329 12495 2332
rect 12437 2323 12495 2329
rect 12912 2304 12940 2332
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 17221 2363 17279 2369
rect 17221 2329 17233 2363
rect 17267 2360 17279 2363
rect 17770 2360 17776 2372
rect 17267 2332 17776 2360
rect 17267 2329 17279 2332
rect 17221 2323 17279 2329
rect 17770 2320 17776 2332
rect 17828 2320 17834 2372
rect 18966 2320 18972 2372
rect 19024 2360 19030 2372
rect 20533 2363 20591 2369
rect 20533 2360 20545 2363
rect 19024 2332 20545 2360
rect 19024 2320 19030 2332
rect 20533 2329 20545 2332
rect 20579 2360 20591 2363
rect 21726 2360 21732 2372
rect 20579 2332 21732 2360
rect 20579 2329 20591 2332
rect 20533 2323 20591 2329
rect 21726 2320 21732 2332
rect 21784 2320 21790 2372
rect 22388 2360 22416 2459
rect 23400 2440 23428 2468
rect 23845 2465 23857 2499
rect 23891 2496 23903 2499
rect 24213 2499 24271 2505
rect 24213 2496 24225 2499
rect 23891 2468 24225 2496
rect 23891 2465 23903 2468
rect 23845 2459 23903 2465
rect 24213 2465 24225 2468
rect 24259 2465 24271 2499
rect 24489 2499 24547 2505
rect 24489 2496 24501 2499
rect 24213 2459 24271 2465
rect 24320 2468 24501 2496
rect 23382 2428 23388 2440
rect 23295 2400 23388 2428
rect 23382 2388 23388 2400
rect 23440 2428 23446 2440
rect 24320 2428 24348 2468
rect 24489 2465 24501 2468
rect 24535 2465 24547 2499
rect 25424 2496 25452 2592
rect 27341 2567 27399 2573
rect 27341 2533 27353 2567
rect 27387 2564 27399 2567
rect 28166 2564 28172 2576
rect 27387 2536 28028 2564
rect 28127 2536 28172 2564
rect 27387 2533 27399 2536
rect 27341 2527 27399 2533
rect 25628 2499 25686 2505
rect 25628 2496 25640 2499
rect 25424 2468 25640 2496
rect 24489 2459 24547 2465
rect 25628 2465 25640 2468
rect 25674 2465 25686 2499
rect 27430 2496 27436 2508
rect 25628 2459 25686 2465
rect 26620 2468 27436 2496
rect 23440 2400 24348 2428
rect 24765 2431 24823 2437
rect 23440 2388 23446 2400
rect 24765 2397 24777 2431
rect 24811 2428 24823 2431
rect 26142 2428 26148 2440
rect 24811 2400 26148 2428
rect 24811 2397 24823 2400
rect 24765 2391 24823 2397
rect 26142 2388 26148 2400
rect 26200 2388 26206 2440
rect 26620 2369 26648 2468
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 28000 2505 28028 2536
rect 28166 2524 28172 2536
rect 28224 2524 28230 2576
rect 28994 2524 29000 2576
rect 29052 2564 29058 2576
rect 29089 2567 29147 2573
rect 29089 2564 29101 2567
rect 29052 2536 29101 2564
rect 29052 2524 29058 2536
rect 29089 2533 29101 2536
rect 29135 2533 29147 2567
rect 29089 2527 29147 2533
rect 27985 2499 28043 2505
rect 27985 2465 27997 2499
rect 28031 2496 28043 2499
rect 28626 2496 28632 2508
rect 28031 2468 28632 2496
rect 28031 2465 28043 2468
rect 27985 2459 28043 2465
rect 28626 2456 28632 2468
rect 28684 2456 28690 2508
rect 29564 2496 29592 2592
rect 30466 2564 30472 2576
rect 30427 2536 30472 2564
rect 30466 2524 30472 2536
rect 30524 2524 30530 2576
rect 30929 2567 30987 2573
rect 30929 2533 30941 2567
rect 30975 2564 30987 2567
rect 31202 2564 31208 2576
rect 30975 2536 31208 2564
rect 30975 2533 30987 2536
rect 30929 2527 30987 2533
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29564 2468 29745 2496
rect 29733 2465 29745 2468
rect 29779 2465 29791 2499
rect 29733 2459 29791 2465
rect 30285 2499 30343 2505
rect 30285 2465 30297 2499
rect 30331 2496 30343 2499
rect 30944 2496 30972 2527
rect 31202 2524 31208 2536
rect 31260 2524 31266 2576
rect 31347 2564 31375 2604
rect 31478 2592 31484 2644
rect 31536 2632 31542 2644
rect 32585 2635 32643 2641
rect 32585 2632 32597 2635
rect 31536 2604 32597 2632
rect 31536 2592 31542 2604
rect 32585 2601 32597 2604
rect 32631 2601 32643 2635
rect 34054 2632 34060 2644
rect 34015 2604 34060 2632
rect 32585 2595 32643 2601
rect 34054 2592 34060 2604
rect 34112 2592 34118 2644
rect 34974 2632 34980 2644
rect 34935 2604 34980 2632
rect 34974 2592 34980 2604
rect 35032 2592 35038 2644
rect 35618 2592 35624 2644
rect 35676 2632 35682 2644
rect 35897 2635 35955 2641
rect 35897 2632 35909 2635
rect 35676 2604 35909 2632
rect 35676 2592 35682 2604
rect 35897 2601 35909 2604
rect 35943 2601 35955 2635
rect 35897 2595 35955 2601
rect 31757 2567 31815 2573
rect 31757 2564 31769 2567
rect 31347 2536 31769 2564
rect 31347 2505 31375 2536
rect 31757 2533 31769 2536
rect 31803 2533 31815 2567
rect 31757 2527 31815 2533
rect 30331 2468 30972 2496
rect 31332 2499 31390 2505
rect 30331 2465 30343 2468
rect 30285 2459 30343 2465
rect 31332 2465 31344 2499
rect 31378 2465 31390 2499
rect 31332 2459 31390 2465
rect 33648 2499 33706 2505
rect 33648 2465 33660 2499
rect 33694 2496 33706 2499
rect 34072 2496 34100 2592
rect 33694 2468 34100 2496
rect 35504 2499 35562 2505
rect 33694 2465 33706 2468
rect 33648 2459 33706 2465
rect 35504 2465 35516 2499
rect 35550 2496 35562 2499
rect 35636 2496 35664 2592
rect 35550 2468 35664 2496
rect 36516 2499 36574 2505
rect 35550 2465 35562 2468
rect 35504 2459 35562 2465
rect 36516 2465 36528 2499
rect 36562 2496 36574 2499
rect 36906 2496 36912 2508
rect 36562 2468 36912 2496
rect 36562 2465 36574 2468
rect 36516 2459 36574 2465
rect 36906 2456 36912 2468
rect 36964 2456 36970 2508
rect 31435 2431 31493 2437
rect 31435 2397 31447 2431
rect 31481 2428 31493 2431
rect 31754 2428 31760 2440
rect 31481 2400 31760 2428
rect 31481 2397 31493 2400
rect 31435 2391 31493 2397
rect 31754 2388 31760 2400
rect 31812 2388 31818 2440
rect 31941 2431 31999 2437
rect 31941 2397 31953 2431
rect 31987 2428 31999 2431
rect 33735 2431 33793 2437
rect 33735 2428 33747 2431
rect 31987 2400 33747 2428
rect 31987 2397 31999 2400
rect 31941 2391 31999 2397
rect 33735 2397 33747 2400
rect 33781 2397 33793 2431
rect 33735 2391 33793 2397
rect 26605 2363 26663 2369
rect 26605 2360 26617 2363
rect 22388 2332 26617 2360
rect 26605 2329 26617 2332
rect 26651 2329 26663 2363
rect 26605 2323 26663 2329
rect 31202 2320 31208 2372
rect 31260 2360 31266 2372
rect 32125 2363 32183 2369
rect 32125 2360 32137 2363
rect 31260 2332 32137 2360
rect 31260 2320 31266 2332
rect 32125 2329 32137 2332
rect 32171 2360 32183 2363
rect 32858 2360 32864 2372
rect 32171 2332 32864 2360
rect 32171 2329 32183 2332
rect 32125 2323 32183 2329
rect 32858 2320 32864 2332
rect 32916 2360 32922 2372
rect 33045 2363 33103 2369
rect 33045 2360 33057 2363
rect 32916 2332 33057 2360
rect 32916 2320 32922 2332
rect 33045 2329 33057 2332
rect 33091 2329 33103 2363
rect 33045 2323 33103 2329
rect 35575 2363 35633 2369
rect 35575 2329 35587 2363
rect 35621 2360 35633 2363
rect 36078 2360 36084 2372
rect 35621 2332 36084 2360
rect 35621 2329 35633 2332
rect 35575 2323 35633 2329
rect 36078 2320 36084 2332
rect 36136 2320 36142 2372
rect 8260 2264 9674 2292
rect 11471 2295 11529 2301
rect 8260 2252 8266 2264
rect 11471 2261 11483 2295
rect 11517 2292 11529 2295
rect 12250 2292 12256 2304
rect 11517 2264 12256 2292
rect 11517 2261 11529 2264
rect 11471 2255 11529 2261
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 12618 2252 12624 2304
rect 12676 2292 12682 2304
rect 12759 2295 12817 2301
rect 12759 2292 12771 2295
rect 12676 2264 12771 2292
rect 12676 2252 12682 2264
rect 12759 2261 12771 2264
rect 12805 2261 12817 2295
rect 12894 2292 12900 2304
rect 12855 2264 12900 2292
rect 12759 2255 12817 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 12986 2252 12992 2304
rect 13044 2292 13050 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13044 2264 13645 2292
rect 13044 2252 13050 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 13817 2295 13875 2301
rect 13817 2261 13829 2295
rect 13863 2292 13875 2295
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 13863 2264 14381 2292
rect 13863 2261 13875 2264
rect 13817 2255 13875 2261
rect 14369 2261 14381 2264
rect 14415 2292 14427 2295
rect 14642 2292 14648 2304
rect 14415 2264 14648 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 14826 2292 14832 2304
rect 14787 2264 14832 2292
rect 14826 2252 14832 2264
rect 14884 2292 14890 2304
rect 15654 2292 15660 2304
rect 14884 2264 15660 2292
rect 14884 2252 14890 2264
rect 15654 2252 15660 2264
rect 15712 2292 15718 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15712 2264 15761 2292
rect 15712 2252 15718 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 25731 2295 25789 2301
rect 25731 2261 25743 2295
rect 25777 2292 25789 2295
rect 26510 2292 26516 2304
rect 25777 2264 26516 2292
rect 25777 2261 25789 2264
rect 25731 2255 25789 2261
rect 26510 2252 26516 2264
rect 26568 2252 26574 2304
rect 27522 2252 27528 2304
rect 27580 2292 27586 2304
rect 31941 2295 31999 2301
rect 31941 2292 31953 2295
rect 27580 2264 31953 2292
rect 27580 2252 27586 2264
rect 31941 2261 31953 2264
rect 31987 2261 31999 2295
rect 31941 2255 31999 2261
rect 35986 2252 35992 2304
rect 36044 2292 36050 2304
rect 36587 2295 36645 2301
rect 36587 2292 36599 2295
rect 36044 2264 36599 2292
rect 36044 2252 36050 2264
rect 36587 2261 36599 2264
rect 36633 2261 36645 2295
rect 36587 2255 36645 2261
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 112 12928 164 12980
rect 39580 12928 39632 12980
rect 5356 12656 5408 12708
rect 16764 12724 16816 12776
rect 32220 12724 32272 12776
rect 1584 12588 1636 12640
rect 3792 12588 3844 12640
rect 5172 12588 5224 12640
rect 5448 12631 5500 12640
rect 5448 12597 5457 12631
rect 5457 12597 5491 12631
rect 5491 12597 5500 12631
rect 5448 12588 5500 12597
rect 11888 12588 11940 12640
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 1032 12384 1084 12436
rect 5356 12316 5408 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 112 12112 164 12164
rect 6184 12248 6236 12300
rect 10508 12248 10560 12300
rect 12256 12248 12308 12300
rect 13452 12248 13504 12300
rect 4620 12112 4672 12164
rect 2136 12044 2188 12096
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 4344 12044 4396 12096
rect 7472 12044 7524 12096
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 11796 12044 11848 12096
rect 14096 12044 14148 12096
rect 14280 12087 14332 12096
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 2504 11840 2556 11892
rect 5448 11840 5500 11892
rect 5540 11840 5592 11892
rect 14096 11883 14148 11892
rect 20 11772 72 11824
rect 3700 11772 3752 11824
rect 1400 11704 1452 11756
rect 7104 11704 7156 11756
rect 14096 11849 14105 11883
rect 14105 11849 14139 11883
rect 14139 11849 14148 11883
rect 14096 11840 14148 11849
rect 15476 11772 15528 11824
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 2320 11679 2372 11688
rect 2320 11645 2329 11679
rect 2329 11645 2363 11679
rect 2363 11645 2372 11679
rect 2320 11636 2372 11645
rect 4712 11636 4764 11688
rect 4896 11636 4948 11688
rect 5540 11636 5592 11688
rect 4068 11568 4120 11620
rect 5448 11568 5500 11620
rect 10600 11636 10652 11688
rect 2044 11500 2096 11552
rect 4620 11500 4672 11552
rect 6184 11500 6236 11552
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 10508 11500 10560 11552
rect 11520 11500 11572 11552
rect 13360 11636 13412 11688
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 12256 11568 12308 11620
rect 14096 11568 14148 11620
rect 17316 11636 17368 11688
rect 19248 11636 19300 11688
rect 15016 11611 15068 11620
rect 15016 11577 15025 11611
rect 15025 11577 15059 11611
rect 15059 11577 15068 11611
rect 15016 11568 15068 11577
rect 15752 11568 15804 11620
rect 22008 11568 22060 11620
rect 12072 11500 12124 11552
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12440 11500 12492 11509
rect 13452 11500 13504 11552
rect 18788 11500 18840 11552
rect 19248 11500 19300 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 19524 11296 19576 11348
rect 35624 11339 35676 11348
rect 35624 11305 35633 11339
rect 35633 11305 35667 11339
rect 35667 11305 35676 11339
rect 35624 11296 35676 11305
rect 4712 11228 4764 11280
rect 1768 11160 1820 11212
rect 2320 11203 2372 11212
rect 2320 11169 2329 11203
rect 2329 11169 2363 11203
rect 2363 11169 2372 11203
rect 2320 11160 2372 11169
rect 3884 11160 3936 11212
rect 5264 11160 5316 11212
rect 6092 11203 6144 11212
rect 6092 11169 6101 11203
rect 6101 11169 6135 11203
rect 6135 11169 6144 11203
rect 6092 11160 6144 11169
rect 7104 11203 7156 11212
rect 7104 11169 7113 11203
rect 7113 11169 7147 11203
rect 7147 11169 7156 11203
rect 7104 11160 7156 11169
rect 8576 11160 8628 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 11244 11160 11296 11212
rect 11704 11160 11756 11212
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 16672 11160 16724 11212
rect 18512 11160 18564 11212
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 22652 11160 22704 11212
rect 26976 11160 27028 11212
rect 34152 11160 34204 11212
rect 34612 11160 34664 11212
rect 35440 11203 35492 11212
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 2228 11092 2280 11144
rect 12808 11092 12860 11144
rect 15200 11092 15252 11144
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 3608 11024 3660 11076
rect 6460 11024 6512 11076
rect 12164 11024 12216 11076
rect 1768 10999 1820 11008
rect 1768 10965 1777 10999
rect 1777 10965 1811 10999
rect 1811 10965 1820 10999
rect 1768 10956 1820 10965
rect 3516 10956 3568 11008
rect 4804 10956 4856 11008
rect 6368 10956 6420 11008
rect 13084 10956 13136 11008
rect 18972 10956 19024 11008
rect 19800 10956 19852 11008
rect 24492 10956 24544 11008
rect 29092 10956 29144 11008
rect 36176 10956 36228 11008
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 940 10752 992 10804
rect 4528 10795 4580 10804
rect 4528 10761 4537 10795
rect 4537 10761 4571 10795
rect 4571 10761 4580 10795
rect 4528 10752 4580 10761
rect 5264 10752 5316 10804
rect 6276 10752 6328 10804
rect 10416 10752 10468 10804
rect 18512 10795 18564 10804
rect 11612 10684 11664 10736
rect 14096 10684 14148 10736
rect 2136 10616 2188 10668
rect 7104 10616 7156 10668
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 11244 10616 11296 10668
rect 2504 10548 2556 10600
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 5264 10548 5316 10600
rect 5632 10591 5684 10600
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 3976 10480 4028 10532
rect 9496 10548 9548 10600
rect 12900 10616 12952 10668
rect 12256 10548 12308 10600
rect 12348 10480 12400 10532
rect 2780 10412 2832 10464
rect 3884 10412 3936 10464
rect 4528 10412 4580 10464
rect 6092 10412 6144 10464
rect 7288 10412 7340 10464
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 9680 10412 9732 10464
rect 10232 10412 10284 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12072 10412 12124 10464
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 18512 10761 18521 10795
rect 18521 10761 18555 10795
rect 18555 10761 18564 10795
rect 18512 10752 18564 10761
rect 22652 10795 22704 10804
rect 22652 10761 22661 10795
rect 22661 10761 22695 10795
rect 22695 10761 22704 10795
rect 22652 10752 22704 10761
rect 26240 10795 26292 10804
rect 26240 10761 26249 10795
rect 26249 10761 26283 10795
rect 26283 10761 26292 10795
rect 26240 10752 26292 10761
rect 35440 10752 35492 10804
rect 35624 10727 35676 10736
rect 35624 10693 35633 10727
rect 35633 10693 35667 10727
rect 35667 10693 35676 10727
rect 35624 10684 35676 10693
rect 17684 10616 17736 10668
rect 19248 10616 19300 10668
rect 14832 10523 14884 10532
rect 14832 10489 14841 10523
rect 14841 10489 14875 10523
rect 14875 10489 14884 10523
rect 14832 10480 14884 10489
rect 16488 10548 16540 10600
rect 17960 10591 18012 10600
rect 17960 10557 17969 10591
rect 17969 10557 18003 10591
rect 18003 10557 18012 10591
rect 17960 10548 18012 10557
rect 18328 10548 18380 10600
rect 20260 10548 20312 10600
rect 28080 10616 28132 10668
rect 35348 10616 35400 10668
rect 16580 10523 16632 10532
rect 16580 10489 16589 10523
rect 16589 10489 16623 10523
rect 16623 10489 16632 10523
rect 16580 10480 16632 10489
rect 18604 10480 18656 10532
rect 25044 10548 25096 10600
rect 26240 10548 26292 10600
rect 26608 10548 26660 10600
rect 27988 10548 28040 10600
rect 23020 10480 23072 10532
rect 28632 10480 28684 10532
rect 12716 10455 12768 10464
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 16672 10412 16724 10464
rect 17132 10412 17184 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 20076 10412 20128 10464
rect 22100 10412 22152 10464
rect 25964 10412 26016 10464
rect 26976 10412 27028 10464
rect 27252 10412 27304 10464
rect 33048 10412 33100 10464
rect 33692 10455 33744 10464
rect 33692 10421 33701 10455
rect 33701 10421 33735 10455
rect 33735 10421 33744 10455
rect 33692 10412 33744 10421
rect 34612 10412 34664 10464
rect 35164 10412 35216 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 3516 10251 3568 10260
rect 3516 10217 3525 10251
rect 3525 10217 3559 10251
rect 3559 10217 3568 10251
rect 3516 10208 3568 10217
rect 6736 10251 6788 10260
rect 3148 10140 3200 10192
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 6920 10208 6972 10260
rect 13268 10208 13320 10260
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 27252 10208 27304 10260
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 1768 10072 1820 10124
rect 2412 10072 2464 10124
rect 2688 10072 2740 10124
rect 4436 10140 4488 10192
rect 6828 10140 6880 10192
rect 10600 10140 10652 10192
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 2320 10004 2372 10056
rect 3884 10004 3936 10056
rect 6000 10072 6052 10124
rect 6920 10115 6972 10124
rect 6920 10081 6929 10115
rect 6929 10081 6963 10115
rect 6963 10081 6972 10115
rect 6920 10072 6972 10081
rect 6552 10004 6604 10056
rect 9404 10072 9456 10124
rect 10232 10072 10284 10124
rect 11612 10072 11664 10124
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 12624 9936 12676 9988
rect 2504 9868 2556 9920
rect 3240 9868 3292 9920
rect 4620 9868 4672 9920
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 12992 10140 13044 10192
rect 27436 10183 27488 10192
rect 27436 10149 27445 10183
rect 27445 10149 27479 10183
rect 27479 10149 27488 10183
rect 27436 10140 27488 10149
rect 13268 10072 13320 10124
rect 12808 9936 12860 9988
rect 15476 9936 15528 9988
rect 16488 10072 16540 10124
rect 17776 10115 17828 10124
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 17868 10072 17920 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 20812 10072 20864 10124
rect 22376 10072 22428 10124
rect 22928 10115 22980 10124
rect 22928 10081 22937 10115
rect 22937 10081 22971 10115
rect 22971 10081 22980 10115
rect 22928 10072 22980 10081
rect 24400 10115 24452 10124
rect 24400 10081 24409 10115
rect 24409 10081 24443 10115
rect 24443 10081 24452 10115
rect 24400 10072 24452 10081
rect 25504 10072 25556 10124
rect 28724 10072 28776 10124
rect 33508 10115 33560 10124
rect 33508 10081 33526 10115
rect 33526 10081 33560 10115
rect 35440 10208 35492 10260
rect 35716 10208 35768 10260
rect 33508 10072 33560 10081
rect 34704 10072 34756 10124
rect 35900 10072 35952 10124
rect 36084 10072 36136 10124
rect 18512 10047 18564 10056
rect 16304 10004 16356 10013
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 21548 10004 21600 10056
rect 27160 10004 27212 10056
rect 29184 10004 29236 10056
rect 18236 9936 18288 9988
rect 27068 9936 27120 9988
rect 35348 9936 35400 9988
rect 37464 10004 37516 10056
rect 36544 9936 36596 9988
rect 13176 9868 13228 9920
rect 14188 9868 14240 9920
rect 15292 9868 15344 9920
rect 19708 9868 19760 9920
rect 20168 9868 20220 9920
rect 21272 9868 21324 9920
rect 21456 9868 21508 9920
rect 21824 9868 21876 9920
rect 23388 9868 23440 9920
rect 24768 9868 24820 9920
rect 28172 9868 28224 9920
rect 35440 9868 35492 9920
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 3884 9664 3936 9716
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 8208 9707 8260 9716
rect 6552 9664 6604 9673
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 3976 9596 4028 9648
rect 6000 9596 6052 9648
rect 6920 9596 6972 9648
rect 3516 9528 3568 9580
rect 3700 9528 3752 9580
rect 3884 9528 3936 9580
rect 5632 9528 5684 9580
rect 7564 9528 7616 9580
rect 8668 9528 8720 9580
rect 1676 9460 1728 9512
rect 2412 9460 2464 9512
rect 2504 9503 2556 9512
rect 2504 9469 2513 9503
rect 2513 9469 2547 9503
rect 2547 9469 2556 9503
rect 2504 9460 2556 9469
rect 2136 9435 2188 9444
rect 2136 9401 2145 9435
rect 2145 9401 2179 9435
rect 2179 9401 2188 9435
rect 2136 9392 2188 9401
rect 2688 9324 2740 9376
rect 3792 9460 3844 9512
rect 4160 9460 4212 9512
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5908 9460 5960 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 10692 9460 10744 9512
rect 11612 9664 11664 9716
rect 11796 9707 11848 9716
rect 11796 9673 11805 9707
rect 11805 9673 11839 9707
rect 11839 9673 11848 9707
rect 15476 9707 15528 9716
rect 11796 9664 11848 9673
rect 15476 9673 15485 9707
rect 15485 9673 15519 9707
rect 15519 9673 15528 9707
rect 15476 9664 15528 9673
rect 16488 9664 16540 9716
rect 17500 9707 17552 9716
rect 17500 9673 17509 9707
rect 17509 9673 17543 9707
rect 17543 9673 17552 9707
rect 17500 9664 17552 9673
rect 17776 9664 17828 9716
rect 19340 9707 19392 9716
rect 19340 9673 19349 9707
rect 19349 9673 19383 9707
rect 19383 9673 19392 9707
rect 19340 9664 19392 9673
rect 20812 9664 20864 9716
rect 21640 9664 21692 9716
rect 22376 9707 22428 9716
rect 22376 9673 22385 9707
rect 22385 9673 22419 9707
rect 22419 9673 22428 9707
rect 22376 9664 22428 9673
rect 26608 9664 26660 9716
rect 32220 9707 32272 9716
rect 13176 9596 13228 9648
rect 25504 9639 25556 9648
rect 12716 9528 12768 9580
rect 13728 9528 13780 9580
rect 15660 9528 15712 9580
rect 13544 9460 13596 9512
rect 3424 9392 3476 9444
rect 3700 9435 3752 9444
rect 3700 9401 3709 9435
rect 3709 9401 3743 9435
rect 3743 9401 3752 9435
rect 3700 9392 3752 9401
rect 3976 9324 4028 9376
rect 6000 9324 6052 9376
rect 7012 9435 7064 9444
rect 7012 9401 7021 9435
rect 7021 9401 7055 9435
rect 7055 9401 7064 9435
rect 7012 9392 7064 9401
rect 12532 9392 12584 9444
rect 13268 9392 13320 9444
rect 13820 9435 13872 9444
rect 13820 9401 13829 9435
rect 13829 9401 13863 9435
rect 13863 9401 13872 9435
rect 13820 9392 13872 9401
rect 18236 9460 18288 9512
rect 20536 9528 20588 9580
rect 25504 9605 25513 9639
rect 25513 9605 25547 9639
rect 25547 9605 25556 9639
rect 25504 9596 25556 9605
rect 27344 9596 27396 9648
rect 18880 9460 18932 9512
rect 19984 9460 20036 9512
rect 20168 9503 20220 9512
rect 20168 9469 20177 9503
rect 20177 9469 20211 9503
rect 20211 9469 20220 9503
rect 20168 9460 20220 9469
rect 24124 9503 24176 9512
rect 24124 9469 24133 9503
rect 24133 9469 24167 9503
rect 24167 9469 24176 9503
rect 24124 9460 24176 9469
rect 27252 9528 27304 9580
rect 8300 9324 8352 9376
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 12716 9324 12768 9376
rect 12992 9324 13044 9376
rect 16120 9435 16172 9444
rect 16120 9401 16129 9435
rect 16129 9401 16163 9435
rect 16163 9401 16172 9435
rect 16672 9435 16724 9444
rect 16120 9392 16172 9401
rect 16672 9401 16681 9435
rect 16681 9401 16715 9435
rect 16715 9401 16724 9435
rect 16672 9392 16724 9401
rect 21456 9435 21508 9444
rect 21456 9401 21465 9435
rect 21465 9401 21499 9435
rect 21499 9401 21508 9435
rect 21456 9392 21508 9401
rect 21548 9435 21600 9444
rect 21548 9401 21557 9435
rect 21557 9401 21591 9435
rect 21591 9401 21600 9435
rect 21548 9392 21600 9401
rect 23664 9392 23716 9444
rect 24860 9435 24912 9444
rect 24860 9401 24869 9435
rect 24869 9401 24903 9435
rect 24903 9401 24912 9435
rect 24860 9392 24912 9401
rect 29828 9503 29880 9512
rect 29828 9469 29837 9503
rect 29837 9469 29871 9503
rect 29871 9469 29880 9503
rect 29828 9460 29880 9469
rect 30288 9503 30340 9512
rect 30288 9469 30297 9503
rect 30297 9469 30331 9503
rect 30331 9469 30340 9503
rect 32220 9673 32229 9707
rect 32229 9673 32263 9707
rect 32263 9673 32272 9707
rect 32220 9664 32272 9673
rect 33508 9707 33560 9716
rect 33508 9673 33517 9707
rect 33517 9673 33551 9707
rect 33551 9673 33560 9707
rect 33508 9664 33560 9673
rect 35532 9707 35584 9716
rect 35532 9673 35541 9707
rect 35541 9673 35575 9707
rect 35575 9673 35584 9707
rect 35532 9664 35584 9673
rect 35900 9707 35952 9716
rect 35900 9673 35909 9707
rect 35909 9673 35943 9707
rect 35943 9673 35952 9707
rect 35900 9664 35952 9673
rect 37648 9664 37700 9716
rect 33600 9528 33652 9580
rect 35532 9528 35584 9580
rect 30288 9460 30340 9469
rect 27436 9392 27488 9444
rect 28080 9435 28132 9444
rect 15936 9324 15988 9376
rect 17868 9367 17920 9376
rect 17868 9333 17877 9367
rect 17877 9333 17911 9367
rect 17911 9333 17920 9367
rect 17868 9324 17920 9333
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 22468 9324 22520 9376
rect 22928 9367 22980 9376
rect 22928 9333 22937 9367
rect 22937 9333 22971 9367
rect 22971 9333 22980 9367
rect 22928 9324 22980 9333
rect 23388 9324 23440 9376
rect 26700 9324 26752 9376
rect 26884 9367 26936 9376
rect 26884 9333 26893 9367
rect 26893 9333 26927 9367
rect 26927 9333 26936 9367
rect 26884 9324 26936 9333
rect 28080 9401 28089 9435
rect 28089 9401 28123 9435
rect 28123 9401 28132 9435
rect 28080 9392 28132 9401
rect 32404 9392 32456 9444
rect 36452 9503 36504 9512
rect 36452 9469 36461 9503
rect 36461 9469 36495 9503
rect 36495 9469 36504 9503
rect 36452 9460 36504 9469
rect 28724 9324 28776 9376
rect 30656 9324 30708 9376
rect 32588 9367 32640 9376
rect 32588 9333 32597 9367
rect 32597 9333 32631 9367
rect 32631 9333 32640 9367
rect 32588 9324 32640 9333
rect 33232 9324 33284 9376
rect 33508 9324 33560 9376
rect 34704 9367 34756 9376
rect 34704 9333 34713 9367
rect 34713 9333 34747 9367
rect 34747 9333 34756 9367
rect 34704 9324 34756 9333
rect 37464 9367 37516 9376
rect 37464 9333 37473 9367
rect 37473 9333 37507 9367
rect 37507 9333 37516 9367
rect 37464 9324 37516 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1676 9120 1728 9172
rect 2504 9120 2556 9172
rect 3424 9163 3476 9172
rect 3424 9129 3433 9163
rect 3433 9129 3467 9163
rect 3467 9129 3476 9163
rect 3424 9120 3476 9129
rect 3516 9120 3568 9172
rect 4896 9120 4948 9172
rect 5540 9120 5592 9172
rect 2320 9095 2372 9104
rect 2320 9061 2329 9095
rect 2329 9061 2363 9095
rect 2363 9061 2372 9095
rect 2320 9052 2372 9061
rect 2872 9052 2924 9104
rect 3700 9052 3752 9104
rect 4252 9095 4304 9104
rect 4252 9061 4261 9095
rect 4261 9061 4295 9095
rect 4295 9061 4304 9095
rect 4252 9052 4304 9061
rect 7380 9095 7432 9104
rect 7380 9061 7389 9095
rect 7389 9061 7423 9095
rect 7423 9061 7432 9095
rect 7380 9052 7432 9061
rect 1676 8984 1728 9036
rect 5724 8984 5776 9036
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 10600 9120 10652 9172
rect 11520 9163 11572 9172
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 16120 9120 16172 9172
rect 18236 9120 18288 9172
rect 18696 9163 18748 9172
rect 18696 9129 18705 9163
rect 18705 9129 18739 9163
rect 18739 9129 18748 9163
rect 18696 9120 18748 9129
rect 20076 9163 20128 9172
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 21456 9120 21508 9172
rect 24400 9163 24452 9172
rect 24400 9129 24409 9163
rect 24409 9129 24443 9163
rect 24443 9129 24452 9163
rect 24400 9120 24452 9129
rect 26700 9120 26752 9172
rect 28632 9163 28684 9172
rect 28632 9129 28641 9163
rect 28641 9129 28675 9163
rect 28675 9129 28684 9163
rect 28632 9120 28684 9129
rect 33048 9120 33100 9172
rect 33324 9120 33376 9172
rect 34704 9120 34756 9172
rect 38660 9120 38712 9172
rect 11888 9052 11940 9104
rect 13452 9052 13504 9104
rect 17408 9052 17460 9104
rect 18052 9052 18104 9104
rect 18880 9052 18932 9104
rect 21272 9095 21324 9104
rect 10416 8984 10468 9036
rect 10692 8984 10744 9036
rect 14832 8984 14884 9036
rect 17776 8984 17828 9036
rect 21272 9061 21281 9095
rect 21281 9061 21315 9095
rect 21315 9061 21324 9095
rect 21272 9052 21324 9061
rect 21364 9095 21416 9104
rect 21364 9061 21373 9095
rect 21373 9061 21407 9095
rect 21407 9061 21416 9095
rect 27344 9095 27396 9104
rect 21364 9052 21416 9061
rect 27344 9061 27353 9095
rect 27353 9061 27387 9095
rect 27387 9061 27396 9095
rect 27344 9052 27396 9061
rect 27528 9052 27580 9104
rect 27712 9052 27764 9104
rect 29000 9095 29052 9104
rect 29000 9061 29009 9095
rect 29009 9061 29043 9095
rect 29043 9061 29052 9095
rect 29000 9052 29052 9061
rect 34152 9052 34204 9104
rect 35624 9095 35676 9104
rect 35624 9061 35633 9095
rect 35633 9061 35667 9095
rect 35667 9061 35676 9095
rect 35624 9052 35676 9061
rect 3608 8916 3660 8968
rect 4804 8916 4856 8968
rect 4988 8916 5040 8968
rect 6092 8959 6144 8968
rect 3056 8848 3108 8900
rect 4620 8848 4672 8900
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 11980 8959 12032 8968
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 13084 8916 13136 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 8576 8848 8628 8900
rect 9036 8848 9088 8900
rect 11612 8848 11664 8900
rect 13636 8848 13688 8900
rect 20168 8984 20220 9036
rect 22744 9027 22796 9036
rect 22744 8993 22753 9027
rect 22753 8993 22787 9027
rect 22787 8993 22796 9027
rect 22744 8984 22796 8993
rect 23940 8984 23992 9036
rect 24124 8984 24176 9036
rect 25228 8984 25280 9036
rect 25412 9027 25464 9036
rect 25412 8993 25421 9027
rect 25421 8993 25455 9027
rect 25455 8993 25464 9027
rect 25412 8984 25464 8993
rect 30380 9027 30432 9036
rect 30380 8993 30389 9027
rect 30389 8993 30423 9027
rect 30423 8993 30432 9027
rect 30380 8984 30432 8993
rect 32312 9027 32364 9036
rect 32312 8993 32321 9027
rect 32321 8993 32355 9027
rect 32355 8993 32364 9027
rect 32312 8984 32364 8993
rect 32680 9027 32732 9036
rect 32680 8993 32689 9027
rect 32689 8993 32723 9027
rect 32723 8993 32732 9027
rect 32680 8984 32732 8993
rect 1768 8780 1820 8832
rect 4436 8780 4488 8832
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 8760 8780 8812 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 16304 8780 16356 8832
rect 16672 8780 16724 8832
rect 19248 8916 19300 8968
rect 21732 8916 21784 8968
rect 22192 8916 22244 8968
rect 25596 8959 25648 8968
rect 25596 8925 25605 8959
rect 25605 8925 25639 8959
rect 25639 8925 25648 8959
rect 25596 8916 25648 8925
rect 28080 8916 28132 8968
rect 28540 8916 28592 8968
rect 28632 8916 28684 8968
rect 29184 8959 29236 8968
rect 29184 8925 29193 8959
rect 29193 8925 29227 8959
rect 29227 8925 29236 8959
rect 29184 8916 29236 8925
rect 32864 8959 32916 8968
rect 32864 8925 32873 8959
rect 32873 8925 32907 8959
rect 32907 8925 32916 8959
rect 32864 8916 32916 8925
rect 33232 8916 33284 8968
rect 33968 8959 34020 8968
rect 33968 8925 33977 8959
rect 33977 8925 34011 8959
rect 34011 8925 34020 8959
rect 33968 8916 34020 8925
rect 34060 8916 34112 8968
rect 35348 8916 35400 8968
rect 36268 8916 36320 8968
rect 19984 8848 20036 8900
rect 23388 8848 23440 8900
rect 26700 8848 26752 8900
rect 36820 8848 36872 8900
rect 21456 8780 21508 8832
rect 23112 8780 23164 8832
rect 24400 8780 24452 8832
rect 27160 8823 27212 8832
rect 27160 8789 27169 8823
rect 27169 8789 27203 8823
rect 27203 8789 27212 8823
rect 27160 8780 27212 8789
rect 31392 8780 31444 8832
rect 33140 8780 33192 8832
rect 33324 8780 33376 8832
rect 34980 8823 35032 8832
rect 34980 8789 34989 8823
rect 34989 8789 35023 8823
rect 35023 8789 35032 8823
rect 34980 8780 35032 8789
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 3700 8508 3752 8560
rect 4252 8576 4304 8628
rect 4804 8576 4856 8628
rect 7380 8576 7432 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 8668 8619 8720 8628
rect 8668 8585 8677 8619
rect 8677 8585 8711 8619
rect 8711 8585 8720 8619
rect 8668 8576 8720 8585
rect 10692 8576 10744 8628
rect 4436 8508 4488 8560
rect 7288 8508 7340 8560
rect 1584 8440 1636 8492
rect 1860 8440 1912 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 10416 8551 10468 8560
rect 10416 8517 10425 8551
rect 10425 8517 10459 8551
rect 10459 8517 10468 8551
rect 10416 8508 10468 8517
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 3056 8347 3108 8356
rect 1584 8304 1636 8313
rect 3056 8313 3065 8347
rect 3065 8313 3099 8347
rect 3099 8313 3108 8347
rect 3056 8304 3108 8313
rect 5356 8347 5408 8356
rect 2872 8279 2924 8288
rect 2872 8245 2881 8279
rect 2881 8245 2915 8279
rect 2915 8245 2924 8279
rect 2872 8236 2924 8245
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 8668 8372 8720 8424
rect 11520 8576 11572 8628
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 19616 8576 19668 8628
rect 21272 8576 21324 8628
rect 22744 8619 22796 8628
rect 22744 8585 22753 8619
rect 22753 8585 22787 8619
rect 22787 8585 22796 8619
rect 22744 8576 22796 8585
rect 23940 8619 23992 8628
rect 23940 8585 23949 8619
rect 23949 8585 23983 8619
rect 23983 8585 23992 8619
rect 23940 8576 23992 8585
rect 25228 8576 25280 8628
rect 27804 8576 27856 8628
rect 29000 8576 29052 8628
rect 32680 8576 32732 8628
rect 35624 8576 35676 8628
rect 36268 8619 36320 8628
rect 36268 8585 36277 8619
rect 36277 8585 36311 8619
rect 36311 8585 36320 8619
rect 36268 8576 36320 8585
rect 36636 8619 36688 8628
rect 36636 8585 36645 8619
rect 36645 8585 36679 8619
rect 36679 8585 36688 8619
rect 36636 8576 36688 8585
rect 13084 8508 13136 8560
rect 17776 8508 17828 8560
rect 19064 8508 19116 8560
rect 19248 8551 19300 8560
rect 19248 8517 19257 8551
rect 19257 8517 19291 8551
rect 19291 8517 19300 8551
rect 19248 8508 19300 8517
rect 20260 8508 20312 8560
rect 28448 8508 28500 8560
rect 35900 8508 35952 8560
rect 11980 8440 12032 8492
rect 16488 8440 16540 8492
rect 18052 8440 18104 8492
rect 19708 8440 19760 8492
rect 20076 8440 20128 8492
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 21732 8440 21784 8492
rect 27712 8483 27764 8492
rect 15200 8415 15252 8424
rect 10968 8347 11020 8356
rect 10968 8313 10977 8347
rect 10977 8313 11011 8347
rect 11011 8313 11020 8347
rect 10968 8304 11020 8313
rect 12348 8304 12400 8356
rect 3424 8236 3476 8288
rect 4252 8236 4304 8288
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 5724 8236 5776 8288
rect 7288 8236 7340 8288
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 11980 8236 12032 8288
rect 12900 8304 12952 8356
rect 13084 8236 13136 8288
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 16856 8372 16908 8424
rect 14648 8304 14700 8356
rect 18420 8347 18472 8356
rect 18420 8313 18429 8347
rect 18429 8313 18463 8347
rect 18463 8313 18472 8347
rect 18420 8304 18472 8313
rect 14740 8236 14792 8288
rect 15660 8236 15712 8288
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 16948 8236 17000 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 19616 8279 19668 8288
rect 19616 8245 19625 8279
rect 19625 8245 19659 8279
rect 19659 8245 19668 8279
rect 21272 8372 21324 8424
rect 23388 8372 23440 8424
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 29184 8440 29236 8492
rect 33324 8483 33376 8492
rect 33324 8449 33333 8483
rect 33333 8449 33367 8483
rect 33367 8449 33376 8483
rect 33324 8440 33376 8449
rect 34060 8440 34112 8492
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 24308 8415 24360 8424
rect 24308 8381 24317 8415
rect 24317 8381 24351 8415
rect 24351 8381 24360 8415
rect 24308 8372 24360 8381
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 25872 8415 25924 8424
rect 25872 8381 25881 8415
rect 25881 8381 25915 8415
rect 25915 8381 25924 8415
rect 25872 8372 25924 8381
rect 31392 8372 31444 8424
rect 33140 8372 33192 8424
rect 21548 8347 21600 8356
rect 21548 8313 21557 8347
rect 21557 8313 21591 8347
rect 21591 8313 21600 8347
rect 21548 8304 21600 8313
rect 22192 8304 22244 8356
rect 27804 8347 27856 8356
rect 20812 8279 20864 8288
rect 19616 8236 19668 8245
rect 20812 8245 20821 8279
rect 20821 8245 20855 8279
rect 20855 8245 20864 8279
rect 20812 8236 20864 8245
rect 27804 8313 27813 8347
rect 27813 8313 27847 8347
rect 27847 8313 27856 8347
rect 27804 8304 27856 8313
rect 28540 8304 28592 8356
rect 29368 8347 29420 8356
rect 29368 8313 29377 8347
rect 29377 8313 29411 8347
rect 29411 8313 29420 8347
rect 29368 8304 29420 8313
rect 26792 8236 26844 8288
rect 26976 8236 27028 8288
rect 27528 8236 27580 8288
rect 32588 8304 32640 8356
rect 34612 8304 34664 8356
rect 30380 8279 30432 8288
rect 30380 8245 30389 8279
rect 30389 8245 30423 8279
rect 30423 8245 30432 8279
rect 30380 8236 30432 8245
rect 32312 8236 32364 8288
rect 34244 8279 34296 8288
rect 34244 8245 34253 8279
rect 34253 8245 34287 8279
rect 34287 8245 34296 8279
rect 34244 8236 34296 8245
rect 34520 8236 34572 8288
rect 38016 8415 38068 8424
rect 38016 8381 38025 8415
rect 38025 8381 38059 8415
rect 38059 8381 38068 8415
rect 38016 8372 38068 8381
rect 37372 8236 37424 8288
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 1584 8032 1636 8084
rect 2872 8032 2924 8084
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3608 8032 3660 8084
rect 6736 8032 6788 8084
rect 6920 8032 6972 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 8944 8032 8996 8084
rect 10600 8032 10652 8084
rect 10968 8032 11020 8084
rect 12532 8032 12584 8084
rect 14832 8032 14884 8084
rect 15660 8075 15712 8084
rect 15660 8041 15669 8075
rect 15669 8041 15703 8075
rect 15703 8041 15712 8075
rect 15660 8032 15712 8041
rect 17408 8032 17460 8084
rect 19248 8032 19300 8084
rect 19708 8032 19760 8084
rect 22100 8075 22152 8084
rect 22100 8041 22109 8075
rect 22109 8041 22143 8075
rect 22143 8041 22152 8075
rect 22100 8032 22152 8041
rect 22192 8032 22244 8084
rect 23756 8032 23808 8084
rect 24308 8075 24360 8084
rect 24308 8041 24317 8075
rect 24317 8041 24351 8075
rect 24351 8041 24360 8075
rect 24308 8032 24360 8041
rect 25872 8075 25924 8084
rect 25872 8041 25881 8075
rect 25881 8041 25915 8075
rect 25915 8041 25924 8075
rect 25872 8032 25924 8041
rect 26792 8032 26844 8084
rect 27436 8075 27488 8084
rect 27436 8041 27445 8075
rect 27445 8041 27479 8075
rect 27479 8041 27488 8075
rect 27436 8032 27488 8041
rect 27988 8032 28040 8084
rect 1676 8007 1728 8016
rect 1676 7973 1685 8007
rect 1685 7973 1719 8007
rect 1719 7973 1728 8007
rect 1676 7964 1728 7973
rect 2320 7964 2372 8016
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 5264 7964 5316 8016
rect 2228 7896 2280 7948
rect 4896 7896 4948 7948
rect 7288 7964 7340 8016
rect 4344 7828 4396 7880
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 11152 7964 11204 8016
rect 12900 8007 12952 8016
rect 12900 7973 12909 8007
rect 12909 7973 12943 8007
rect 12943 7973 12952 8007
rect 12900 7964 12952 7973
rect 13544 7964 13596 8016
rect 16488 8007 16540 8016
rect 16488 7973 16497 8007
rect 16497 7973 16531 8007
rect 16531 7973 16540 8007
rect 16488 7964 16540 7973
rect 17132 8007 17184 8016
rect 17132 7973 17141 8007
rect 17141 7973 17175 8007
rect 17175 7973 17184 8007
rect 17132 7964 17184 7973
rect 17224 8007 17276 8016
rect 17224 7973 17233 8007
rect 17233 7973 17267 8007
rect 17267 7973 17276 8007
rect 17776 8007 17828 8016
rect 17224 7964 17276 7973
rect 17776 7973 17785 8007
rect 17785 7973 17819 8007
rect 17819 7973 17828 8007
rect 17776 7964 17828 7973
rect 21272 8007 21324 8016
rect 21272 7973 21281 8007
rect 21281 7973 21315 8007
rect 21315 7973 21324 8007
rect 21272 7964 21324 7973
rect 22836 8007 22888 8016
rect 22836 7973 22845 8007
rect 22845 7973 22879 8007
rect 22879 7973 22888 8007
rect 22836 7964 22888 7973
rect 25228 7964 25280 8016
rect 12348 7896 12400 7948
rect 15016 7896 15068 7948
rect 18696 7896 18748 7948
rect 20812 7896 20864 7948
rect 24676 7896 24728 7948
rect 25412 7939 25464 7948
rect 25412 7905 25421 7939
rect 25421 7905 25455 7939
rect 25455 7905 25464 7939
rect 25412 7896 25464 7905
rect 27344 7964 27396 8016
rect 28632 8007 28684 8016
rect 28632 7973 28641 8007
rect 28641 7973 28675 8007
rect 28675 7973 28684 8007
rect 28632 7964 28684 7973
rect 33508 8032 33560 8084
rect 33968 8032 34020 8084
rect 34428 8032 34480 8084
rect 35900 8075 35952 8084
rect 32588 7964 32640 8016
rect 33048 7964 33100 8016
rect 34244 7964 34296 8016
rect 34704 7964 34756 8016
rect 35900 8041 35909 8075
rect 35909 8041 35943 8075
rect 35943 8041 35952 8075
rect 35900 8032 35952 8041
rect 38016 7964 38068 8016
rect 30472 7939 30524 7948
rect 30472 7905 30481 7939
rect 30481 7905 30515 7939
rect 30515 7905 30524 7939
rect 30472 7896 30524 7905
rect 31300 7896 31352 7948
rect 11704 7828 11756 7880
rect 12624 7828 12676 7880
rect 14740 7828 14792 7880
rect 19984 7828 20036 7880
rect 21824 7828 21876 7880
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 24124 7828 24176 7880
rect 24768 7871 24820 7880
rect 24768 7837 24777 7871
rect 24777 7837 24811 7871
rect 24811 7837 24820 7871
rect 24768 7828 24820 7837
rect 27620 7828 27672 7880
rect 28540 7871 28592 7880
rect 28540 7837 28549 7871
rect 28549 7837 28583 7871
rect 28583 7837 28592 7871
rect 28540 7828 28592 7837
rect 30012 7828 30064 7880
rect 32496 7828 32548 7880
rect 5816 7803 5868 7812
rect 5816 7769 5825 7803
rect 5825 7769 5859 7803
rect 5859 7769 5868 7803
rect 5816 7760 5868 7769
rect 6368 7760 6420 7812
rect 9128 7760 9180 7812
rect 9956 7760 10008 7812
rect 13084 7760 13136 7812
rect 16856 7803 16908 7812
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5264 7692 5316 7701
rect 5908 7692 5960 7744
rect 6644 7692 6696 7744
rect 8668 7735 8720 7744
rect 8668 7701 8677 7735
rect 8677 7701 8711 7735
rect 8711 7701 8720 7735
rect 8668 7692 8720 7701
rect 13544 7692 13596 7744
rect 16856 7769 16865 7803
rect 16865 7769 16899 7803
rect 16899 7769 16908 7803
rect 16856 7760 16908 7769
rect 24584 7760 24636 7812
rect 30288 7760 30340 7812
rect 30380 7760 30432 7812
rect 34152 7896 34204 7948
rect 36452 7939 36504 7948
rect 36452 7905 36461 7939
rect 36461 7905 36495 7939
rect 36495 7905 36504 7939
rect 36452 7896 36504 7905
rect 34980 7871 35032 7880
rect 34980 7837 34989 7871
rect 34989 7837 35023 7871
rect 35023 7837 35032 7871
rect 34980 7828 35032 7837
rect 35624 7871 35676 7880
rect 35624 7837 35633 7871
rect 35633 7837 35667 7871
rect 35667 7837 35676 7871
rect 35624 7828 35676 7837
rect 36360 7760 36412 7812
rect 36636 7803 36688 7812
rect 36636 7769 36645 7803
rect 36645 7769 36679 7803
rect 36679 7769 36688 7803
rect 36636 7760 36688 7769
rect 18420 7692 18472 7744
rect 18880 7692 18932 7744
rect 27528 7692 27580 7744
rect 29368 7692 29420 7744
rect 33048 7735 33100 7744
rect 33048 7701 33057 7735
rect 33057 7701 33091 7735
rect 33091 7701 33100 7735
rect 33048 7692 33100 7701
rect 34980 7692 35032 7744
rect 36820 7692 36872 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 3332 7488 3384 7540
rect 4252 7488 4304 7540
rect 5264 7488 5316 7540
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 12900 7488 12952 7540
rect 15660 7488 15712 7540
rect 16948 7488 17000 7540
rect 17132 7488 17184 7540
rect 19616 7488 19668 7540
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 21916 7488 21968 7540
rect 24676 7488 24728 7540
rect 26976 7531 27028 7540
rect 26976 7497 26985 7531
rect 26985 7497 27019 7531
rect 27019 7497 27028 7531
rect 26976 7488 27028 7497
rect 27620 7531 27672 7540
rect 27620 7497 27629 7531
rect 27629 7497 27663 7531
rect 27663 7497 27672 7531
rect 27620 7488 27672 7497
rect 28632 7531 28684 7540
rect 28632 7497 28641 7531
rect 28641 7497 28675 7531
rect 28675 7497 28684 7531
rect 28632 7488 28684 7497
rect 32496 7531 32548 7540
rect 32496 7497 32505 7531
rect 32505 7497 32539 7531
rect 32539 7497 32548 7531
rect 32496 7488 32548 7497
rect 33048 7531 33100 7540
rect 33048 7497 33057 7531
rect 33057 7497 33091 7531
rect 33091 7497 33100 7531
rect 33048 7488 33100 7497
rect 34152 7488 34204 7540
rect 36452 7488 36504 7540
rect 2228 7420 2280 7472
rect 3884 7420 3936 7472
rect 9496 7420 9548 7472
rect 12624 7420 12676 7472
rect 1676 7352 1728 7404
rect 3148 7284 3200 7336
rect 4068 7352 4120 7404
rect 6000 7352 6052 7404
rect 6368 7352 6420 7404
rect 8300 7352 8352 7404
rect 9220 7352 9272 7404
rect 10508 7352 10560 7404
rect 12164 7352 12216 7404
rect 5356 7259 5408 7268
rect 5356 7225 5365 7259
rect 5365 7225 5399 7259
rect 5399 7225 5408 7259
rect 5908 7259 5960 7268
rect 5356 7216 5408 7225
rect 5908 7225 5917 7259
rect 5917 7225 5951 7259
rect 5951 7225 5960 7259
rect 5908 7216 5960 7225
rect 2228 7148 2280 7200
rect 3976 7148 4028 7200
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 11612 7284 11664 7336
rect 7288 7216 7340 7268
rect 8484 7259 8536 7268
rect 8484 7225 8493 7259
rect 8493 7225 8527 7259
rect 8527 7225 8536 7259
rect 8484 7216 8536 7225
rect 9128 7216 9180 7268
rect 8116 7148 8168 7200
rect 11152 7148 11204 7200
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 14740 7284 14792 7336
rect 17776 7420 17828 7472
rect 20536 7420 20588 7472
rect 22744 7420 22796 7472
rect 27160 7420 27212 7472
rect 28908 7420 28960 7472
rect 16488 7352 16540 7404
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 18144 7352 18196 7404
rect 19892 7352 19944 7404
rect 22100 7352 22152 7404
rect 23756 7395 23808 7404
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 23756 7352 23808 7361
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 25596 7352 25648 7404
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 26332 7352 26384 7404
rect 26792 7352 26844 7404
rect 29184 7352 29236 7404
rect 25412 7284 25464 7336
rect 16028 7216 16080 7268
rect 16120 7259 16172 7268
rect 16120 7225 16129 7259
rect 16129 7225 16163 7259
rect 16163 7225 16172 7259
rect 17868 7259 17920 7268
rect 16120 7216 16172 7225
rect 17868 7225 17877 7259
rect 17877 7225 17911 7259
rect 17911 7225 17920 7259
rect 17868 7216 17920 7225
rect 19248 7216 19300 7268
rect 12900 7191 12952 7200
rect 12164 7148 12216 7157
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 17132 7191 17184 7200
rect 17132 7157 17141 7191
rect 17141 7157 17175 7191
rect 17175 7157 17184 7191
rect 17132 7148 17184 7157
rect 19340 7191 19392 7200
rect 19340 7157 19349 7191
rect 19349 7157 19383 7191
rect 19383 7157 19392 7191
rect 19340 7148 19392 7157
rect 21916 7259 21968 7268
rect 21916 7225 21925 7259
rect 21925 7225 21959 7259
rect 21959 7225 21968 7259
rect 22836 7259 22888 7268
rect 21916 7216 21968 7225
rect 22836 7225 22845 7259
rect 22845 7225 22879 7259
rect 22879 7225 22888 7259
rect 22836 7216 22888 7225
rect 23756 7216 23808 7268
rect 22560 7148 22612 7200
rect 23204 7148 23256 7200
rect 26332 7216 26384 7268
rect 28264 7327 28316 7336
rect 28264 7293 28273 7327
rect 28273 7293 28307 7327
rect 28307 7293 28316 7327
rect 28264 7284 28316 7293
rect 34612 7420 34664 7472
rect 31392 7395 31444 7404
rect 31392 7361 31401 7395
rect 31401 7361 31435 7395
rect 31435 7361 31444 7395
rect 31392 7352 31444 7361
rect 33508 7352 33560 7404
rect 35900 7352 35952 7404
rect 31300 7327 31352 7336
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 28448 7216 28500 7268
rect 29460 7259 29512 7268
rect 29460 7225 29469 7259
rect 29469 7225 29503 7259
rect 29503 7225 29512 7259
rect 30012 7259 30064 7268
rect 29460 7216 29512 7225
rect 30012 7225 30021 7259
rect 30021 7225 30055 7259
rect 30055 7225 30064 7259
rect 30012 7216 30064 7225
rect 33048 7216 33100 7268
rect 25872 7191 25924 7200
rect 25872 7157 25881 7191
rect 25881 7157 25915 7191
rect 25915 7157 25924 7191
rect 25872 7148 25924 7157
rect 30288 7191 30340 7200
rect 30288 7157 30297 7191
rect 30297 7157 30331 7191
rect 30331 7157 30340 7191
rect 30288 7148 30340 7157
rect 30472 7148 30524 7200
rect 32496 7148 32548 7200
rect 34980 7216 35032 7268
rect 35624 7259 35676 7268
rect 34704 7191 34756 7200
rect 34704 7157 34713 7191
rect 34713 7157 34747 7191
rect 34747 7157 34756 7191
rect 34704 7148 34756 7157
rect 34796 7148 34848 7200
rect 35624 7225 35633 7259
rect 35633 7225 35667 7259
rect 35667 7225 35676 7259
rect 35624 7216 35676 7225
rect 36360 7352 36412 7404
rect 36820 7395 36872 7404
rect 36820 7361 36829 7395
rect 36829 7361 36863 7395
rect 36863 7361 36872 7395
rect 36820 7352 36872 7361
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 1860 6944 1912 6996
rect 2136 6987 2188 6996
rect 2136 6953 2145 6987
rect 2145 6953 2179 6987
rect 2179 6953 2188 6987
rect 2136 6944 2188 6953
rect 2228 6944 2280 6996
rect 2872 6944 2924 6996
rect 4344 6987 4396 6996
rect 4344 6953 4353 6987
rect 4353 6953 4387 6987
rect 4387 6953 4396 6987
rect 4344 6944 4396 6953
rect 5356 6944 5408 6996
rect 6000 6987 6052 6996
rect 6000 6953 6009 6987
rect 6009 6953 6043 6987
rect 6043 6953 6052 6987
rect 6000 6944 6052 6953
rect 8300 6944 8352 6996
rect 10508 6944 10560 6996
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 14740 6944 14792 6996
rect 15016 6944 15068 6996
rect 16396 6944 16448 6996
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 18696 6944 18748 6996
rect 19892 6944 19944 6996
rect 22560 6944 22612 6996
rect 23204 6987 23256 6996
rect 23204 6953 23213 6987
rect 23213 6953 23247 6987
rect 23247 6953 23256 6987
rect 23204 6944 23256 6953
rect 23756 6944 23808 6996
rect 26056 6987 26108 6996
rect 26056 6953 26065 6987
rect 26065 6953 26099 6987
rect 26099 6953 26108 6987
rect 26056 6944 26108 6953
rect 27528 6944 27580 6996
rect 28540 6944 28592 6996
rect 28632 6944 28684 6996
rect 29184 6944 29236 6996
rect 29460 6944 29512 6996
rect 30656 6944 30708 6996
rect 31576 6944 31628 6996
rect 34152 6987 34204 6996
rect 34152 6953 34161 6987
rect 34161 6953 34195 6987
rect 34195 6953 34204 6987
rect 34152 6944 34204 6953
rect 34704 6944 34756 6996
rect 3056 6876 3108 6928
rect 4712 6876 4764 6928
rect 6368 6919 6420 6928
rect 6368 6885 6377 6919
rect 6377 6885 6411 6919
rect 6411 6885 6420 6919
rect 6368 6876 6420 6885
rect 7472 6876 7524 6928
rect 8024 6876 8076 6928
rect 8484 6876 8536 6928
rect 11152 6876 11204 6928
rect 12900 6876 12952 6928
rect 13544 6919 13596 6928
rect 13544 6885 13553 6919
rect 13553 6885 13587 6919
rect 13587 6885 13596 6919
rect 13544 6876 13596 6885
rect 16948 6876 17000 6928
rect 17868 6876 17920 6928
rect 18880 6919 18932 6928
rect 18880 6885 18889 6919
rect 18889 6885 18923 6919
rect 18923 6885 18932 6919
rect 18880 6876 18932 6885
rect 18972 6876 19024 6928
rect 22468 6876 22520 6928
rect 24400 6876 24452 6928
rect 28816 6876 28868 6928
rect 35440 6919 35492 6928
rect 35440 6885 35449 6919
rect 35449 6885 35483 6919
rect 35483 6885 35492 6919
rect 35440 6876 35492 6885
rect 35992 6876 36044 6928
rect 36360 6876 36412 6928
rect 2044 6808 2096 6860
rect 5908 6808 5960 6860
rect 9588 6808 9640 6860
rect 11060 6851 11112 6860
rect 11060 6817 11069 6851
rect 11069 6817 11103 6851
rect 11103 6817 11112 6851
rect 11060 6808 11112 6817
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 15476 6808 15528 6860
rect 16580 6808 16632 6860
rect 20260 6808 20312 6860
rect 5448 6740 5500 6792
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 12440 6740 12492 6792
rect 8208 6672 8260 6724
rect 10232 6715 10284 6724
rect 10232 6681 10241 6715
rect 10241 6681 10275 6715
rect 10275 6681 10284 6715
rect 13360 6740 13412 6792
rect 15384 6740 15436 6792
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 20720 6740 20772 6792
rect 22744 6808 22796 6860
rect 26608 6808 26660 6860
rect 32128 6851 32180 6860
rect 32128 6817 32137 6851
rect 32137 6817 32171 6851
rect 32171 6817 32180 6851
rect 32128 6808 32180 6817
rect 32680 6851 32732 6860
rect 32680 6817 32689 6851
rect 32689 6817 32723 6851
rect 32723 6817 32732 6851
rect 32680 6808 32732 6817
rect 34612 6808 34664 6860
rect 22376 6740 22428 6792
rect 10232 6672 10284 6681
rect 13636 6672 13688 6724
rect 27804 6783 27856 6792
rect 27804 6749 27813 6783
rect 27813 6749 27847 6783
rect 27847 6749 27856 6783
rect 27804 6740 27856 6749
rect 29552 6783 29604 6792
rect 29552 6749 29561 6783
rect 29561 6749 29595 6783
rect 29595 6749 29604 6783
rect 29552 6740 29604 6749
rect 31300 6740 31352 6792
rect 33784 6783 33836 6792
rect 33784 6749 33793 6783
rect 33793 6749 33827 6783
rect 33827 6749 33836 6783
rect 33784 6740 33836 6749
rect 35256 6740 35308 6792
rect 112 6604 164 6656
rect 3516 6604 3568 6656
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 9036 6604 9088 6656
rect 9496 6604 9548 6656
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 17132 6604 17184 6656
rect 17868 6604 17920 6656
rect 20168 6604 20220 6656
rect 22284 6604 22336 6656
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 27528 6604 27580 6656
rect 33324 6647 33376 6656
rect 33324 6613 33333 6647
rect 33333 6613 33367 6647
rect 33367 6613 33376 6647
rect 33324 6604 33376 6613
rect 34796 6604 34848 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 2044 6400 2096 6452
rect 2136 6264 2188 6316
rect 4896 6400 4948 6452
rect 6276 6400 6328 6452
rect 4620 6332 4672 6384
rect 6368 6332 6420 6384
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 6552 6264 6604 6316
rect 6000 6196 6052 6248
rect 9956 6400 10008 6452
rect 11060 6400 11112 6452
rect 12900 6400 12952 6452
rect 16580 6400 16632 6452
rect 18880 6400 18932 6452
rect 19800 6443 19852 6452
rect 19800 6409 19809 6443
rect 19809 6409 19843 6443
rect 19843 6409 19852 6443
rect 19800 6400 19852 6409
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 13912 6332 13964 6384
rect 18788 6332 18840 6384
rect 12532 6307 12584 6316
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 12532 6273 12541 6307
rect 12541 6273 12575 6307
rect 12575 6273 12584 6307
rect 12532 6264 12584 6273
rect 13544 6264 13596 6316
rect 16396 6264 16448 6316
rect 24400 6400 24452 6452
rect 26884 6400 26936 6452
rect 32312 6400 32364 6452
rect 32680 6400 32732 6452
rect 34152 6400 34204 6452
rect 35992 6443 36044 6452
rect 35992 6409 36001 6443
rect 36001 6409 36035 6443
rect 36035 6409 36044 6443
rect 35992 6400 36044 6409
rect 24676 6332 24728 6384
rect 32128 6375 32180 6384
rect 22376 6307 22428 6316
rect 22376 6273 22385 6307
rect 22385 6273 22419 6307
rect 22419 6273 22428 6307
rect 22376 6264 22428 6273
rect 24860 6264 24912 6316
rect 25228 6307 25280 6316
rect 25228 6273 25237 6307
rect 25237 6273 25271 6307
rect 25271 6273 25280 6307
rect 25228 6264 25280 6273
rect 26608 6264 26660 6316
rect 27528 6264 27580 6316
rect 9220 6196 9272 6205
rect 10232 6239 10284 6248
rect 10232 6205 10241 6239
rect 10241 6205 10275 6239
rect 10275 6205 10284 6239
rect 10232 6196 10284 6205
rect 2228 6128 2280 6180
rect 4160 6128 4212 6180
rect 5356 6171 5408 6180
rect 5356 6137 5365 6171
rect 5365 6137 5399 6171
rect 5399 6137 5408 6171
rect 5356 6128 5408 6137
rect 5540 6128 5592 6180
rect 2964 6103 3016 6112
rect 2964 6069 2973 6103
rect 2973 6069 3007 6103
rect 3007 6069 3016 6103
rect 2964 6060 3016 6069
rect 3792 6060 3844 6112
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 6276 6060 6328 6112
rect 8024 6128 8076 6180
rect 8300 6171 8352 6180
rect 8300 6137 8309 6171
rect 8309 6137 8343 6171
rect 8343 6137 8352 6171
rect 8300 6128 8352 6137
rect 10508 6128 10560 6180
rect 13360 6196 13412 6248
rect 22100 6239 22152 6248
rect 22100 6205 22109 6239
rect 22109 6205 22143 6239
rect 22143 6205 22152 6239
rect 22100 6196 22152 6205
rect 22284 6239 22336 6248
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 14004 6171 14056 6180
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 14004 6137 14013 6171
rect 14013 6137 14047 6171
rect 14047 6137 14056 6171
rect 14004 6128 14056 6137
rect 16212 6128 16264 6180
rect 16948 6128 17000 6180
rect 17868 6171 17920 6180
rect 17868 6137 17877 6171
rect 17877 6137 17911 6171
rect 17911 6137 17920 6171
rect 18788 6171 18840 6180
rect 17868 6128 17920 6137
rect 12164 6060 12216 6069
rect 15476 6060 15528 6112
rect 18788 6137 18797 6171
rect 18797 6137 18831 6171
rect 18831 6137 18840 6171
rect 18788 6128 18840 6137
rect 19432 6171 19484 6180
rect 19432 6137 19441 6171
rect 19441 6137 19475 6171
rect 19475 6137 19484 6171
rect 19432 6128 19484 6137
rect 19524 6060 19576 6112
rect 20260 6060 20312 6112
rect 20444 6171 20496 6180
rect 20444 6137 20453 6171
rect 20453 6137 20487 6171
rect 20487 6137 20496 6171
rect 20996 6171 21048 6180
rect 20444 6128 20496 6137
rect 20996 6137 21005 6171
rect 21005 6137 21039 6171
rect 21039 6137 21048 6171
rect 20996 6128 21048 6137
rect 23756 6196 23808 6248
rect 24768 6196 24820 6248
rect 29736 6239 29788 6248
rect 29736 6205 29745 6239
rect 29745 6205 29779 6239
rect 29779 6205 29788 6239
rect 29736 6196 29788 6205
rect 32128 6341 32137 6375
rect 32137 6341 32171 6375
rect 32171 6341 32180 6375
rect 32128 6332 32180 6341
rect 35072 6332 35124 6384
rect 33324 6307 33376 6316
rect 33324 6273 33333 6307
rect 33333 6273 33367 6307
rect 33367 6273 33376 6307
rect 33324 6264 33376 6273
rect 33692 6264 33744 6316
rect 35440 6264 35492 6316
rect 31208 6196 31260 6248
rect 31576 6239 31628 6248
rect 31576 6205 31585 6239
rect 31585 6205 31619 6239
rect 31619 6205 31628 6239
rect 31576 6196 31628 6205
rect 25412 6128 25464 6180
rect 20720 6060 20772 6112
rect 22560 6060 22612 6112
rect 22744 6060 22796 6112
rect 23480 6103 23532 6112
rect 23480 6069 23489 6103
rect 23489 6069 23523 6103
rect 23523 6069 23532 6103
rect 23480 6060 23532 6069
rect 25872 6060 25924 6112
rect 26148 6103 26200 6112
rect 26148 6069 26157 6103
rect 26157 6069 26191 6103
rect 26191 6069 26200 6103
rect 26148 6060 26200 6069
rect 26884 6128 26936 6180
rect 27252 6128 27304 6180
rect 27804 6128 27856 6180
rect 31852 6171 31904 6180
rect 28816 6060 28868 6112
rect 31852 6137 31861 6171
rect 31861 6137 31895 6171
rect 31895 6137 31904 6171
rect 31852 6128 31904 6137
rect 30380 6103 30432 6112
rect 30380 6069 30389 6103
rect 30389 6069 30423 6103
rect 30423 6069 30432 6103
rect 30380 6060 30432 6069
rect 33048 6103 33100 6112
rect 33048 6069 33057 6103
rect 33057 6069 33091 6103
rect 33091 6069 33100 6103
rect 35992 6128 36044 6180
rect 36544 6171 36596 6180
rect 36544 6137 36553 6171
rect 36553 6137 36587 6171
rect 36587 6137 36596 6171
rect 36544 6128 36596 6137
rect 33048 6060 33100 6069
rect 35900 6060 35952 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 2688 5856 2740 5908
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 5356 5856 5408 5908
rect 7472 5899 7524 5908
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 8300 5856 8352 5908
rect 12440 5856 12492 5908
rect 13544 5856 13596 5908
rect 14648 5899 14700 5908
rect 2228 5788 2280 5840
rect 4160 5788 4212 5840
rect 5264 5788 5316 5840
rect 6276 5831 6328 5840
rect 6276 5797 6285 5831
rect 6285 5797 6319 5831
rect 6319 5797 6328 5831
rect 6276 5788 6328 5797
rect 7288 5788 7340 5840
rect 1952 5763 2004 5772
rect 1952 5729 1961 5763
rect 1961 5729 1995 5763
rect 1995 5729 2004 5763
rect 1952 5720 2004 5729
rect 4620 5720 4672 5772
rect 5356 5763 5408 5772
rect 5356 5729 5365 5763
rect 5365 5729 5399 5763
rect 5399 5729 5408 5763
rect 5356 5720 5408 5729
rect 7196 5720 7248 5772
rect 8116 5720 8168 5772
rect 10416 5788 10468 5840
rect 11152 5788 11204 5840
rect 11980 5788 12032 5840
rect 13360 5788 13412 5840
rect 14004 5788 14056 5840
rect 14648 5865 14657 5899
rect 14657 5865 14691 5899
rect 14691 5865 14700 5899
rect 14648 5856 14700 5865
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 16304 5856 16356 5908
rect 16856 5856 16908 5908
rect 17500 5788 17552 5840
rect 22376 5899 22428 5908
rect 22376 5865 22385 5899
rect 22385 5865 22419 5899
rect 22419 5865 22428 5899
rect 22376 5856 22428 5865
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 15384 5763 15436 5772
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 16028 5720 16080 5772
rect 20444 5788 20496 5840
rect 20536 5788 20588 5840
rect 21640 5831 21692 5840
rect 21640 5797 21649 5831
rect 21649 5797 21683 5831
rect 21683 5797 21692 5831
rect 21640 5788 21692 5797
rect 22652 5788 22704 5840
rect 23480 5856 23532 5908
rect 23756 5899 23808 5908
rect 23756 5865 23765 5899
rect 23765 5865 23799 5899
rect 23799 5865 23808 5899
rect 23756 5856 23808 5865
rect 24400 5899 24452 5908
rect 24400 5865 24409 5899
rect 24409 5865 24443 5899
rect 24443 5865 24452 5899
rect 24400 5856 24452 5865
rect 25228 5899 25280 5908
rect 25228 5865 25237 5899
rect 25237 5865 25271 5899
rect 25271 5865 25280 5899
rect 25228 5856 25280 5865
rect 25412 5856 25464 5908
rect 29552 5856 29604 5908
rect 33048 5856 33100 5908
rect 33784 5899 33836 5908
rect 33784 5865 33793 5899
rect 33793 5865 33827 5899
rect 33827 5865 33836 5899
rect 33784 5856 33836 5865
rect 34152 5856 34204 5908
rect 34796 5899 34848 5908
rect 34796 5865 34805 5899
rect 34805 5865 34839 5899
rect 34839 5865 34848 5899
rect 34796 5856 34848 5865
rect 36544 5856 36596 5908
rect 23848 5788 23900 5840
rect 26700 5831 26752 5840
rect 26700 5797 26709 5831
rect 26709 5797 26743 5831
rect 26743 5797 26752 5831
rect 26700 5788 26752 5797
rect 28264 5831 28316 5840
rect 28264 5797 28273 5831
rect 28273 5797 28307 5831
rect 28307 5797 28316 5831
rect 28264 5788 28316 5797
rect 30380 5788 30432 5840
rect 32496 5831 32548 5840
rect 32496 5797 32499 5831
rect 32499 5797 32533 5831
rect 32533 5797 32548 5831
rect 32496 5788 32548 5797
rect 33140 5788 33192 5840
rect 35900 5788 35952 5840
rect 2780 5652 2832 5704
rect 5448 5652 5500 5704
rect 6368 5652 6420 5704
rect 5908 5584 5960 5636
rect 10508 5652 10560 5704
rect 12256 5652 12308 5704
rect 13544 5652 13596 5704
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 19064 5695 19116 5704
rect 19064 5661 19073 5695
rect 19073 5661 19107 5695
rect 19107 5661 19116 5695
rect 19064 5652 19116 5661
rect 20996 5695 21048 5704
rect 20996 5661 21005 5695
rect 21005 5661 21039 5695
rect 21039 5661 21048 5695
rect 20996 5652 21048 5661
rect 21916 5652 21968 5704
rect 22284 5652 22336 5704
rect 32864 5720 32916 5772
rect 24032 5695 24084 5704
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 25964 5652 26016 5704
rect 27252 5695 27304 5704
rect 27252 5661 27261 5695
rect 27261 5661 27295 5695
rect 27295 5661 27304 5695
rect 27252 5652 27304 5661
rect 28172 5695 28224 5704
rect 28172 5661 28181 5695
rect 28181 5661 28215 5695
rect 28215 5661 28224 5695
rect 28172 5652 28224 5661
rect 28356 5652 28408 5704
rect 12532 5584 12584 5636
rect 13728 5584 13780 5636
rect 21824 5584 21876 5636
rect 22100 5584 22152 5636
rect 7288 5516 7340 5568
rect 10968 5559 11020 5568
rect 10968 5525 10977 5559
rect 10977 5525 11011 5559
rect 11011 5525 11020 5559
rect 10968 5516 11020 5525
rect 11336 5559 11388 5568
rect 11336 5525 11345 5559
rect 11345 5525 11379 5559
rect 11379 5525 11388 5559
rect 11336 5516 11388 5525
rect 13544 5516 13596 5568
rect 15844 5559 15896 5568
rect 15844 5525 15853 5559
rect 15853 5525 15887 5559
rect 15887 5525 15896 5559
rect 15844 5516 15896 5525
rect 19616 5559 19668 5568
rect 19616 5525 19625 5559
rect 19625 5525 19659 5559
rect 19659 5525 19668 5559
rect 19616 5516 19668 5525
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 21456 5516 21508 5568
rect 24952 5559 25004 5568
rect 24952 5525 24961 5559
rect 24961 5525 24995 5559
rect 24995 5525 25004 5559
rect 24952 5516 25004 5525
rect 26056 5516 26108 5568
rect 27068 5516 27120 5568
rect 28172 5516 28224 5568
rect 30472 5652 30524 5704
rect 31576 5652 31628 5704
rect 32404 5652 32456 5704
rect 33876 5695 33928 5704
rect 33876 5661 33885 5695
rect 33885 5661 33919 5695
rect 33919 5661 33928 5695
rect 33876 5652 33928 5661
rect 35992 5695 36044 5704
rect 35992 5661 36001 5695
rect 36001 5661 36035 5695
rect 36035 5661 36044 5695
rect 35992 5652 36044 5661
rect 28632 5516 28684 5568
rect 29736 5516 29788 5568
rect 33048 5559 33100 5568
rect 33048 5525 33057 5559
rect 33057 5525 33091 5559
rect 33091 5525 33100 5559
rect 33048 5516 33100 5525
rect 35256 5516 35308 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 1492 5312 1544 5364
rect 2964 5312 3016 5364
rect 5448 5355 5500 5364
rect 5448 5321 5457 5355
rect 5457 5321 5491 5355
rect 5491 5321 5500 5355
rect 5448 5312 5500 5321
rect 6460 5355 6512 5364
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 7196 5355 7248 5364
rect 7196 5321 7205 5355
rect 7205 5321 7239 5355
rect 7239 5321 7248 5355
rect 7196 5312 7248 5321
rect 8300 5312 8352 5364
rect 6276 5244 6328 5296
rect 3792 5176 3844 5228
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 9772 5312 9824 5364
rect 10416 5355 10468 5364
rect 10416 5321 10425 5355
rect 10425 5321 10459 5355
rect 10459 5321 10468 5355
rect 10416 5312 10468 5321
rect 12624 5355 12676 5364
rect 12624 5321 12633 5355
rect 12633 5321 12667 5355
rect 12667 5321 12676 5355
rect 12624 5312 12676 5321
rect 13084 5312 13136 5364
rect 15292 5312 15344 5364
rect 16212 5312 16264 5364
rect 17500 5312 17552 5364
rect 18696 5312 18748 5364
rect 22744 5312 22796 5364
rect 24952 5312 25004 5364
rect 26700 5312 26752 5364
rect 28264 5312 28316 5364
rect 28356 5312 28408 5364
rect 31024 5355 31076 5364
rect 31024 5321 31033 5355
rect 31033 5321 31067 5355
rect 31067 5321 31076 5355
rect 31024 5312 31076 5321
rect 31300 5312 31352 5364
rect 33876 5312 33928 5364
rect 35900 5355 35952 5364
rect 35900 5321 35909 5355
rect 35909 5321 35943 5355
rect 35943 5321 35952 5355
rect 35900 5312 35952 5321
rect 2596 5108 2648 5160
rect 2872 5108 2924 5160
rect 3976 5108 4028 5160
rect 2504 5083 2556 5092
rect 2504 5049 2513 5083
rect 2513 5049 2547 5083
rect 2547 5049 2556 5083
rect 2504 5040 2556 5049
rect 4160 5083 4212 5092
rect 4160 5049 4169 5083
rect 4169 5049 4203 5083
rect 4203 5049 4212 5083
rect 4160 5040 4212 5049
rect 6736 5108 6788 5160
rect 9404 5108 9456 5160
rect 10600 5176 10652 5228
rect 11980 5176 12032 5228
rect 11152 5151 11204 5160
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 11520 5151 11572 5160
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 8116 5040 8168 5092
rect 19064 5244 19116 5296
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 15384 5176 15436 5185
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 19248 5219 19300 5228
rect 19248 5185 19257 5219
rect 19257 5185 19291 5219
rect 19291 5185 19300 5219
rect 19248 5176 19300 5185
rect 19616 5176 19668 5228
rect 21456 5244 21508 5296
rect 21640 5287 21692 5296
rect 21640 5253 21649 5287
rect 21649 5253 21683 5287
rect 21683 5253 21692 5287
rect 21640 5244 21692 5253
rect 26884 5244 26936 5296
rect 34704 5244 34756 5296
rect 36636 5244 36688 5296
rect 23480 5176 23532 5228
rect 24860 5176 24912 5228
rect 26056 5219 26108 5228
rect 26056 5185 26065 5219
rect 26065 5185 26099 5219
rect 26099 5185 26108 5219
rect 26056 5176 26108 5185
rect 26148 5176 26200 5228
rect 15200 5151 15252 5160
rect 15200 5117 15209 5151
rect 15209 5117 15243 5151
rect 15243 5117 15252 5151
rect 15200 5108 15252 5117
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 24308 5108 24360 5160
rect 9496 5015 9548 5024
rect 9496 4981 9505 5015
rect 9505 4981 9539 5015
rect 9539 4981 9548 5015
rect 9496 4972 9548 4981
rect 10784 4972 10836 5024
rect 15844 5040 15896 5092
rect 19340 5040 19392 5092
rect 19708 5040 19760 5092
rect 16948 4972 17000 5024
rect 17684 5015 17736 5024
rect 17684 4981 17693 5015
rect 17693 4981 17727 5015
rect 17727 4981 17736 5015
rect 17684 4972 17736 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 20536 4972 20588 5024
rect 24400 5040 24452 5092
rect 22284 4972 22336 5024
rect 22560 5015 22612 5024
rect 22560 4981 22569 5015
rect 22569 4981 22603 5015
rect 22603 4981 22612 5015
rect 22560 4972 22612 4981
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 27068 5176 27120 5228
rect 27252 5219 27304 5228
rect 27252 5185 27261 5219
rect 27261 5185 27295 5219
rect 27295 5185 27304 5219
rect 27252 5176 27304 5185
rect 28172 5176 28224 5228
rect 31852 5176 31904 5228
rect 32956 5176 33008 5228
rect 30840 5151 30892 5160
rect 30840 5117 30849 5151
rect 30849 5117 30883 5151
rect 30883 5117 30892 5151
rect 30840 5108 30892 5117
rect 31576 5108 31628 5160
rect 29092 5040 29144 5092
rect 30196 5040 30248 5092
rect 32496 5040 32548 5092
rect 34152 5176 34204 5228
rect 35072 5176 35124 5228
rect 35348 5219 35400 5228
rect 35348 5185 35357 5219
rect 35357 5185 35391 5219
rect 35391 5185 35400 5219
rect 35348 5176 35400 5185
rect 35992 5176 36044 5228
rect 35072 5083 35124 5092
rect 35072 5049 35081 5083
rect 35081 5049 35115 5083
rect 35115 5049 35124 5083
rect 35072 5040 35124 5049
rect 36176 5040 36228 5092
rect 36636 5083 36688 5092
rect 36636 5049 36645 5083
rect 36645 5049 36679 5083
rect 36679 5049 36688 5083
rect 36636 5040 36688 5049
rect 30472 4972 30524 5024
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 1952 4768 2004 4820
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 6092 4768 6144 4820
rect 8116 4768 8168 4820
rect 12164 4811 12216 4820
rect 2504 4700 2556 4752
rect 3976 4700 4028 4752
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 3148 4564 3200 4616
rect 8484 4632 8536 4684
rect 9220 4700 9272 4752
rect 10140 4700 10192 4752
rect 10968 4700 11020 4752
rect 12164 4777 12173 4811
rect 12173 4777 12207 4811
rect 12207 4777 12216 4811
rect 12164 4768 12216 4777
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 13084 4768 13136 4820
rect 13452 4768 13504 4820
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 14188 4768 14240 4820
rect 16948 4768 17000 4820
rect 18144 4768 18196 4820
rect 20536 4768 20588 4820
rect 21916 4811 21968 4820
rect 21916 4777 21925 4811
rect 21925 4777 21959 4811
rect 21959 4777 21968 4811
rect 21916 4768 21968 4777
rect 24308 4811 24360 4820
rect 24308 4777 24317 4811
rect 24317 4777 24351 4811
rect 24351 4777 24360 4811
rect 24308 4768 24360 4777
rect 25964 4768 26016 4820
rect 29092 4768 29144 4820
rect 32588 4811 32640 4820
rect 32588 4777 32597 4811
rect 32597 4777 32631 4811
rect 32631 4777 32640 4811
rect 32588 4768 32640 4777
rect 32956 4811 33008 4820
rect 32956 4777 32965 4811
rect 32965 4777 32999 4811
rect 32999 4777 33008 4811
rect 32956 4768 33008 4777
rect 34980 4811 35032 4820
rect 34980 4777 34989 4811
rect 34989 4777 35023 4811
rect 35023 4777 35032 4811
rect 34980 4768 35032 4777
rect 35072 4768 35124 4820
rect 36176 4768 36228 4820
rect 11980 4700 12032 4752
rect 13728 4743 13780 4752
rect 13728 4709 13737 4743
rect 13737 4709 13771 4743
rect 13771 4709 13780 4743
rect 13728 4700 13780 4709
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 7472 4564 7524 4616
rect 8024 4564 8076 4616
rect 9496 4564 9548 4616
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 11060 4564 11112 4616
rect 14648 4564 14700 4616
rect 15108 4564 15160 4616
rect 17500 4700 17552 4752
rect 17684 4700 17736 4752
rect 19708 4700 19760 4752
rect 20812 4700 20864 4752
rect 21640 4743 21692 4752
rect 21640 4709 21649 4743
rect 21649 4709 21683 4743
rect 21683 4709 21692 4743
rect 21640 4700 21692 4709
rect 24032 4743 24084 4752
rect 24032 4709 24041 4743
rect 24041 4709 24075 4743
rect 24075 4709 24084 4743
rect 24032 4700 24084 4709
rect 26700 4743 26752 4752
rect 26700 4709 26709 4743
rect 26709 4709 26743 4743
rect 26743 4709 26752 4743
rect 26700 4700 26752 4709
rect 28264 4743 28316 4752
rect 28264 4709 28273 4743
rect 28273 4709 28307 4743
rect 28307 4709 28316 4743
rect 28264 4700 28316 4709
rect 34152 4700 34204 4752
rect 34888 4700 34940 4752
rect 18512 4632 18564 4684
rect 23388 4675 23440 4684
rect 23388 4641 23397 4675
rect 23397 4641 23431 4675
rect 23431 4641 23440 4675
rect 23388 4632 23440 4641
rect 23664 4632 23716 4684
rect 16672 4564 16724 4616
rect 21272 4564 21324 4616
rect 22560 4564 22612 4616
rect 24768 4632 24820 4684
rect 30380 4632 30432 4684
rect 31024 4675 31076 4684
rect 31024 4641 31033 4675
rect 31033 4641 31067 4675
rect 31067 4641 31076 4675
rect 31024 4632 31076 4641
rect 35256 4632 35308 4684
rect 35440 4743 35492 4752
rect 35440 4709 35449 4743
rect 35449 4709 35483 4743
rect 35483 4709 35492 4743
rect 35440 4700 35492 4709
rect 35808 4632 35860 4684
rect 25136 4564 25188 4616
rect 25964 4564 26016 4616
rect 27252 4564 27304 4616
rect 28172 4607 28224 4616
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 32128 4607 32180 4616
rect 2872 4496 2924 4548
rect 4252 4496 4304 4548
rect 4712 4539 4764 4548
rect 4712 4505 4721 4539
rect 4721 4505 4755 4539
rect 4755 4505 4764 4539
rect 4712 4496 4764 4505
rect 11152 4496 11204 4548
rect 17960 4496 18012 4548
rect 23020 4496 23072 4548
rect 23296 4496 23348 4548
rect 27160 4539 27212 4548
rect 27160 4505 27169 4539
rect 27169 4505 27203 4539
rect 27203 4505 27212 4539
rect 32128 4573 32137 4607
rect 32137 4573 32171 4607
rect 32171 4573 32180 4607
rect 32128 4564 32180 4573
rect 33968 4564 34020 4616
rect 35164 4607 35216 4616
rect 35164 4573 35173 4607
rect 35173 4573 35207 4607
rect 35207 4573 35216 4607
rect 35164 4564 35216 4573
rect 27160 4496 27212 4505
rect 28816 4496 28868 4548
rect 2780 4428 2832 4480
rect 9036 4471 9088 4480
rect 9036 4437 9045 4471
rect 9045 4437 9079 4471
rect 9079 4437 9088 4471
rect 9036 4428 9088 4437
rect 9404 4471 9456 4480
rect 9404 4437 9413 4471
rect 9413 4437 9447 4471
rect 9447 4437 9456 4471
rect 9404 4428 9456 4437
rect 10968 4428 11020 4480
rect 12992 4428 13044 4480
rect 13820 4428 13872 4480
rect 15200 4428 15252 4480
rect 16488 4428 16540 4480
rect 16948 4428 17000 4480
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17316 4428 17368 4437
rect 18328 4428 18380 4480
rect 19156 4428 19208 4480
rect 31484 4471 31536 4480
rect 31484 4437 31493 4471
rect 31493 4437 31527 4471
rect 31527 4437 31536 4471
rect 31484 4428 31536 4437
rect 34612 4428 34664 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 2504 4267 2556 4276
rect 2504 4233 2513 4267
rect 2513 4233 2547 4267
rect 2547 4233 2556 4267
rect 2504 4224 2556 4233
rect 1492 4063 1544 4072
rect 1492 4029 1501 4063
rect 1501 4029 1535 4063
rect 1535 4029 1544 4063
rect 2320 4156 2372 4208
rect 2872 4156 2924 4208
rect 4712 4224 4764 4276
rect 3976 4199 4028 4208
rect 3976 4165 3985 4199
rect 3985 4165 4019 4199
rect 4019 4165 4028 4199
rect 3976 4156 4028 4165
rect 5632 4156 5684 4208
rect 5816 4156 5868 4208
rect 6736 4224 6788 4276
rect 6828 4224 6880 4276
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 11520 4224 11572 4276
rect 15752 4224 15804 4276
rect 16120 4224 16172 4276
rect 17132 4224 17184 4276
rect 18144 4224 18196 4276
rect 19708 4224 19760 4276
rect 20812 4224 20864 4276
rect 21272 4267 21324 4276
rect 21272 4233 21281 4267
rect 21281 4233 21315 4267
rect 21315 4233 21324 4267
rect 21272 4224 21324 4233
rect 23388 4224 23440 4276
rect 23664 4224 23716 4276
rect 24400 4224 24452 4276
rect 6552 4156 6604 4208
rect 9864 4156 9916 4208
rect 10232 4156 10284 4208
rect 11336 4199 11388 4208
rect 11336 4165 11345 4199
rect 11345 4165 11379 4199
rect 11379 4165 11388 4199
rect 11336 4156 11388 4165
rect 11980 4156 12032 4208
rect 12716 4199 12768 4208
rect 12716 4165 12725 4199
rect 12725 4165 12759 4199
rect 12759 4165 12768 4199
rect 12716 4156 12768 4165
rect 13820 4156 13872 4208
rect 16488 4199 16540 4208
rect 16488 4165 16512 4199
rect 16512 4165 16540 4199
rect 16488 4156 16540 4165
rect 17868 4156 17920 4208
rect 18328 4199 18380 4208
rect 18328 4165 18337 4199
rect 18337 4165 18371 4199
rect 18371 4165 18380 4199
rect 18328 4156 18380 4165
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 3884 4088 3936 4140
rect 5448 4088 5500 4140
rect 7472 4088 7524 4140
rect 13084 4088 13136 4140
rect 16304 4088 16356 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 1492 4020 1544 4029
rect 6092 4020 6144 4072
rect 9680 4020 9732 4072
rect 10968 4020 11020 4072
rect 2780 3995 2832 4004
rect 2780 3961 2789 3995
rect 2789 3961 2823 3995
rect 2823 3961 2832 3995
rect 2780 3952 2832 3961
rect 2228 3884 2280 3936
rect 4896 3995 4948 4004
rect 4896 3961 4905 3995
rect 4905 3961 4939 3995
rect 4939 3961 4948 3995
rect 4896 3952 4948 3961
rect 5264 3927 5316 3936
rect 5264 3893 5273 3927
rect 5273 3893 5307 3927
rect 5307 3893 5316 3927
rect 5264 3884 5316 3893
rect 7932 3952 7984 4004
rect 8116 3952 8168 4004
rect 11060 3952 11112 4004
rect 8300 3884 8352 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 10508 3884 10560 3936
rect 13636 4020 13688 4072
rect 13912 4020 13964 4072
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 15200 4020 15252 4072
rect 15660 4020 15712 4072
rect 11796 3952 11848 4004
rect 14648 3952 14700 4004
rect 14924 3995 14976 4004
rect 14924 3961 14933 3995
rect 14933 3961 14967 3995
rect 14967 3961 14976 3995
rect 14924 3952 14976 3961
rect 15292 3952 15344 4004
rect 18144 4020 18196 4072
rect 21364 4156 21416 4208
rect 22284 4156 22336 4208
rect 23204 4156 23256 4208
rect 24676 4156 24728 4208
rect 21088 4088 21140 4140
rect 19892 4020 19944 4072
rect 20628 4020 20680 4072
rect 21732 4063 21784 4072
rect 21732 4029 21741 4063
rect 21741 4029 21775 4063
rect 21775 4029 21784 4063
rect 21732 4020 21784 4029
rect 22284 4063 22336 4072
rect 22284 4029 22293 4063
rect 22293 4029 22327 4063
rect 22327 4029 22336 4063
rect 22284 4020 22336 4029
rect 16580 3952 16632 4004
rect 17500 3952 17552 4004
rect 12992 3884 13044 3936
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 19708 3884 19760 3936
rect 26240 4224 26292 4276
rect 26700 4224 26752 4276
rect 28264 4224 28316 4276
rect 31024 4224 31076 4276
rect 34612 4267 34664 4276
rect 24860 4156 24912 4208
rect 30380 4156 30432 4208
rect 24952 4063 25004 4072
rect 24952 4029 24961 4063
rect 24961 4029 24995 4063
rect 24995 4029 25004 4063
rect 24952 4020 25004 4029
rect 28908 4088 28960 4140
rect 29552 4088 29604 4140
rect 29368 4063 29420 4072
rect 29368 4029 29377 4063
rect 29377 4029 29411 4063
rect 29411 4029 29420 4063
rect 29368 4020 29420 4029
rect 31208 4156 31260 4208
rect 31392 4088 31444 4140
rect 32588 4063 32640 4072
rect 28356 3952 28408 4004
rect 32588 4029 32597 4063
rect 32597 4029 32631 4063
rect 32631 4029 32640 4063
rect 32588 4020 32640 4029
rect 30104 3995 30156 4004
rect 30104 3961 30113 3995
rect 30113 3961 30147 3995
rect 30147 3961 30156 3995
rect 30104 3952 30156 3961
rect 31484 3952 31536 4004
rect 33600 4156 33652 4208
rect 34152 4156 34204 4208
rect 34612 4233 34621 4267
rect 34621 4233 34655 4267
rect 34655 4233 34664 4267
rect 34612 4224 34664 4233
rect 34888 4224 34940 4276
rect 35440 4224 35492 4276
rect 35992 4224 36044 4276
rect 36728 4224 36780 4276
rect 35348 4156 35400 4208
rect 36452 4063 36504 4072
rect 36452 4029 36461 4063
rect 36461 4029 36495 4063
rect 36495 4029 36504 4063
rect 37004 4063 37056 4072
rect 36452 4020 36504 4029
rect 37004 4029 37013 4063
rect 37013 4029 37047 4063
rect 37047 4029 37056 4063
rect 37004 4020 37056 4029
rect 37372 4020 37424 4072
rect 33324 3995 33376 4004
rect 22008 3927 22060 3936
rect 22008 3893 22017 3927
rect 22017 3893 22051 3927
rect 22051 3893 22060 3927
rect 22008 3884 22060 3893
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 26148 3927 26200 3936
rect 26148 3893 26157 3927
rect 26157 3893 26191 3927
rect 26191 3893 26200 3927
rect 26148 3884 26200 3893
rect 27344 3884 27396 3936
rect 28172 3884 28224 3936
rect 29000 3927 29052 3936
rect 29000 3893 29009 3927
rect 29009 3893 29043 3927
rect 29043 3893 29052 3927
rect 29000 3884 29052 3893
rect 29092 3884 29144 3936
rect 33324 3961 33333 3995
rect 33333 3961 33367 3995
rect 33367 3961 33376 3995
rect 33324 3952 33376 3961
rect 33140 3884 33192 3936
rect 33968 3927 34020 3936
rect 33968 3893 33977 3927
rect 33977 3893 34011 3927
rect 34011 3893 34020 3927
rect 33968 3884 34020 3893
rect 34612 3884 34664 3936
rect 35440 3952 35492 4004
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 2780 3723 2832 3732
rect 2780 3689 2789 3723
rect 2789 3689 2823 3723
rect 2823 3689 2832 3723
rect 2780 3680 2832 3689
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 1676 3612 1728 3664
rect 2504 3612 2556 3664
rect 4252 3680 4304 3732
rect 6736 3680 6788 3732
rect 8024 3680 8076 3732
rect 8300 3680 8352 3732
rect 9220 3680 9272 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 11060 3723 11112 3732
rect 11060 3689 11069 3723
rect 11069 3689 11103 3723
rect 11103 3689 11112 3723
rect 11060 3680 11112 3689
rect 11888 3680 11940 3732
rect 13636 3680 13688 3732
rect 14004 3680 14056 3732
rect 18328 3680 18380 3732
rect 18972 3723 19024 3732
rect 18972 3689 18981 3723
rect 18981 3689 19015 3723
rect 19015 3689 19024 3723
rect 18972 3680 19024 3689
rect 19524 3680 19576 3732
rect 20812 3680 20864 3732
rect 3700 3544 3752 3596
rect 4620 3587 4672 3596
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 6368 3612 6420 3664
rect 6828 3612 6880 3664
rect 8116 3612 8168 3664
rect 8760 3612 8812 3664
rect 12992 3612 13044 3664
rect 13084 3612 13136 3664
rect 13820 3655 13872 3664
rect 13820 3621 13829 3655
rect 13829 3621 13863 3655
rect 13863 3621 13872 3655
rect 13820 3612 13872 3621
rect 6276 3544 6328 3596
rect 6736 3544 6788 3596
rect 9588 3544 9640 3596
rect 11060 3587 11112 3596
rect 11060 3553 11069 3587
rect 11069 3553 11103 3587
rect 11103 3553 11112 3587
rect 11060 3544 11112 3553
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 11796 3587 11848 3596
rect 11796 3553 11805 3587
rect 11805 3553 11839 3587
rect 11839 3553 11848 3587
rect 11796 3544 11848 3553
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 5816 3476 5868 3528
rect 9036 3476 9088 3528
rect 10876 3476 10928 3528
rect 13912 3544 13964 3596
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 18052 3612 18104 3664
rect 18236 3655 18288 3664
rect 18236 3621 18245 3655
rect 18245 3621 18279 3655
rect 18279 3621 18288 3655
rect 18236 3612 18288 3621
rect 19892 3655 19944 3664
rect 19892 3621 19901 3655
rect 19901 3621 19935 3655
rect 19935 3621 19944 3655
rect 19892 3612 19944 3621
rect 18972 3544 19024 3596
rect 19616 3587 19668 3596
rect 19616 3553 19625 3587
rect 19625 3553 19659 3587
rect 19659 3553 19668 3587
rect 19616 3544 19668 3553
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 14648 3476 14700 3528
rect 16672 3476 16724 3528
rect 17132 3476 17184 3528
rect 22008 3680 22060 3732
rect 22744 3723 22796 3732
rect 22744 3689 22753 3723
rect 22753 3689 22787 3723
rect 22787 3689 22796 3723
rect 22744 3680 22796 3689
rect 23480 3680 23532 3732
rect 25136 3723 25188 3732
rect 23664 3612 23716 3664
rect 24216 3655 24268 3664
rect 24216 3621 24225 3655
rect 24225 3621 24259 3655
rect 24259 3621 24268 3655
rect 24216 3612 24268 3621
rect 25136 3689 25145 3723
rect 25145 3689 25179 3723
rect 25179 3689 25188 3723
rect 25136 3680 25188 3689
rect 25964 3723 26016 3732
rect 25964 3689 25973 3723
rect 25973 3689 26007 3723
rect 26007 3689 26016 3723
rect 25964 3680 26016 3689
rect 26240 3723 26292 3732
rect 26240 3689 26249 3723
rect 26249 3689 26283 3723
rect 26283 3689 26292 3723
rect 26240 3680 26292 3689
rect 28080 3723 28132 3732
rect 28080 3689 28089 3723
rect 28089 3689 28123 3723
rect 28123 3689 28132 3723
rect 28080 3680 28132 3689
rect 29092 3680 29144 3732
rect 30104 3723 30156 3732
rect 30104 3689 30113 3723
rect 30113 3689 30147 3723
rect 30147 3689 30156 3723
rect 30104 3680 30156 3689
rect 26056 3612 26108 3664
rect 26884 3612 26936 3664
rect 27344 3655 27396 3664
rect 27344 3621 27353 3655
rect 27353 3621 27387 3655
rect 27387 3621 27396 3655
rect 27344 3612 27396 3621
rect 28356 3612 28408 3664
rect 31484 3680 31536 3732
rect 10140 3408 10192 3460
rect 12624 3408 12676 3460
rect 16488 3408 16540 3460
rect 17868 3408 17920 3460
rect 21272 3476 21324 3528
rect 24400 3476 24452 3528
rect 23112 3408 23164 3460
rect 24124 3408 24176 3460
rect 26332 3476 26384 3528
rect 26792 3476 26844 3528
rect 28172 3519 28224 3528
rect 28172 3485 28181 3519
rect 28181 3485 28215 3519
rect 28215 3485 28224 3519
rect 28172 3476 28224 3485
rect 25412 3408 25464 3460
rect 29460 3408 29512 3460
rect 30196 3408 30248 3460
rect 31208 3612 31260 3664
rect 30380 3544 30432 3596
rect 31852 3544 31904 3596
rect 33600 3612 33652 3664
rect 36268 3612 36320 3664
rect 33324 3544 33376 3596
rect 35164 3519 35216 3528
rect 35164 3485 35173 3519
rect 35173 3485 35207 3519
rect 35207 3485 35216 3519
rect 35164 3476 35216 3485
rect 35900 3476 35952 3528
rect 35624 3408 35676 3460
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 5080 3340 5132 3392
rect 5448 3340 5500 3392
rect 8024 3340 8076 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 13820 3340 13872 3392
rect 14740 3340 14792 3392
rect 15108 3340 15160 3392
rect 15568 3383 15620 3392
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 16304 3340 16356 3392
rect 18052 3340 18104 3392
rect 18328 3340 18380 3392
rect 21732 3383 21784 3392
rect 21732 3349 21741 3383
rect 21741 3349 21775 3383
rect 21775 3349 21784 3383
rect 21732 3340 21784 3349
rect 24400 3340 24452 3392
rect 24952 3340 25004 3392
rect 27436 3340 27488 3392
rect 29368 3383 29420 3392
rect 29368 3349 29377 3383
rect 29377 3349 29411 3383
rect 29411 3349 29420 3383
rect 29368 3340 29420 3349
rect 31484 3383 31536 3392
rect 31484 3349 31493 3383
rect 31493 3349 31527 3383
rect 31527 3349 31536 3383
rect 31484 3340 31536 3349
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 4620 3136 4672 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 8116 3179 8168 3188
rect 6276 3136 6328 3145
rect 1768 3000 1820 3052
rect 3240 3068 3292 3120
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 5724 3000 5776 3052
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2504 2864 2556 2916
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5448 2975 5500 2984
rect 5264 2932 5316 2941
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 9496 3136 9548 3188
rect 9956 3136 10008 3188
rect 10508 3179 10560 3188
rect 10508 3145 10517 3179
rect 10517 3145 10551 3179
rect 10551 3145 10560 3179
rect 10508 3136 10560 3145
rect 12716 3136 12768 3188
rect 13176 3136 13228 3188
rect 16120 3136 16172 3188
rect 8944 3068 8996 3120
rect 13268 3068 13320 3120
rect 13728 3068 13780 3120
rect 15200 3068 15252 3120
rect 16488 3068 16540 3120
rect 17132 3068 17184 3120
rect 20812 3136 20864 3188
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 21824 3179 21876 3188
rect 21824 3145 21833 3179
rect 21833 3145 21867 3179
rect 21867 3145 21876 3179
rect 21824 3136 21876 3145
rect 22744 3136 22796 3188
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 24216 3179 24268 3188
rect 23480 3136 23532 3145
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 26056 3179 26108 3188
rect 26056 3145 26065 3179
rect 26065 3145 26099 3179
rect 26099 3145 26108 3179
rect 26056 3136 26108 3145
rect 28356 3136 28408 3188
rect 30196 3136 30248 3188
rect 30288 3136 30340 3188
rect 31852 3179 31904 3188
rect 27160 3111 27212 3120
rect 27160 3077 27169 3111
rect 27169 3077 27203 3111
rect 27203 3077 27212 3111
rect 27160 3068 27212 3077
rect 11612 3000 11664 3052
rect 16028 3043 16080 3052
rect 7932 2932 7984 2984
rect 8852 2932 8904 2984
rect 10508 2932 10560 2984
rect 12532 2975 12584 2984
rect 12532 2941 12541 2975
rect 12541 2941 12575 2975
rect 12575 2941 12584 2975
rect 12532 2932 12584 2941
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 16028 3009 16037 3043
rect 16037 3009 16071 3043
rect 16071 3009 16080 3043
rect 16028 3000 16080 3009
rect 16764 3000 16816 3052
rect 19616 3000 19668 3052
rect 14004 2975 14056 2984
rect 12716 2932 12768 2941
rect 14004 2941 14013 2975
rect 14013 2941 14047 2975
rect 14047 2941 14056 2975
rect 14004 2932 14056 2941
rect 14188 2932 14240 2984
rect 14740 2932 14792 2984
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 18052 2975 18104 2984
rect 9496 2864 9548 2916
rect 9680 2864 9732 2916
rect 4712 2839 4764 2848
rect 2044 2796 2096 2805
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 6276 2796 6328 2848
rect 8024 2796 8076 2848
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 30012 3043 30064 3052
rect 30012 3009 30021 3043
rect 30021 3009 30055 3043
rect 30055 3009 30064 3043
rect 30012 3000 30064 3009
rect 17776 2864 17828 2916
rect 19616 2864 19668 2916
rect 19800 2864 19852 2916
rect 21824 2864 21876 2916
rect 23388 2932 23440 2984
rect 24768 2975 24820 2984
rect 24768 2941 24777 2975
rect 24777 2941 24811 2975
rect 24811 2941 24820 2975
rect 24768 2932 24820 2941
rect 28080 2932 28132 2984
rect 31852 3145 31861 3179
rect 31861 3145 31895 3179
rect 31895 3145 31904 3179
rect 31852 3136 31904 3145
rect 32312 3179 32364 3188
rect 32312 3145 32321 3179
rect 32321 3145 32355 3179
rect 32355 3145 32364 3179
rect 32312 3136 32364 3145
rect 33324 3136 33376 3188
rect 34704 3179 34756 3188
rect 34704 3145 34713 3179
rect 34713 3145 34747 3179
rect 34747 3145 34756 3179
rect 34704 3136 34756 3145
rect 35900 3179 35952 3188
rect 35900 3145 35909 3179
rect 35909 3145 35943 3179
rect 35943 3145 35952 3179
rect 35900 3136 35952 3145
rect 36268 3179 36320 3188
rect 36268 3145 36277 3179
rect 36277 3145 36311 3179
rect 36311 3145 36320 3179
rect 36268 3136 36320 3145
rect 33600 3068 33652 3120
rect 33784 3068 33836 3120
rect 31576 3043 31628 3052
rect 31576 3009 31585 3043
rect 31585 3009 31619 3043
rect 31619 3009 31628 3043
rect 31576 3000 31628 3009
rect 33140 3043 33192 3052
rect 33140 3009 33149 3043
rect 33149 3009 33183 3043
rect 33183 3009 33192 3043
rect 34980 3043 35032 3052
rect 33140 3000 33192 3009
rect 34980 3009 34989 3043
rect 34989 3009 35023 3043
rect 35023 3009 35032 3043
rect 34980 3000 35032 3009
rect 35440 3000 35492 3052
rect 35808 3000 35860 3052
rect 31208 2932 31260 2984
rect 32312 2932 32364 2984
rect 32864 2975 32916 2984
rect 32864 2941 32873 2975
rect 32873 2941 32907 2975
rect 32907 2941 32916 2975
rect 32864 2932 32916 2941
rect 37004 2932 37056 2984
rect 24400 2864 24452 2916
rect 13728 2796 13780 2848
rect 14096 2796 14148 2848
rect 14648 2796 14700 2848
rect 15568 2796 15620 2848
rect 18328 2796 18380 2848
rect 19524 2796 19576 2848
rect 29092 2864 29144 2916
rect 28172 2796 28224 2848
rect 29460 2907 29512 2916
rect 29460 2873 29469 2907
rect 29469 2873 29503 2907
rect 29503 2873 29512 2907
rect 29460 2864 29512 2873
rect 32128 2864 32180 2916
rect 34704 2796 34756 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 2044 2635 2096 2644
rect 2044 2601 2053 2635
rect 2053 2601 2087 2635
rect 2087 2601 2096 2635
rect 2044 2592 2096 2601
rect 2228 2567 2280 2576
rect 2228 2533 2237 2567
rect 2237 2533 2271 2567
rect 2271 2533 2280 2567
rect 2228 2524 2280 2533
rect 4712 2592 4764 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 9312 2592 9364 2644
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 12808 2592 12860 2644
rect 13268 2635 13320 2644
rect 13268 2601 13277 2635
rect 13277 2601 13311 2635
rect 13311 2601 13320 2635
rect 13268 2592 13320 2601
rect 14004 2592 14056 2644
rect 14740 2592 14792 2644
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 4804 2524 4856 2576
rect 8852 2567 8904 2576
rect 3332 2456 3384 2508
rect 5080 2456 5132 2508
rect 5448 2456 5500 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 8484 2456 8536 2508
rect 8852 2533 8861 2567
rect 8861 2533 8895 2567
rect 8895 2533 8904 2567
rect 8852 2524 8904 2533
rect 9956 2567 10008 2576
rect 9956 2533 9965 2567
rect 9965 2533 9999 2567
rect 9999 2533 10008 2567
rect 9956 2524 10008 2533
rect 11060 2524 11112 2576
rect 2228 2388 2280 2440
rect 1584 2320 1636 2372
rect 6276 2388 6328 2440
rect 9312 2388 9364 2440
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 4988 2363 5040 2372
rect 4988 2329 4997 2363
rect 4997 2329 5031 2363
rect 5031 2329 5040 2363
rect 4988 2320 5040 2329
rect 5448 2252 5500 2304
rect 9404 2320 9456 2372
rect 12532 2456 12584 2508
rect 13728 2456 13780 2508
rect 13912 2456 13964 2508
rect 15200 2456 15252 2508
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 16580 2456 16632 2465
rect 17316 2592 17368 2644
rect 17592 2635 17644 2644
rect 17592 2601 17601 2635
rect 17601 2601 17635 2635
rect 17635 2601 17644 2635
rect 17592 2592 17644 2601
rect 21364 2635 21416 2644
rect 21364 2601 21373 2635
rect 21373 2601 21407 2635
rect 21407 2601 21416 2635
rect 21364 2592 21416 2601
rect 18328 2567 18380 2576
rect 18328 2533 18337 2567
rect 18337 2533 18371 2567
rect 18371 2533 18380 2567
rect 18328 2524 18380 2533
rect 19800 2524 19852 2576
rect 17960 2456 18012 2508
rect 19156 2456 19208 2508
rect 24768 2592 24820 2644
rect 25412 2635 25464 2644
rect 25412 2601 25421 2635
rect 25421 2601 25455 2635
rect 25455 2601 25464 2635
rect 25412 2592 25464 2601
rect 26332 2635 26384 2644
rect 26332 2601 26341 2635
rect 26341 2601 26375 2635
rect 26375 2601 26384 2635
rect 26332 2592 26384 2601
rect 29460 2592 29512 2644
rect 29552 2635 29604 2644
rect 29552 2601 29561 2635
rect 29561 2601 29595 2635
rect 29595 2601 29604 2635
rect 29552 2592 29604 2601
rect 30012 2592 30064 2644
rect 24860 2524 24912 2576
rect 18144 2388 18196 2440
rect 8208 2252 8260 2304
rect 16120 2320 16172 2372
rect 17776 2320 17828 2372
rect 18972 2320 19024 2372
rect 21732 2320 21784 2372
rect 23388 2431 23440 2440
rect 23388 2397 23397 2431
rect 23397 2397 23431 2431
rect 23431 2397 23440 2431
rect 28172 2567 28224 2576
rect 27436 2499 27488 2508
rect 23388 2388 23440 2397
rect 26148 2388 26200 2440
rect 27436 2465 27445 2499
rect 27445 2465 27479 2499
rect 27479 2465 27488 2499
rect 27436 2456 27488 2465
rect 28172 2533 28181 2567
rect 28181 2533 28215 2567
rect 28215 2533 28224 2567
rect 28172 2524 28224 2533
rect 29000 2524 29052 2576
rect 28632 2456 28684 2508
rect 30472 2567 30524 2576
rect 30472 2533 30481 2567
rect 30481 2533 30515 2567
rect 30515 2533 30524 2567
rect 30472 2524 30524 2533
rect 31208 2524 31260 2576
rect 31484 2592 31536 2644
rect 34060 2635 34112 2644
rect 34060 2601 34069 2635
rect 34069 2601 34103 2635
rect 34103 2601 34112 2635
rect 34060 2592 34112 2601
rect 34980 2635 35032 2644
rect 34980 2601 34989 2635
rect 34989 2601 35023 2635
rect 35023 2601 35032 2635
rect 34980 2592 35032 2601
rect 35624 2592 35676 2644
rect 36912 2499 36964 2508
rect 36912 2465 36921 2499
rect 36921 2465 36955 2499
rect 36955 2465 36964 2499
rect 36912 2456 36964 2465
rect 31760 2388 31812 2440
rect 31208 2320 31260 2372
rect 32864 2320 32916 2372
rect 36084 2320 36136 2372
rect 12256 2252 12308 2304
rect 12624 2252 12676 2304
rect 12900 2295 12952 2304
rect 12900 2261 12909 2295
rect 12909 2261 12943 2295
rect 12943 2261 12952 2295
rect 12900 2252 12952 2261
rect 12992 2252 13044 2304
rect 14648 2252 14700 2304
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 15660 2252 15712 2304
rect 26516 2252 26568 2304
rect 27528 2252 27580 2304
rect 35992 2252 36044 2304
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
<< metal2 >>
rect 6642 15586 6698 16000
rect 19982 15586 20038 16000
rect 33322 15586 33378 16000
rect 6288 15558 6698 15586
rect 938 15056 994 15065
rect 938 14991 994 15000
rect 110 13800 166 13809
rect 110 13735 166 13744
rect 124 12986 152 13735
rect 112 12980 164 12986
rect 112 12922 164 12928
rect 112 12164 164 12170
rect 112 12106 164 12112
rect 20 11824 72 11830
rect 20 11766 72 11772
rect 32 10305 60 11766
rect 124 11121 152 12106
rect 110 11112 166 11121
rect 110 11047 166 11056
rect 952 10810 980 14991
rect 1030 14240 1086 14249
rect 1030 14175 1086 14184
rect 1044 12442 1072 14175
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 1032 12436 1084 12442
rect 1032 12378 1084 12384
rect 1490 12336 1546 12345
rect 1400 12300 1452 12306
rect 1490 12271 1546 12280
rect 1400 12242 1452 12248
rect 1412 11762 1440 12242
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 940 10804 992 10810
rect 940 10746 992 10752
rect 18 10296 74 10305
rect 18 10231 74 10240
rect 112 6656 164 6662
rect 112 6598 164 6604
rect 124 2281 152 6598
rect 1504 5370 1532 12271
rect 1596 8498 1624 12582
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2148 11694 2176 12038
rect 2332 11694 2360 12038
rect 2516 11898 2544 12242
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 11014 1808 11154
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 10130 1808 10950
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1688 9518 1716 10066
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9178 1716 9454
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 8090 1624 8298
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1688 8022 1716 8978
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1688 7410 1716 7958
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 110 2272 166 2281
rect 110 2207 166 2216
rect 1504 1057 1532 4014
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1596 2378 1624 3470
rect 1688 3194 1716 3606
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1780 3058 1808 8774
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 7002 1900 8434
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1964 5778 1992 9998
rect 2056 6866 2084 11494
rect 2148 10674 2176 11630
rect 2332 11218 2360 11630
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 2148 7002 2176 9386
rect 2240 7954 2268 11086
rect 2332 10062 2360 11154
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2424 9908 2452 10066
rect 2516 9926 2544 10542
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2332 9880 2452 9908
rect 2504 9920 2556 9926
rect 2332 9217 2360 9880
rect 2504 9862 2556 9868
rect 2516 9518 2544 9862
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2318 9208 2374 9217
rect 2318 9143 2374 9152
rect 2332 9110 2360 9143
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2424 8634 2452 9454
rect 2516 9178 2544 9454
rect 2700 9382 2728 10066
rect 2688 9376 2740 9382
rect 2686 9344 2688 9353
rect 2740 9344 2742 9353
rect 2686 9279 2742 9288
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2240 7478 2268 7890
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2228 7200 2280 7206
rect 2332 7188 2360 7958
rect 2280 7160 2360 7188
rect 2228 7142 2280 7148
rect 2240 7002 2268 7142
rect 2318 7032 2374 7041
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2228 6996 2280 7002
rect 2318 6967 2374 6976
rect 2228 6938 2280 6944
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 6458 2084 6802
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2148 6322 2176 6938
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2240 6186 2268 6938
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2240 5846 2268 6122
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1964 4826 1992 5714
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2332 4214 2360 6967
rect 2700 6066 2728 9279
rect 2608 6038 2728 6066
rect 2608 5166 2636 6038
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2516 4758 2544 5034
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2516 4282 2544 4694
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2650 2084 2790
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2240 2582 2268 3878
rect 2516 3670 2544 4218
rect 2700 4146 2728 5850
rect 2792 5710 2820 10406
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 2962 10024 3018 10033
rect 2962 9959 3018 9968
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2884 8294 2912 9046
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 8090 2912 8230
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2884 7002 2912 8026
rect 2976 7993 3004 9959
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3068 8362 3096 8842
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2962 7984 3018 7993
rect 2962 7919 3018 7928
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 3068 6934 3096 8298
rect 3160 7342 3188 10134
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2976 5370 3004 6054
rect 3252 5914 3280 9862
rect 3344 9625 3372 10542
rect 3528 10266 3556 10950
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3330 9616 3386 9625
rect 3528 9586 3556 10202
rect 3330 9551 3386 9560
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3436 9178 3464 9386
rect 3424 9172 3476 9178
rect 3344 9132 3424 9160
rect 3344 7546 3372 9132
rect 3424 9114 3476 9120
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 8090 3464 8230
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3528 6662 3556 9114
rect 3620 8974 3648 11018
rect 3712 9586 3740 11766
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3804 9518 3832 12582
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3896 10470 3924 11154
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 10169 3924 10406
rect 3882 10160 3938 10169
rect 3882 10095 3938 10104
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3896 9722 3924 9998
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3988 9654 4016 10474
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3712 9110 3740 9386
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 8090 3648 8910
rect 3712 8566 3740 9046
rect 3896 8888 3924 9522
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3804 8860 3924 8888
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3804 7970 3832 8860
rect 3882 8800 3938 8809
rect 3882 8735 3938 8744
rect 3620 7942 3832 7970
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3238 5808 3294 5817
rect 3238 5743 3294 5752
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2884 4554 2912 5102
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2792 4010 2820 4422
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2792 3738 2820 3946
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 2922 2544 3334
rect 2884 3058 2912 4150
rect 3160 3738 3188 4558
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3252 3126 3280 5743
rect 3620 3641 3648 7942
rect 3896 7478 3924 8735
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3988 7206 4016 9318
rect 4080 7410 4108 11562
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 4172 7041 4200 9454
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4264 8634 4292 9046
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 8294 4292 8570
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4264 7546 4292 7958
rect 4356 7886 4384 12038
rect 4632 11558 4660 12106
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4620 11552 4672 11558
rect 4526 11520 4582 11529
rect 4620 11494 4672 11500
rect 4526 11455 4582 11464
rect 4540 10810 4568 11455
rect 4632 11132 4660 11494
rect 4724 11286 4752 11630
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 4632 11104 4752 11132
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4448 8838 4476 10134
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8566 4476 8774
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4158 7032 4214 7041
rect 4356 7002 4384 7822
rect 4158 6967 4214 6976
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5234 3832 6054
rect 4172 5846 4200 6122
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3804 4826 3832 5170
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3988 4758 4016 5102
rect 4172 5098 4200 5782
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3988 4214 4016 4694
rect 4540 4593 4568 10406
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 8906 4660 9862
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4724 7936 4752 11104
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4816 8974 4844 10950
rect 4908 9178 4936 11630
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 4816 8634 4844 8910
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5000 8294 5028 8910
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4896 7948 4948 7954
rect 4724 7908 4896 7936
rect 4896 7890 4948 7896
rect 4712 6928 4764 6934
rect 4632 6888 4712 6916
rect 4632 6390 4660 6888
rect 4712 6870 4764 6876
rect 4908 6458 4936 7890
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4632 6118 4660 6326
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5778 4660 6054
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4526 4584 4582 4593
rect 4252 4548 4304 4554
rect 4526 4519 4582 4528
rect 4712 4548 4764 4554
rect 4252 4490 4304 4496
rect 4712 4490 4764 4496
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 3738 3924 4082
rect 4264 3738 4292 4490
rect 4724 4282 4752 4490
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4908 4010 4936 5170
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 3606 3632 3662 3641
rect 3606 3567 3662 3576
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 3712 3194 3740 3538
rect 4632 3194 4660 3538
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4724 2650 4752 2790
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 2228 2576 2280 2582
rect 2228 2518 2280 2524
rect 4804 2576 4856 2582
rect 4908 2564 4936 3946
rect 4856 2536 4936 2564
rect 4804 2518 4856 2524
rect 2240 2446 2268 2518
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1490 1048 1546 1057
rect 1490 983 1546 992
rect 1122 96 1178 480
rect 3344 82 3372 2450
rect 5000 2378 5028 8230
rect 5092 3398 5120 9454
rect 5184 6304 5212 12582
rect 5368 12374 5396 12650
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5460 11898 5488 12582
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5460 11801 5488 11834
rect 5446 11792 5502 11801
rect 5446 11727 5502 11736
rect 5552 11694 5580 11834
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5276 10810 5304 11154
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5276 10713 5304 10746
rect 5262 10704 5318 10713
rect 5262 10639 5318 10648
rect 5276 10606 5304 10639
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8498 5304 8774
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5276 8022 5304 8434
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5264 7744 5316 7750
rect 5368 7732 5396 8298
rect 5316 7704 5396 7732
rect 5264 7686 5316 7692
rect 5276 7546 5304 7686
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 7002 5396 7210
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5264 6316 5316 6322
rect 5184 6276 5264 6304
rect 5264 6258 5316 6264
rect 5276 5846 5304 6258
rect 5368 6186 5396 6938
rect 5460 6798 5488 11562
rect 6196 11558 6224 12242
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6090 11248 6146 11257
rect 6090 11183 6092 11192
rect 6144 11183 6146 11192
rect 6092 11154 6144 11160
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5644 9586 5672 10542
rect 6104 10470 6132 11154
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9654 6040 10066
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5538 9208 5594 9217
rect 5538 9143 5540 9152
rect 5592 9143 5594 9152
rect 5540 9114 5592 9120
rect 5552 8378 5580 9114
rect 5644 8498 5672 9522
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5920 9042 5948 9454
rect 6012 9382 6040 9590
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5552 8350 5672 8378
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5368 5914 5396 6122
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5840 5316 5846
rect 5460 5794 5488 6734
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5264 5782 5316 5788
rect 5368 5778 5488 5794
rect 5356 5772 5488 5778
rect 5408 5766 5488 5772
rect 5356 5714 5408 5720
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5370 5488 5646
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5552 4154 5580 6122
rect 5644 4214 5672 8350
rect 5736 8294 5764 8978
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5460 4146 5580 4154
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5448 4140 5580 4146
rect 5500 4126 5580 4140
rect 5448 4082 5500 4088
rect 5736 4049 5764 8230
rect 5814 8120 5870 8129
rect 5814 8055 5870 8064
rect 5828 7818 5856 8055
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5920 7750 5948 8978
rect 6012 8537 6040 9318
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 5998 8528 6054 8537
rect 5998 8463 6054 8472
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 6866 5948 7210
rect 6012 7002 6040 7346
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5920 5642 5948 6802
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5722 4040 5778 4049
rect 5722 3975 5778 3984
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5092 2514 5120 2994
rect 5276 2990 5304 3878
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3097 5488 3334
rect 5446 3088 5502 3097
rect 5736 3058 5764 3975
rect 5828 3534 5856 4150
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5446 3023 5502 3032
rect 5724 3052 5776 3058
rect 5460 2990 5488 3023
rect 5724 2994 5776 3000
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 5276 1873 5304 2926
rect 5460 2514 5488 2926
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5460 2310 5488 2450
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5262 1864 5318 1873
rect 5262 1799 5318 1808
rect 3422 82 3478 480
rect 3344 54 3478 82
rect 5460 82 5488 2246
rect 6012 1193 6040 6190
rect 6104 4826 6132 8910
rect 6196 7177 6224 11494
rect 6288 10810 6316 15558
rect 6642 15520 6698 15558
rect 19628 15558 20038 15586
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11218 7144 11698
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6380 7970 6408 10950
rect 6288 7942 6408 7970
rect 6182 7168 6238 7177
rect 6182 7103 6238 7112
rect 6288 6798 6316 7942
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6380 7410 6408 7754
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6458 6316 6734
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6380 6390 6408 6870
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6288 5846 6316 6054
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6288 5302 6316 5782
rect 6368 5704 6420 5710
rect 6472 5692 6500 11018
rect 7116 10674 7144 11154
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 9722 6592 9998
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6748 8090 6776 10202
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6564 6322 6592 6734
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6656 6225 6684 7686
rect 6642 6216 6698 6225
rect 6642 6151 6698 6160
rect 6420 5664 6500 5692
rect 6368 5646 6420 5652
rect 6472 5370 6500 5664
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6104 4078 6132 4762
rect 6748 4690 6776 5102
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6564 4214 6592 4626
rect 6748 4282 6776 4626
rect 6840 4282 6868 10134
rect 6932 10130 6960 10202
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6932 9654 6960 10066
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7012 9444 7064 9450
rect 6932 9404 7012 9432
rect 6932 8838 6960 9404
rect 7012 9386 7064 9392
rect 7300 8974 7328 10406
rect 7392 10169 7420 11494
rect 7378 10160 7434 10169
rect 7378 10095 7434 10104
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8090 6960 8774
rect 7300 8566 7328 8910
rect 7392 8634 7420 9046
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7300 8022 7328 8230
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7300 7274 7328 7958
rect 7378 7848 7434 7857
rect 7378 7783 7434 7792
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7300 6662 7328 7210
rect 7392 7177 7420 7783
rect 7378 7168 7434 7177
rect 7378 7103 7434 7112
rect 7484 6934 7512 12038
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 8588 10674 8616 11154
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 7576 10577 7604 10610
rect 9496 10600 9548 10606
rect 7562 10568 7618 10577
rect 9496 10542 9548 10548
rect 7562 10503 7618 10512
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 8220 9722 8248 10406
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 7576 8974 7604 9522
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8036 8090 8064 8570
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 8312 7410 8340 9318
rect 8588 8906 8616 9454
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8680 8634 8708 9522
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8668 8424 8720 8430
rect 8772 8412 8800 8774
rect 8720 8384 8800 8412
rect 8668 8366 8720 8372
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 5846 7328 6598
rect 7484 5914 7512 6870
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8036 6186 8064 6870
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 5370 7236 5714
rect 7300 5574 7328 5782
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 8036 5080 8064 5850
rect 8128 5778 8156 7142
rect 8312 7002 8340 7346
rect 8496 7274 8524 7890
rect 8680 7750 8708 8366
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8220 6322 8248 6666
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5914 8340 6122
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8312 5370 8340 5850
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8116 5092 8168 5098
rect 8036 5052 8116 5080
rect 8116 5034 8168 5040
rect 8128 4826 8156 5034
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6748 3738 6776 4218
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6288 3194 6316 3538
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6288 2446 6316 2790
rect 6380 2650 6408 3606
rect 6748 3602 6776 3674
rect 6840 3670 6868 4218
rect 7484 4146 7512 4558
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 7944 3380 7972 3946
rect 8036 3738 8064 4558
rect 8128 4010 8156 4762
rect 8496 4690 8524 6870
rect 8680 6497 8708 7686
rect 8666 6488 8722 6497
rect 8666 6423 8722 6432
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8680 4154 8708 6423
rect 8496 4126 8708 4154
rect 8864 4154 8892 10406
rect 9126 10024 9182 10033
rect 9126 9959 9182 9968
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 8090 8984 8230
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 9048 7342 9076 8842
rect 9140 7818 9168 9959
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6662 9076 7278
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8864 4126 8984 4154
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3738 8340 3878
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8024 3392 8076 3398
rect 7944 3352 8024 3380
rect 8024 3334 8076 3340
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7944 2650 7972 2926
rect 8036 2854 8064 3334
rect 8128 3194 8156 3606
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8496 2514 8524 4126
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3670 8800 3878
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8956 3126 8984 4126
rect 9048 3534 9076 4422
rect 9140 3777 9168 7210
rect 9232 6254 9260 7346
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9232 4282 9260 4694
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9218 4176 9274 4185
rect 9218 4111 9274 4120
rect 9126 3768 9182 3777
rect 9232 3738 9260 4111
rect 9126 3703 9182 3712
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8864 2582 8892 2926
rect 9324 2650 9352 10406
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9416 9382 9444 10066
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9416 8945 9444 9318
rect 9402 8936 9458 8945
rect 9402 8871 9458 8880
rect 9416 6361 9444 8871
rect 9508 7478 9536 10542
rect 9692 10470 9720 11154
rect 10428 10810 10456 12038
rect 10520 11558 10548 12242
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 10232 10464 10284 10470
rect 10520 10418 10548 11494
rect 10232 10406 10284 10412
rect 10244 10130 10272 10406
rect 10428 10390 10548 10418
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10244 9722 10272 10066
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10244 9625 10272 9658
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10428 9042 10456 10390
rect 10612 10198 10640 11630
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11256 10674 11284 11154
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 10470 11284 10610
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10612 9518 10640 10134
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8566 10456 8978
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9968 7546 9996 7754
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9402 6352 9458 6361
rect 9402 6287 9458 6296
rect 9404 5160 9456 5166
rect 9508 5148 9536 6598
rect 9600 6118 9628 6802
rect 9968 6458 9996 7482
rect 10520 7410 10548 9318
rect 10612 9178 10640 9454
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10704 9042 10732 9454
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8090 10640 8910
rect 10704 8634 10732 8978
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 8090 11008 8298
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10520 7002 10548 7346
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 11072 6866 11100 9998
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11164 7206 11192 7958
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6934 11192 7142
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10244 6254 10272 6666
rect 11072 6458 11100 6802
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9600 5273 9628 6054
rect 9784 5370 9812 6054
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9586 5264 9642 5273
rect 9586 5199 9642 5208
rect 9456 5120 9536 5148
rect 9404 5102 9456 5108
rect 9416 4486 9444 5102
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4622 9536 4966
rect 9496 4616 9548 4622
rect 9600 4593 9628 5199
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 9772 4616 9824 4622
rect 9496 4558 9548 4564
rect 9586 4584 9642 4593
rect 9772 4558 9824 4564
rect 9586 4519 9642 4528
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6932 1601 6960 2450
rect 9324 2446 9352 2586
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9416 2378 9444 4422
rect 9784 4185 9812 4558
rect 9864 4208 9916 4214
rect 9770 4176 9826 4185
rect 9864 4150 9916 4156
rect 9770 4111 9826 4120
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3194 9536 3334
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9496 2916 9548 2922
rect 9600 2904 9628 3538
rect 9692 2922 9720 4014
rect 9876 3738 9904 4150
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10152 3466 10180 4694
rect 10244 4214 10272 6190
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10428 5370 10456 5782
rect 10520 5710 10548 6122
rect 11164 6118 11192 6870
rect 11256 6769 11284 10406
rect 11532 9178 11560 11494
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11624 10130 11652 10678
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11624 9722 11652 10066
rect 11716 9926 11744 11154
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9761 11744 9862
rect 11702 9752 11758 9761
rect 11612 9716 11664 9722
rect 11808 9722 11836 12038
rect 11702 9687 11758 9696
rect 11796 9716 11848 9722
rect 11612 9658 11664 9664
rect 11796 9658 11848 9664
rect 11900 9194 11928 12582
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 12268 11626 12296 12242
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12072 11552 12124 11558
rect 12268 11529 12296 11562
rect 12440 11552 12492 11558
rect 12072 11494 12124 11500
rect 12254 11520 12310 11529
rect 12084 11393 12112 11494
rect 12440 11494 12492 11500
rect 12254 11455 12310 11464
rect 12070 11384 12126 11393
rect 12070 11319 12126 11328
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11808 9166 11928 9194
rect 11532 8634 11560 9114
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11612 8900 11664 8906
rect 11612 8842 11664 8848
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11624 7342 11652 8842
rect 11716 7886 11744 8910
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11242 6760 11298 6769
rect 11242 6695 11298 6704
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5846 11192 6054
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10520 5545 10548 5646
rect 10968 5568 11020 5574
rect 10506 5536 10562 5545
rect 10968 5510 11020 5516
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 10506 5471 10562 5480
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10612 5137 10640 5170
rect 10598 5128 10654 5137
rect 10598 5063 10654 5072
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10506 4040 10562 4049
rect 10506 3975 10562 3984
rect 10520 3942 10548 3975
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9548 2876 9628 2904
rect 9680 2916 9732 2922
rect 9496 2858 9548 2864
rect 9680 2858 9732 2864
rect 9508 2650 9536 2858
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9968 2582 9996 3130
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10152 2446 10180 3402
rect 10520 3194 10548 3878
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10520 2990 10548 3130
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 6918 1592 6974 1601
rect 6918 1527 6974 1536
rect 5998 1184 6054 1193
rect 5998 1119 6054 1128
rect 5814 82 5870 480
rect 5460 54 5870 82
rect 1122 0 1178 40
rect 3422 0 3478 54
rect 5814 0 5870 54
rect 8114 82 8170 480
rect 8220 82 8248 2246
rect 8114 54 8248 82
rect 10506 82 10562 480
rect 10796 82 10824 4966
rect 10980 4758 11008 5510
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10980 4078 11008 4422
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10980 3584 11008 4014
rect 11072 4010 11100 4558
rect 11164 4554 11192 5102
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11348 4214 11376 5510
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4282 11560 5102
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11808 4010 11836 9166
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11900 8276 11928 9046
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 8498 12020 8910
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11980 8288 12032 8294
rect 11900 8248 11980 8276
rect 11980 8230 12032 8236
rect 11992 7002 12020 8230
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11072 3738 11100 3946
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11808 3602 11836 3946
rect 11900 3738 11928 6054
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11992 5234 12020 5782
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11992 4758 12020 5170
rect 12084 5166 12112 10406
rect 12176 7410 12204 11018
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 6118 12204 7142
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12176 4826 12204 6054
rect 12268 5710 12296 10542
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12360 8362 12388 10474
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12360 7954 12388 8298
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12452 6798 12480 11494
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9450 12572 9862
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12544 8090 12572 9386
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12636 7886 12664 9930
rect 12728 9586 12756 10406
rect 12820 9994 12848 11086
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7478 12664 7822
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12452 5914 12480 6734
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6322 12572 6598
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12452 4826 12480 5714
rect 12544 5642 12572 6258
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 11992 4214 12020 4694
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11060 3596 11112 3602
rect 10980 3556 11060 3584
rect 11060 3538 11112 3544
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 2650 10916 3470
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11072 2582 11100 3538
rect 11624 3058 11652 3538
rect 12636 3466 12664 5306
rect 12728 4214 12756 9318
rect 12820 8838 12848 9930
rect 12808 8832 12860 8838
rect 12912 8809 12940 10610
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 13004 9382 13032 10134
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13096 8974 13124 10950
rect 13268 10260 13320 10266
rect 13372 10248 13400 11630
rect 13464 11558 13492 12242
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14108 11898 14136 12038
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14108 11626 14136 11834
rect 14292 11694 14320 12038
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 10266 13492 11494
rect 14108 11218 14136 11562
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 13320 10220 13400 10248
rect 13268 10202 13320 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 9654 13216 9862
rect 13176 9648 13228 9654
rect 13176 9590 13228 9596
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12808 8774 12860 8780
rect 12898 8800 12954 8809
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12820 4154 12848 8774
rect 12898 8735 12954 8744
rect 13096 8566 13124 8910
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12912 8022 12940 8298
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12912 7546 12940 7958
rect 13096 7818 13124 8230
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6934 12940 7142
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12912 6458 12940 6870
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13084 5364 13136 5370
rect 13188 5352 13216 9590
rect 13280 9450 13308 10066
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13372 6798 13400 10220
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8634 13492 9046
rect 13556 8974 13584 9454
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13556 8022 13584 8910
rect 13648 8906 13676 11154
rect 14108 10742 14136 11154
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14108 10266 14136 10678
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14200 9926 14228 10542
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13740 7834 13768 9522
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13464 7806 13768 7834
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13372 5846 13400 6190
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13136 5324 13216 5352
rect 13084 5306 13136 5312
rect 13464 4826 13492 7806
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 6934 13584 7686
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13556 6322 13584 6870
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13556 5710 13584 5850
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13556 5166 13584 5510
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12820 4126 12940 4154
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 12544 2990 12572 3334
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 12544 2514 12572 2926
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12636 2394 12664 3402
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12728 3097 12756 3130
rect 12714 3088 12770 3097
rect 12714 3023 12770 3032
rect 12728 2990 12756 3023
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12820 2650 12848 3538
rect 12912 3516 12940 4126
rect 13004 3942 13032 4422
rect 13096 4146 13124 4762
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3670 13032 3878
rect 13096 3670 13124 4082
rect 13556 3942 13584 5102
rect 13648 4078 13676 6666
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13740 4758 13768 5578
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13832 4486 13860 9386
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14844 9042 14872 10474
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13648 3738 13676 4014
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13832 3670 13860 4150
rect 13924 4078 13952 6326
rect 14186 6216 14242 6225
rect 14004 6180 14056 6186
rect 14186 6151 14242 6160
rect 14004 6122 14056 6128
rect 14016 5846 14044 6122
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14016 4826 14044 5782
rect 14200 4826 14228 6151
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14660 5914 14688 8298
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 7993 14780 8230
rect 14844 8090 14872 8978
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14738 7984 14794 7993
rect 15028 7954 15056 11562
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 8430 15240 11086
rect 15488 9994 15516 11766
rect 15752 11620 15804 11626
rect 15752 11562 15804 11568
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 14738 7919 14794 7928
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14752 7342 14780 7822
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14752 7002 14780 7278
rect 15028 7002 15056 7890
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15304 6866 15332 9862
rect 15488 9722 15516 9930
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15672 9586 15700 11086
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15672 8294 15700 9114
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 8090 15700 8230
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15672 7546 15700 8026
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13820 3664 13872 3670
rect 14016 3641 14044 3674
rect 13820 3606 13872 3612
rect 14002 3632 14058 3641
rect 13176 3528 13228 3534
rect 12912 3488 13176 3516
rect 13176 3470 13228 3476
rect 13188 3194 13216 3470
rect 13832 3398 13860 3606
rect 13912 3596 13964 3602
rect 14002 3567 14058 3576
rect 13912 3538 13964 3544
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13280 2650 13308 3062
rect 13740 2854 13768 3062
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13740 2514 13768 2790
rect 13924 2514 13952 3538
rect 14200 2990 14228 4762
rect 14660 4622 14688 5850
rect 15396 5778 15424 6734
rect 15488 6497 15516 6802
rect 15474 6488 15530 6497
rect 15474 6423 15530 6432
rect 15488 6118 15516 6423
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15384 5772 15436 5778
rect 15212 5732 15384 5760
rect 15212 5166 15240 5732
rect 15384 5714 15436 5720
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15304 4690 15332 5306
rect 15488 5273 15516 6054
rect 15658 5536 15714 5545
rect 15764 5522 15792 11562
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 10130 16528 10542
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16316 9674 16344 9998
rect 16500 9722 16528 10066
rect 16488 9716 16540 9722
rect 16316 9646 16436 9674
rect 16488 9658 16540 9664
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15714 5494 15792 5522
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15658 5471 15714 5480
rect 15474 5264 15530 5273
rect 15384 5228 15436 5234
rect 15672 5234 15700 5471
rect 15474 5199 15530 5208
rect 15660 5228 15712 5234
rect 15384 5170 15436 5176
rect 15660 5170 15712 5176
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 14738 4312 14794 4321
rect 14738 4247 14794 4256
rect 14648 4004 14700 4010
rect 14752 3992 14780 4247
rect 15120 4078 15148 4558
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4078 15240 4422
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 14700 3964 14780 3992
rect 14924 4004 14976 4010
rect 14648 3946 14700 3952
rect 14924 3946 14976 3952
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14016 2650 14044 2926
rect 14660 2854 14688 3470
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14752 2990 14780 3334
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 12636 2366 13032 2394
rect 12636 2310 12664 2366
rect 13004 2310 13032 2366
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 12268 1329 12296 2246
rect 12254 1320 12310 1329
rect 12254 1255 12310 1264
rect 10506 54 10824 82
rect 12806 82 12862 480
rect 12912 82 12940 2246
rect 14108 1601 14136 2790
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 14660 2310 14688 2790
rect 14752 2650 14780 2926
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 1873 14872 2246
rect 14830 1864 14886 1873
rect 14830 1799 14886 1808
rect 14094 1592 14150 1601
rect 14094 1527 14150 1536
rect 12806 54 12940 82
rect 14936 82 14964 3946
rect 15120 3398 15148 4014
rect 15304 4010 15332 4626
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15396 3913 15424 5170
rect 15856 5098 15884 5510
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15752 4276 15804 4282
rect 15948 4264 15976 9318
rect 16132 9178 16160 9386
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7274 16160 8230
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16040 5778 16068 7210
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16224 5914 16252 6122
rect 16316 5914 16344 8774
rect 16408 7002 16436 9646
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16500 8022 16528 8434
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16500 7410 16528 7958
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16408 6322 16436 6938
rect 16592 6866 16620 10474
rect 16684 10470 16712 11154
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 9450 16712 10406
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16684 8838 16712 9386
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16684 7410 16712 8774
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16592 6458 16620 6802
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 16224 5370 16252 5850
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16120 4276 16172 4282
rect 15948 4236 16120 4264
rect 15752 4218 15804 4224
rect 16120 4218 16172 4224
rect 15764 4185 15792 4218
rect 15750 4176 15806 4185
rect 15750 4111 15806 4120
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 15672 3602 15700 4014
rect 16132 3942 16160 4218
rect 16500 4214 16528 4422
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16026 3768 16082 3777
rect 16026 3703 16082 3712
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15212 2650 15240 3062
rect 15580 2854 15608 3334
rect 16040 3058 16068 3703
rect 16132 3194 16160 3878
rect 16316 3398 16344 4082
rect 16500 3466 16528 4150
rect 16684 4146 16712 4558
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15212 2514 15240 2586
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15672 2310 15700 2926
rect 16132 2378 16160 3130
rect 16500 3126 16528 3402
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16592 2689 16620 3946
rect 16684 3534 16712 4082
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16776 3058 16804 12718
rect 17314 11792 17370 11801
rect 17314 11727 17370 11736
rect 17328 11694 17356 11727
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19260 11558 19288 11630
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 18510 11248 18566 11257
rect 18510 11183 18512 11192
rect 18564 11183 18566 11192
rect 18512 11154 18564 11160
rect 18524 10810 18552 11154
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18524 10713 18552 10746
rect 18326 10704 18382 10713
rect 17684 10668 17736 10674
rect 18326 10639 18382 10648
rect 18510 10704 18566 10713
rect 18510 10639 18566 10648
rect 17684 10610 17736 10616
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16868 7818 16896 8366
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16960 7546 16988 8230
rect 17144 8022 17172 10406
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17420 8294 17448 9046
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 8090 17448 8230
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17144 7546 17172 7958
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16960 6934 16988 7482
rect 17132 7200 17184 7206
rect 17236 7188 17264 7958
rect 17184 7160 17264 7188
rect 17132 7142 17184 7148
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 16960 6186 16988 6870
rect 17144 6662 17172 7142
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16868 5166 16896 5850
rect 17512 5846 17540 9658
rect 17696 9024 17724 10610
rect 18340 10606 18368 10639
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17788 9722 17816 10066
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17880 9382 17908 10066
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17776 9036 17828 9042
rect 17696 8996 17776 9024
rect 17776 8978 17828 8984
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17788 8022 17816 8502
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17880 7868 17908 9318
rect 17972 8537 18000 10542
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18248 9518 18276 9930
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 17958 8528 18014 8537
rect 18064 8498 18092 9046
rect 17958 8463 18014 8472
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 17788 7840 17908 7868
rect 17788 7478 17816 7840
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17500 5840 17552 5846
rect 17500 5782 17552 5788
rect 17512 5370 17540 5782
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 16960 4826 16988 4966
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16960 4486 16988 4762
rect 17696 4758 17724 4966
rect 17500 4752 17552 4758
rect 17500 4694 17552 4700
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17144 4282 17172 4422
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17144 3126 17172 3470
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16578 2680 16634 2689
rect 17328 2650 17356 4422
rect 17512 4049 17540 4694
rect 17498 4040 17554 4049
rect 17554 3984 17632 3992
rect 17498 3975 17500 3984
rect 17552 3964 17632 3984
rect 17500 3946 17552 3952
rect 17512 3915 17540 3946
rect 17604 2650 17632 3964
rect 17788 2922 17816 7414
rect 18156 7410 18184 9318
rect 18248 9178 18276 9454
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18432 7750 18460 8298
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17880 6934 17908 7210
rect 18156 7002 18184 7346
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17880 6186 17908 6598
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18234 5128 18290 5137
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17880 3466 17908 4150
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 16578 2615 16634 2624
rect 17316 2644 17368 2650
rect 16592 2514 16620 2615
rect 17316 2586 17368 2592
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 17788 2378 17816 2858
rect 17972 2514 18000 4490
rect 18064 3670 18092 5102
rect 18234 5063 18290 5072
rect 18248 5030 18276 5063
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18156 4282 18184 4762
rect 18524 4690 18552 9998
rect 18616 5692 18644 10474
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18708 7954 18736 9114
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7002 18736 7890
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18800 6798 18828 11494
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18892 9110 18920 9454
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 6934 18920 7686
rect 18984 6934 19012 10950
rect 19260 10674 19288 11494
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19444 10452 19472 11154
rect 19536 11121 19564 11290
rect 19522 11112 19578 11121
rect 19522 11047 19578 11056
rect 19524 10464 19576 10470
rect 19444 10424 19524 10452
rect 19524 10406 19576 10412
rect 19536 10169 19564 10406
rect 19522 10160 19578 10169
rect 19340 10124 19392 10130
rect 19522 10095 19578 10104
rect 19340 10066 19392 10072
rect 19352 9897 19380 10066
rect 19338 9888 19394 9897
rect 19338 9823 19394 9832
rect 19352 9722 19380 9823
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8566 19288 8910
rect 19628 8634 19656 15558
rect 19982 15520 20038 15558
rect 33060 15558 33378 15586
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 32220 12776 32272 12782
rect 32220 12718 32272 12724
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18800 6390 18828 6734
rect 18892 6458 18920 6870
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18788 6180 18840 6186
rect 18984 6168 19012 6870
rect 18840 6140 19012 6168
rect 18788 6122 18840 6128
rect 19076 5710 19104 8502
rect 19720 8498 19748 9862
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19260 7274 19288 8026
rect 19628 7546 19656 8230
rect 19720 8090 19748 8434
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 18696 5704 18748 5710
rect 18616 5664 18696 5692
rect 18696 5646 18748 5652
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 18708 5370 18736 5646
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 19076 5302 19104 5646
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18340 4214 18368 4422
rect 18328 4208 18380 4214
rect 19168 4185 19196 4422
rect 18328 4150 18380 4156
rect 19154 4176 19210 4185
rect 19154 4111 19210 4120
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18234 4040 18290 4049
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 2990 18092 3334
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15198 82 15254 480
rect 14936 54 15254 82
rect 8114 0 8170 54
rect 10506 0 10562 54
rect 12806 0 12862 54
rect 15198 0 15254 54
rect 17590 82 17646 480
rect 17972 82 18000 2450
rect 18156 2446 18184 4014
rect 18234 3975 18290 3984
rect 18248 3670 18276 3975
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18340 3398 18368 3674
rect 18984 3641 19012 3674
rect 18970 3632 19026 3641
rect 18970 3567 18972 3576
rect 19024 3567 19026 3576
rect 18972 3538 19024 3544
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 2990 18368 3334
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18340 2582 18368 2790
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18984 2378 19012 3538
rect 19168 2514 19196 4111
rect 19260 4060 19288 5170
rect 19352 5098 19380 7142
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 6186 19472 6734
rect 19812 6458 19840 10950
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 7410 19932 9318
rect 19996 8906 20024 9454
rect 20088 9178 20116 10406
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9518 20208 9862
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19996 7886 20024 8842
rect 20088 8498 20116 9114
rect 20180 9042 20208 9454
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19904 7002 19932 7346
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 20180 6662 20208 8978
rect 20272 8566 20300 10542
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 9722 20852 10066
rect 21548 10056 21600 10062
rect 21548 9998 21600 10004
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20548 8498 20576 9522
rect 21284 9110 21312 9862
rect 21468 9450 21496 9862
rect 21560 9450 21588 9998
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21468 9178 21496 9386
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21364 9104 21416 9110
rect 21364 9046 21416 9052
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21284 8634 21312 9046
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20548 7478 20576 8434
rect 21272 8424 21324 8430
rect 21376 8412 21404 9046
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21468 8498 21496 8774
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21324 8384 21404 8412
rect 21272 8366 21324 8372
rect 21560 8362 21588 9386
rect 21652 8673 21680 9658
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21638 8664 21694 8673
rect 21638 8599 21694 8608
rect 21744 8498 21772 8910
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21548 8356 21600 8362
rect 21548 8298 21600 8304
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20824 7954 20852 8230
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21284 7546 21312 7958
rect 21836 7886 21864 9862
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 21928 7274 21956 7482
rect 21916 7268 21968 7274
rect 21916 7210 21968 7216
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 20272 6118 20300 6802
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19536 4321 19564 6054
rect 20456 5846 20484 6122
rect 20732 6118 20760 6734
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20996 6180 21048 6186
rect 20996 6122 21048 6128
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19628 5234 19656 5510
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19720 4758 19748 5034
rect 20548 5030 20576 5782
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4826 20576 4966
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 19708 4752 19760 4758
rect 19708 4694 19760 4700
rect 19522 4312 19578 4321
rect 19720 4282 19748 4694
rect 19522 4247 19578 4256
rect 19708 4276 19760 4282
rect 19260 4032 19472 4060
rect 19444 2836 19472 4032
rect 19536 3738 19564 4247
rect 19708 4218 19760 4224
rect 19720 3942 19748 4218
rect 20640 4078 20668 5510
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 20628 4072 20680 4078
rect 20732 4049 20760 6054
rect 21008 5710 21036 6122
rect 21640 5840 21692 5846
rect 21640 5782 21692 5788
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21468 5302 21496 5510
rect 21652 5302 21680 5782
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21824 5636 21876 5642
rect 21824 5578 21876 5584
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21652 4758 21680 5238
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 20824 4282 20852 4694
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21284 4282 21312 4558
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 21100 4049 21128 4082
rect 20628 4014 20680 4020
rect 20718 4040 20774 4049
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19628 3058 19656 3538
rect 19616 3052 19668 3058
rect 19616 2994 19668 3000
rect 19628 2922 19656 2994
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19524 2848 19576 2854
rect 19444 2808 19524 2836
rect 19524 2790 19576 2796
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 17590 54 18000 82
rect 19720 82 19748 3878
rect 19904 3670 19932 4014
rect 20718 3975 20774 3984
rect 21086 4040 21142 4049
rect 21086 3975 21142 3984
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 20824 3194 20852 3674
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 21284 3194 21312 3470
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 19800 2916 19852 2922
rect 19800 2858 19852 2864
rect 19812 2582 19840 2858
rect 21284 2689 21312 3130
rect 21270 2680 21326 2689
rect 21376 2650 21404 4150
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21744 3398 21772 4014
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21270 2615 21326 2624
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 19800 2576 19852 2582
rect 19800 2518 19852 2524
rect 21744 2378 21772 3334
rect 21836 3194 21864 5578
rect 21928 4826 21956 5646
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 22020 4154 22048 11562
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 26976 11212 27028 11218
rect 26976 11154 27028 11160
rect 22664 10810 22692 11154
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 26238 10976 26294 10985
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22374 10568 22430 10577
rect 22374 10503 22430 10512
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22112 8090 22140 10406
rect 22388 10130 22416 10503
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22388 9722 22416 10066
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 22204 8362 22232 8910
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22204 8090 22232 8298
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22112 7410 22140 8026
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22480 6934 22508 9318
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 7002 22600 7142
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22284 6656 22336 6662
rect 22284 6598 22336 6604
rect 22098 6352 22154 6361
rect 22098 6287 22154 6296
rect 22112 6254 22140 6287
rect 22296 6254 22324 6598
rect 22388 6322 22416 6734
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22112 5642 22140 6190
rect 22296 5710 22324 6190
rect 22388 5914 22416 6258
rect 22572 6118 22600 6938
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22664 5846 22692 10746
rect 23020 10532 23072 10538
rect 23020 10474 23072 10480
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 22940 9382 22968 10066
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22756 8634 22784 8978
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22756 8537 22784 8570
rect 22742 8528 22798 8537
rect 22742 8463 22798 8472
rect 22836 8016 22888 8022
rect 22836 7958 22888 7964
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22756 7478 22784 7822
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22756 6866 22784 7414
rect 22848 7274 22876 7958
rect 22836 7268 22888 7274
rect 22836 7210 22888 7216
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22652 5840 22704 5846
rect 22652 5782 22704 5788
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 22296 5030 22324 5646
rect 22756 5370 22784 6054
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22296 4214 22324 4966
rect 22572 4622 22600 4966
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22284 4208 22336 4214
rect 22020 4126 22140 4154
rect 22284 4150 22336 4156
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 22020 3738 22048 3878
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 21836 2922 21864 3130
rect 21824 2916 21876 2922
rect 21824 2858 21876 2864
rect 21732 2372 21784 2378
rect 21732 2314 21784 2320
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 19890 82 19946 480
rect 19720 54 19946 82
rect 22112 82 22140 4126
rect 22296 4078 22324 4150
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22756 3738 22784 5306
rect 23032 4554 23060 10474
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23400 9382 23428 9862
rect 23938 9616 23994 9625
rect 23938 9551 23994 9560
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 23020 4548 23072 4554
rect 23020 4490 23072 4496
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22756 3194 22784 3674
rect 23124 3466 23152 8774
rect 23400 8537 23428 8842
rect 23386 8528 23442 8537
rect 23386 8463 23442 8472
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23216 7002 23244 7142
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23400 6225 23428 8366
rect 23386 6216 23442 6225
rect 23386 6151 23442 6160
rect 23400 4690 23428 6151
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23492 5914 23520 6054
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23492 5234 23520 5850
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23676 4690 23704 9386
rect 23952 9042 23980 9551
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24136 9042 24164 9454
rect 24412 9178 24440 10066
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 23940 9036 23992 9042
rect 23940 8978 23992 8984
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 23952 8634 23980 8978
rect 24412 8838 24440 9114
rect 24400 8832 24452 8838
rect 24400 8774 24452 8780
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23768 7410 23796 8026
rect 23952 7857 23980 8570
rect 24308 8424 24360 8430
rect 24308 8366 24360 8372
rect 24320 8090 24348 8366
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24124 7880 24176 7886
rect 23938 7848 23994 7857
rect 24124 7822 24176 7828
rect 23938 7783 23994 7792
rect 24136 7410 24164 7822
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 23756 7268 23808 7274
rect 23756 7210 23808 7216
rect 23768 7002 23796 7210
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23768 5914 23796 6190
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23860 5846 23888 6598
rect 23848 5840 23900 5846
rect 23848 5782 23900 5788
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24044 4758 24072 5646
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 23388 4684 23440 4690
rect 23216 4644 23388 4672
rect 23216 4214 23244 4644
rect 23388 4626 23440 4632
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 23204 4208 23256 4214
rect 23204 4150 23256 4156
rect 23112 3460 23164 3466
rect 23112 3402 23164 3408
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 23308 2961 23336 4490
rect 23676 4282 23704 4626
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23664 4276 23716 4282
rect 23664 4218 23716 4224
rect 23400 2990 23428 4218
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23492 3194 23520 3674
rect 23676 3670 23704 3878
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 24136 3466 24164 7346
rect 24400 6928 24452 6934
rect 24400 6870 24452 6876
rect 24412 6458 24440 6870
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24412 5914 24440 6394
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 24320 4826 24348 5102
rect 24412 5098 24440 5850
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24412 4282 24440 5034
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24398 3632 24454 3641
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 24228 3194 24256 3606
rect 24398 3567 24454 3576
rect 24412 3534 24440 3567
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 23388 2984 23440 2990
rect 23294 2952 23350 2961
rect 23388 2926 23440 2932
rect 23294 2887 23350 2896
rect 23400 2446 23428 2926
rect 24412 2922 24440 3334
rect 24400 2916 24452 2922
rect 24400 2858 24452 2864
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 22282 82 22338 480
rect 22112 54 22338 82
rect 24504 82 24532 10950
rect 26238 10911 26294 10920
rect 26252 10810 26280 10911
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 25502 10704 25558 10713
rect 25502 10639 25558 10648
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24674 8528 24730 8537
rect 24674 8463 24730 8472
rect 24688 7954 24716 8463
rect 24780 8430 24808 9862
rect 25056 9489 25084 10542
rect 25516 10130 25544 10639
rect 26252 10606 26280 10746
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 25504 10124 25556 10130
rect 25504 10066 25556 10072
rect 25516 9761 25544 10066
rect 25502 9752 25558 9761
rect 25502 9687 25558 9696
rect 25516 9654 25544 9687
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25042 9480 25098 9489
rect 24860 9444 24912 9450
rect 25042 9415 25098 9424
rect 24860 9386 24912 9392
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24584 7812 24636 7818
rect 24584 7754 24636 7760
rect 24596 4049 24624 7754
rect 24688 7546 24716 7890
rect 24780 7886 24808 8366
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24688 6390 24716 7482
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 24688 4672 24716 6326
rect 24780 6254 24808 7822
rect 24872 6322 24900 9386
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25240 8634 25268 8978
rect 25228 8628 25280 8634
rect 25228 8570 25280 8576
rect 25240 8022 25268 8570
rect 25228 8016 25280 8022
rect 25228 7958 25280 7964
rect 25424 7954 25452 8978
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 25424 7342 25452 7890
rect 25608 7410 25636 8910
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25884 8090 25912 8366
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 25240 5914 25268 6258
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 25424 5914 25452 6122
rect 25884 6118 25912 7142
rect 25872 6112 25924 6118
rect 25872 6054 25924 6060
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25976 5710 26004 10406
rect 26620 9722 26648 10542
rect 26988 10470 27016 11154
rect 29092 11008 29144 11014
rect 29092 10950 29144 10956
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 27988 10600 28040 10606
rect 27894 10568 27950 10577
rect 27950 10548 27988 10554
rect 28092 10577 28120 10610
rect 27950 10542 28040 10548
rect 28078 10568 28134 10577
rect 27950 10526 28028 10542
rect 27894 10503 27950 10512
rect 28078 10503 28134 10512
rect 28632 10532 28684 10538
rect 28632 10474 28684 10480
rect 26976 10464 27028 10470
rect 26976 10406 27028 10412
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 26988 10033 27016 10406
rect 27264 10266 27292 10406
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 27160 10056 27212 10062
rect 26974 10024 27030 10033
rect 27160 9998 27212 10004
rect 26974 9959 27030 9968
rect 27068 9988 27120 9994
rect 26608 9716 26660 9722
rect 26608 9658 26660 9664
rect 26620 9081 26648 9658
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26712 9178 26740 9318
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26606 9072 26662 9081
rect 26606 9007 26662 9016
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26068 7002 26096 7346
rect 26344 7274 26372 7346
rect 26332 7268 26384 7274
rect 26332 7210 26384 7216
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26620 6769 26648 6802
rect 26606 6760 26662 6769
rect 26606 6695 26662 6704
rect 26620 6322 26648 6695
rect 26712 6338 26740 8842
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26804 8090 26832 8230
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 26804 7410 26832 8026
rect 26896 7426 26924 9318
rect 26988 8945 27016 9959
rect 27068 9930 27120 9936
rect 26974 8936 27030 8945
rect 26974 8871 27030 8880
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26988 7546 27016 8230
rect 26976 7540 27028 7546
rect 26976 7482 27028 7488
rect 26792 7404 26844 7410
rect 26896 7398 27016 7426
rect 26792 7346 26844 7352
rect 26884 6452 26936 6458
rect 26884 6394 26936 6400
rect 26896 6361 26924 6394
rect 26882 6352 26938 6361
rect 26608 6316 26660 6322
rect 26712 6310 26832 6338
rect 26608 6258 26660 6264
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 24964 5370 24992 5510
rect 24952 5364 25004 5370
rect 24952 5306 25004 5312
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24768 4684 24820 4690
rect 24688 4644 24768 4672
rect 24688 4214 24716 4644
rect 24768 4626 24820 4632
rect 24872 4214 24900 5170
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 24676 4208 24728 4214
rect 24676 4150 24728 4156
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24582 4040 24638 4049
rect 24582 3975 24638 3984
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 24780 2650 24808 2926
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24872 2582 24900 4150
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24964 3398 24992 4014
rect 25148 3738 25176 4558
rect 25424 3913 25452 4966
rect 25976 4826 26004 5646
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 26068 5234 26096 5510
rect 26160 5234 26188 6054
rect 26056 5228 26108 5234
rect 26056 5170 26108 5176
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 25964 4820 26016 4826
rect 25964 4762 26016 4768
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25410 3904 25466 3913
rect 25410 3839 25466 3848
rect 25976 3738 26004 4558
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 26056 3664 26108 3670
rect 26056 3606 26108 3612
rect 25412 3460 25464 3466
rect 25412 3402 25464 3408
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 25424 2650 25452 3402
rect 26068 3194 26096 3606
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 24860 2576 24912 2582
rect 24860 2518 24912 2524
rect 26160 2446 26188 3878
rect 26252 3738 26280 4218
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26344 2650 26372 3470
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26528 1193 26556 2246
rect 26620 1465 26648 6258
rect 26700 5840 26752 5846
rect 26700 5782 26752 5788
rect 26712 5370 26740 5782
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 26700 4752 26752 4758
rect 26700 4694 26752 4700
rect 26712 4282 26740 4694
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26804 3534 26832 6310
rect 26882 6287 26938 6296
rect 26884 6180 26936 6186
rect 26884 6122 26936 6128
rect 26896 5302 26924 6122
rect 26988 5681 27016 7398
rect 26974 5672 27030 5681
rect 26974 5607 27030 5616
rect 27080 5574 27108 9930
rect 27172 8838 27200 9998
rect 27264 9586 27292 10202
rect 27436 10192 27488 10198
rect 27436 10134 27488 10140
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 27252 9580 27304 9586
rect 27252 9522 27304 9528
rect 27356 9110 27384 9590
rect 27448 9450 27476 10134
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 27436 9444 27488 9450
rect 27436 9386 27488 9392
rect 28080 9444 28132 9450
rect 28080 9386 28132 9392
rect 27344 9104 27396 9110
rect 27344 9046 27396 9052
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27172 7478 27200 8774
rect 27356 8022 27384 9046
rect 27448 8090 27476 9386
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 27528 9104 27580 9110
rect 27528 9046 27580 9052
rect 27712 9104 27764 9110
rect 27712 9046 27764 9052
rect 27540 8294 27568 9046
rect 27724 8498 27752 9046
rect 28092 8974 28120 9386
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 27804 8628 27856 8634
rect 27804 8570 27856 8576
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27816 8362 27844 8570
rect 27804 8356 27856 8362
rect 27856 8316 28028 8344
rect 27804 8298 27856 8304
rect 27528 8288 27580 8294
rect 27528 8230 27580 8236
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 28000 8090 28028 8316
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 27344 8016 27396 8022
rect 27344 7958 27396 7964
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27160 7472 27212 7478
rect 27160 7414 27212 7420
rect 27540 7002 27568 7686
rect 27632 7546 27660 7822
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27540 6322 27568 6598
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27252 6180 27304 6186
rect 27252 6122 27304 6128
rect 27264 5710 27292 6122
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 27068 5568 27120 5574
rect 27068 5510 27120 5516
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 26896 3670 26924 5238
rect 27080 5234 27108 5510
rect 27264 5234 27292 5646
rect 27068 5228 27120 5234
rect 27068 5170 27120 5176
rect 27252 5228 27304 5234
rect 27252 5170 27304 5176
rect 27264 4622 27292 5170
rect 27252 4616 27304 4622
rect 27252 4558 27304 4564
rect 27160 4548 27212 4554
rect 27160 4490 27212 4496
rect 26884 3664 26936 3670
rect 26884 3606 26936 3612
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 27172 3126 27200 4490
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27356 3670 27384 3878
rect 27344 3664 27396 3670
rect 27344 3606 27396 3612
rect 27436 3392 27488 3398
rect 27436 3334 27488 3340
rect 27160 3120 27212 3126
rect 27160 3062 27212 3068
rect 27448 2514 27476 3334
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27540 2310 27568 6258
rect 27816 6186 27844 6734
rect 27804 6180 27856 6186
rect 27804 6122 27856 6128
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 28184 5710 28212 9862
rect 28644 9178 28672 10474
rect 28724 10124 28776 10130
rect 28724 10066 28776 10072
rect 28736 9382 28764 10066
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28632 9172 28684 9178
rect 28632 9114 28684 9120
rect 28644 8974 28672 9114
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28448 8560 28500 8566
rect 28262 8528 28318 8537
rect 28448 8502 28500 8508
rect 28262 8463 28318 8472
rect 28276 7449 28304 8463
rect 28460 7993 28488 8502
rect 28552 8362 28580 8910
rect 28540 8356 28592 8362
rect 28540 8298 28592 8304
rect 28446 7984 28502 7993
rect 28446 7919 28502 7928
rect 28552 7886 28580 8298
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28262 7440 28318 7449
rect 28262 7375 28318 7384
rect 28276 7342 28304 7375
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 28448 7268 28500 7274
rect 28448 7210 28500 7216
rect 28264 5840 28316 5846
rect 28264 5782 28316 5788
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28184 5234 28212 5510
rect 28276 5370 28304 5782
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 28368 5370 28396 5646
rect 28460 5556 28488 7210
rect 28552 7002 28580 7822
rect 28644 7546 28672 7958
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 28644 7002 28672 7482
rect 28540 6996 28592 7002
rect 28540 6938 28592 6944
rect 28632 6996 28684 7002
rect 28632 6938 28684 6944
rect 28632 5568 28684 5574
rect 28460 5528 28632 5556
rect 28632 5510 28684 5516
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 28356 5364 28408 5370
rect 28356 5306 28408 5312
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28184 4622 28212 5170
rect 28264 4752 28316 4758
rect 28264 4694 28316 4700
rect 28172 4616 28224 4622
rect 28078 4584 28134 4593
rect 28172 4558 28224 4564
rect 28078 4519 28134 4528
rect 28092 3913 28120 4519
rect 28184 3942 28212 4558
rect 28276 4282 28304 4694
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 28356 4004 28408 4010
rect 28356 3946 28408 3952
rect 28172 3936 28224 3942
rect 28078 3904 28134 3913
rect 27622 3836 27918 3856
rect 28172 3878 28224 3884
rect 28078 3839 28134 3848
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 28092 2990 28120 3674
rect 28368 3670 28396 3946
rect 28356 3664 28408 3670
rect 28356 3606 28408 3612
rect 28172 3528 28224 3534
rect 28172 3470 28224 3476
rect 28080 2984 28132 2990
rect 28080 2926 28132 2932
rect 28184 2854 28212 3470
rect 28368 3194 28396 3606
rect 28356 3188 28408 3194
rect 28356 3130 28408 3136
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 28184 2582 28212 2790
rect 28172 2576 28224 2582
rect 28172 2518 28224 2524
rect 28644 2514 28672 5510
rect 28736 4593 28764 9318
rect 29000 9104 29052 9110
rect 29000 9046 29052 9052
rect 29012 8634 29040 9046
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 28816 6928 28868 6934
rect 28816 6870 28868 6876
rect 28828 6118 28856 6870
rect 28920 6225 28948 7414
rect 28906 6216 28962 6225
rect 28906 6151 28962 6160
rect 28816 6112 28868 6118
rect 28816 6054 28868 6060
rect 28722 4584 28778 4593
rect 28722 4519 28778 4528
rect 28816 4548 28868 4554
rect 28816 4490 28868 4496
rect 28828 3097 28856 4490
rect 28920 4146 28948 6151
rect 29104 5098 29132 10950
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29196 8974 29224 9998
rect 32232 9722 32260 12718
rect 33060 11121 33088 15558
rect 33322 15520 33378 15558
rect 35530 15056 35586 15065
rect 35530 14991 35586 15000
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 34152 11212 34204 11218
rect 34152 11154 34204 11160
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 33046 11112 33102 11121
rect 33046 11047 33102 11056
rect 34164 10985 34192 11154
rect 34150 10976 34206 10985
rect 34150 10911 34206 10920
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 34624 10470 34652 11154
rect 35452 10810 35480 11154
rect 35440 10804 35492 10810
rect 35440 10746 35492 10752
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 35360 10577 35388 10610
rect 35346 10568 35402 10577
rect 35346 10503 35402 10512
rect 33048 10464 33100 10470
rect 33048 10406 33100 10412
rect 33692 10464 33744 10470
rect 33692 10406 33744 10412
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 35164 10464 35216 10470
rect 35164 10406 35216 10412
rect 32220 9716 32272 9722
rect 32220 9658 32272 9664
rect 29826 9616 29882 9625
rect 29826 9551 29882 9560
rect 29840 9518 29868 9551
rect 29828 9512 29880 9518
rect 29828 9454 29880 9460
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 29184 8968 29236 8974
rect 29184 8910 29236 8916
rect 29196 8498 29224 8910
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 29196 7410 29224 8434
rect 29368 8356 29420 8362
rect 29368 8298 29420 8304
rect 29380 7750 29408 8298
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 29196 7002 29224 7346
rect 30024 7274 30052 7822
rect 30300 7818 30328 9454
rect 32404 9444 32456 9450
rect 32404 9386 32456 9392
rect 30656 9376 30708 9382
rect 30656 9318 30708 9324
rect 30380 9036 30432 9042
rect 30380 8978 30432 8984
rect 30392 8294 30420 8978
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 30392 7818 30420 8230
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 30380 7812 30432 7818
rect 30380 7754 30432 7760
rect 29460 7268 29512 7274
rect 29460 7210 29512 7216
rect 30012 7268 30064 7274
rect 30012 7210 30064 7216
rect 29472 7002 29500 7210
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 29460 6996 29512 7002
rect 29460 6938 29512 6944
rect 29552 6792 29604 6798
rect 29552 6734 29604 6740
rect 29564 5914 29592 6734
rect 29736 6248 29788 6254
rect 29736 6190 29788 6196
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29748 5574 29776 6190
rect 29736 5568 29788 5574
rect 29736 5510 29788 5516
rect 29092 5092 29144 5098
rect 29092 5034 29144 5040
rect 29104 4826 29132 5034
rect 29092 4820 29144 4826
rect 29092 4762 29144 4768
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29092 3936 29144 3942
rect 29092 3878 29144 3884
rect 28814 3088 28870 3097
rect 28814 3023 28870 3032
rect 29012 2582 29040 3878
rect 29104 3738 29132 3878
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 29380 3398 29408 4014
rect 29460 3460 29512 3466
rect 29460 3402 29512 3408
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29472 2922 29500 3402
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 29460 2916 29512 2922
rect 29460 2858 29512 2864
rect 29000 2576 29052 2582
rect 29000 2518 29052 2524
rect 28632 2508 28684 2514
rect 28632 2450 28684 2456
rect 27528 2304 27580 2310
rect 27528 2246 27580 2252
rect 26606 1456 26662 1465
rect 26606 1391 26662 1400
rect 26514 1184 26570 1193
rect 26514 1119 26570 1128
rect 24582 82 24638 480
rect 24504 54 24638 82
rect 17590 0 17646 54
rect 19890 0 19946 54
rect 22282 0 22338 54
rect 24582 0 24638 54
rect 26974 82 27030 480
rect 27250 368 27306 377
rect 27250 303 27306 312
rect 27264 82 27292 303
rect 26974 54 27292 82
rect 29104 82 29132 2858
rect 29472 2650 29500 2858
rect 29564 2650 29592 4082
rect 30024 3058 30052 7210
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30196 5092 30248 5098
rect 30196 5034 30248 5040
rect 30104 4004 30156 4010
rect 30104 3946 30156 3952
rect 30116 3738 30144 3946
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 30208 3466 30236 5034
rect 30196 3460 30248 3466
rect 30196 3402 30248 3408
rect 30208 3194 30236 3402
rect 30300 3194 30328 7142
rect 30392 6905 30420 7754
rect 30484 7206 30512 7890
rect 30472 7200 30524 7206
rect 30472 7142 30524 7148
rect 30668 7002 30696 9318
rect 32312 9036 32364 9042
rect 32312 8978 32364 8984
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31404 8430 31432 8774
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 31312 7342 31340 7890
rect 31404 7410 31432 8366
rect 32324 8294 32352 8978
rect 32312 8288 32364 8294
rect 32312 8230 32364 8236
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 30656 6996 30708 7002
rect 30656 6938 30708 6944
rect 30378 6896 30434 6905
rect 30378 6831 30434 6840
rect 31312 6798 31340 7278
rect 31576 6996 31628 7002
rect 31576 6938 31628 6944
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31208 6248 31260 6254
rect 31208 6190 31260 6196
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 30392 5846 30420 6054
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30484 5030 30512 5646
rect 31024 5364 31076 5370
rect 31024 5306 31076 5312
rect 30840 5160 30892 5166
rect 30840 5102 30892 5108
rect 30472 5024 30524 5030
rect 30472 4966 30524 4972
rect 30380 4684 30432 4690
rect 30380 4626 30432 4632
rect 30392 4214 30420 4626
rect 30380 4208 30432 4214
rect 30380 4150 30432 4156
rect 30392 3602 30420 4150
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 30196 3188 30248 3194
rect 30196 3130 30248 3136
rect 30288 3188 30340 3194
rect 30288 3130 30340 3136
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 30024 2650 30052 2994
rect 29460 2644 29512 2650
rect 29460 2586 29512 2592
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 30484 2582 30512 4966
rect 30852 3641 30880 5102
rect 31036 4690 31064 5306
rect 31024 4684 31076 4690
rect 31024 4626 31076 4632
rect 31036 4282 31064 4626
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 31220 4214 31248 6190
rect 31312 5370 31340 6734
rect 31588 6254 31616 6938
rect 32128 6860 32180 6866
rect 32128 6802 32180 6808
rect 32140 6390 32168 6802
rect 32324 6458 32352 8230
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32128 6384 32180 6390
rect 32128 6326 32180 6332
rect 31576 6248 31628 6254
rect 31576 6190 31628 6196
rect 31852 6180 31904 6186
rect 31852 6122 31904 6128
rect 31576 5704 31628 5710
rect 31576 5646 31628 5652
rect 31300 5364 31352 5370
rect 31300 5306 31352 5312
rect 31588 5166 31616 5646
rect 31864 5234 31892 6122
rect 31852 5228 31904 5234
rect 31852 5170 31904 5176
rect 31576 5160 31628 5166
rect 31576 5102 31628 5108
rect 31484 4480 31536 4486
rect 31484 4422 31536 4428
rect 31208 4208 31260 4214
rect 31208 4150 31260 4156
rect 31220 3670 31248 4150
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 31208 3664 31260 3670
rect 30838 3632 30894 3641
rect 31208 3606 31260 3612
rect 30838 3567 30894 3576
rect 31220 2990 31248 3606
rect 31404 3380 31432 4082
rect 31496 4010 31524 4422
rect 31484 4004 31536 4010
rect 31484 3946 31536 3952
rect 31496 3738 31524 3946
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31484 3392 31536 3398
rect 31404 3352 31484 3380
rect 31484 3334 31536 3340
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31220 2582 31248 2926
rect 31496 2650 31524 3334
rect 31588 3058 31616 5102
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 31852 3596 31904 3602
rect 31852 3538 31904 3544
rect 31864 3194 31892 3538
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31576 3052 31628 3058
rect 31576 2994 31628 3000
rect 32140 2922 32168 4558
rect 32324 3194 32352 6394
rect 32416 5710 32444 9386
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 32600 8673 32628 9318
rect 33060 9178 33088 10406
rect 33508 10124 33560 10130
rect 33508 10066 33560 10072
rect 33520 9761 33548 10066
rect 33506 9752 33562 9761
rect 33506 9687 33508 9696
rect 33560 9687 33562 9696
rect 33508 9658 33560 9664
rect 33520 9627 33548 9658
rect 33600 9580 33652 9586
rect 33600 9522 33652 9528
rect 33232 9376 33284 9382
rect 33232 9318 33284 9324
rect 33508 9376 33560 9382
rect 33508 9318 33560 9324
rect 33048 9172 33100 9178
rect 33048 9114 33100 9120
rect 32680 9036 32732 9042
rect 32680 8978 32732 8984
rect 32586 8664 32642 8673
rect 32692 8634 32720 8978
rect 33244 8974 33272 9318
rect 33324 9172 33376 9178
rect 33324 9114 33376 9120
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 33232 8968 33284 8974
rect 33232 8910 33284 8916
rect 32586 8599 32642 8608
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32588 8356 32640 8362
rect 32588 8298 32640 8304
rect 32600 8022 32628 8298
rect 32588 8016 32640 8022
rect 32588 7958 32640 7964
rect 32496 7880 32548 7886
rect 32496 7822 32548 7828
rect 32508 7546 32536 7822
rect 32496 7540 32548 7546
rect 32496 7482 32548 7488
rect 32496 7200 32548 7206
rect 32600 7188 32628 7958
rect 32548 7160 32628 7188
rect 32496 7142 32548 7148
rect 32508 5846 32536 7142
rect 32692 6866 32720 8570
rect 32680 6860 32732 6866
rect 32680 6802 32732 6808
rect 32692 6458 32720 6802
rect 32680 6452 32732 6458
rect 32680 6394 32732 6400
rect 32496 5840 32548 5846
rect 32496 5782 32548 5788
rect 32404 5704 32456 5710
rect 32404 5646 32456 5652
rect 32508 5098 32536 5782
rect 32876 5778 32904 8910
rect 33336 8838 33364 9114
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33324 8832 33376 8838
rect 33324 8774 33376 8780
rect 33152 8430 33180 8774
rect 33336 8498 33364 8774
rect 33324 8492 33376 8498
rect 33324 8434 33376 8440
rect 33140 8424 33192 8430
rect 33140 8366 33192 8372
rect 33520 8090 33548 9318
rect 33612 8945 33640 9522
rect 33598 8936 33654 8945
rect 33598 8871 33654 8880
rect 33704 8401 33732 10406
rect 34704 10124 34756 10130
rect 34704 10066 34756 10072
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34716 9382 34744 10066
rect 34704 9376 34756 9382
rect 34704 9318 34756 9324
rect 34716 9178 34744 9318
rect 34704 9172 34756 9178
rect 34704 9114 34756 9120
rect 34152 9104 34204 9110
rect 34152 9046 34204 9052
rect 33968 8968 34020 8974
rect 33968 8910 34020 8916
rect 34060 8968 34112 8974
rect 34060 8910 34112 8916
rect 33690 8392 33746 8401
rect 33690 8327 33746 8336
rect 33980 8090 34008 8910
rect 34072 8498 34100 8910
rect 34060 8492 34112 8498
rect 34060 8434 34112 8440
rect 34164 8276 34192 9046
rect 34716 8945 34744 9114
rect 34702 8936 34758 8945
rect 34702 8871 34758 8880
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34992 8498 35020 8774
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34244 8288 34296 8294
rect 34164 8248 34244 8276
rect 34244 8230 34296 8236
rect 34520 8288 34572 8294
rect 34520 8230 34572 8236
rect 33508 8084 33560 8090
rect 33508 8026 33560 8032
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 33048 8016 33100 8022
rect 33048 7958 33100 7964
rect 33060 7750 33088 7958
rect 33048 7744 33100 7750
rect 33048 7686 33100 7692
rect 33060 7546 33088 7686
rect 33048 7540 33100 7546
rect 33048 7482 33100 7488
rect 33060 7274 33088 7482
rect 33520 7410 33548 8026
rect 34256 8022 34284 8230
rect 34532 8129 34560 8230
rect 34518 8120 34574 8129
rect 34428 8084 34480 8090
rect 34518 8055 34574 8064
rect 34428 8026 34480 8032
rect 34244 8016 34296 8022
rect 34058 7984 34114 7993
rect 34440 7993 34468 8026
rect 34244 7958 34296 7964
rect 34426 7984 34482 7993
rect 34058 7919 34114 7928
rect 34152 7948 34204 7954
rect 33508 7404 33560 7410
rect 33508 7346 33560 7352
rect 33048 7268 33100 7274
rect 33048 7210 33100 7216
rect 33784 6792 33836 6798
rect 33784 6734 33836 6740
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33336 6322 33364 6598
rect 33324 6316 33376 6322
rect 33324 6258 33376 6264
rect 33692 6316 33744 6322
rect 33692 6258 33744 6264
rect 33048 6112 33100 6118
rect 33048 6054 33100 6060
rect 33060 5914 33088 6054
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 33140 5840 33192 5846
rect 33140 5782 33192 5788
rect 32864 5772 32916 5778
rect 32864 5714 32916 5720
rect 33048 5568 33100 5574
rect 33152 5556 33180 5782
rect 33100 5528 33180 5556
rect 33048 5510 33100 5516
rect 32586 5264 32642 5273
rect 32586 5199 32642 5208
rect 32956 5228 33008 5234
rect 32496 5092 32548 5098
rect 32496 5034 32548 5040
rect 32600 4826 32628 5199
rect 32956 5170 33008 5176
rect 32968 4826 32996 5170
rect 32588 4820 32640 4826
rect 32588 4762 32640 4768
rect 32956 4820 33008 4826
rect 32956 4762 33008 4768
rect 32600 4078 32628 4762
rect 33600 4208 33652 4214
rect 33600 4150 33652 4156
rect 33704 4154 33732 6258
rect 33796 5914 33824 6734
rect 33784 5908 33836 5914
rect 33784 5850 33836 5856
rect 33876 5704 33928 5710
rect 33876 5646 33928 5652
rect 33888 5370 33916 5646
rect 33876 5364 33928 5370
rect 33876 5306 33928 5312
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 33324 4004 33376 4010
rect 33324 3946 33376 3952
rect 33140 3936 33192 3942
rect 33140 3878 33192 3884
rect 32312 3188 32364 3194
rect 32312 3130 32364 3136
rect 32324 2990 32352 3130
rect 33152 3058 33180 3878
rect 33336 3602 33364 3946
rect 33612 3670 33640 4150
rect 33704 4126 33824 4154
rect 33600 3664 33652 3670
rect 33600 3606 33652 3612
rect 33324 3596 33376 3602
rect 33324 3538 33376 3544
rect 33336 3194 33364 3538
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 33612 3126 33640 3606
rect 33796 3126 33824 4126
rect 33980 3942 34008 4558
rect 33968 3936 34020 3942
rect 33968 3878 34020 3884
rect 33600 3120 33652 3126
rect 33600 3062 33652 3068
rect 33784 3120 33836 3126
rect 33784 3062 33836 3068
rect 33140 3052 33192 3058
rect 33140 2994 33192 3000
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 32864 2984 32916 2990
rect 32864 2926 32916 2932
rect 32128 2916 32180 2922
rect 32128 2858 32180 2864
rect 31484 2644 31536 2650
rect 31484 2586 31536 2592
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 31208 2576 31260 2582
rect 31208 2518 31260 2524
rect 31220 2378 31248 2518
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 31208 2372 31260 2378
rect 31208 2314 31260 2320
rect 29366 82 29422 480
rect 29104 54 29422 82
rect 26974 0 27030 54
rect 29366 0 29422 54
rect 31666 82 31722 480
rect 31772 82 31800 2382
rect 32876 2378 32904 2926
rect 34072 2650 34100 7919
rect 34426 7919 34482 7928
rect 34152 7890 34204 7896
rect 34164 7546 34192 7890
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34152 7540 34204 7546
rect 34152 7482 34204 7488
rect 34624 7478 34652 8298
rect 34704 8016 34756 8022
rect 34704 7958 34756 7964
rect 34612 7472 34664 7478
rect 34612 7414 34664 7420
rect 34152 6996 34204 7002
rect 34152 6938 34204 6944
rect 34164 6458 34192 6938
rect 34624 6866 34652 7414
rect 34716 7206 34744 7958
rect 34980 7880 35032 7886
rect 34980 7822 35032 7828
rect 34992 7750 35020 7822
rect 34980 7744 35032 7750
rect 34980 7686 35032 7692
rect 34992 7274 35020 7686
rect 34980 7268 35032 7274
rect 34980 7210 35032 7216
rect 34704 7200 34756 7206
rect 34704 7142 34756 7148
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34716 7002 34744 7142
rect 34704 6996 34756 7002
rect 34704 6938 34756 6944
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34808 6662 34836 7142
rect 34796 6656 34848 6662
rect 34796 6598 34848 6604
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34152 6452 34204 6458
rect 34152 6394 34204 6400
rect 34164 5914 34192 6394
rect 34808 5914 34836 6598
rect 35072 6384 35124 6390
rect 35072 6326 35124 6332
rect 34152 5908 34204 5914
rect 34152 5850 34204 5856
rect 34796 5908 34848 5914
rect 34796 5850 34848 5856
rect 34164 5234 34192 5850
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34704 5296 34756 5302
rect 34704 5238 34756 5244
rect 34152 5228 34204 5234
rect 34152 5170 34204 5176
rect 34164 4758 34192 5170
rect 34152 4752 34204 4758
rect 34152 4694 34204 4700
rect 34164 4214 34192 4694
rect 34612 4480 34664 4486
rect 34612 4422 34664 4428
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 34624 4282 34652 4422
rect 34612 4276 34664 4282
rect 34612 4218 34664 4224
rect 34152 4208 34204 4214
rect 34152 4150 34204 4156
rect 34624 3942 34652 4218
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 34716 3194 34744 5238
rect 35084 5234 35112 6326
rect 35176 5409 35204 10406
rect 35452 10266 35480 10746
rect 35440 10260 35492 10266
rect 35440 10202 35492 10208
rect 35348 9988 35400 9994
rect 35348 9930 35400 9936
rect 35360 8974 35388 9930
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 35452 6934 35480 9862
rect 35544 9722 35572 14991
rect 35714 14240 35770 14249
rect 35714 14175 35770 14184
rect 35622 11520 35678 11529
rect 35622 11455 35678 11464
rect 35636 11354 35664 11455
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 35622 10840 35678 10849
rect 35622 10775 35678 10784
rect 35636 10742 35664 10775
rect 35624 10736 35676 10742
rect 35624 10678 35676 10684
rect 35728 10266 35756 14175
rect 39578 13800 39634 13809
rect 39578 13735 39634 13744
rect 39592 12986 39620 13735
rect 39580 12980 39632 12986
rect 39580 12922 39632 12928
rect 36726 12336 36782 12345
rect 36726 12271 36782 12280
rect 36176 11008 36228 11014
rect 36176 10950 36228 10956
rect 36082 10704 36138 10713
rect 36082 10639 36138 10648
rect 35716 10260 35768 10266
rect 35716 10202 35768 10208
rect 36096 10130 36124 10639
rect 35900 10124 35952 10130
rect 35900 10066 35952 10072
rect 36084 10124 36136 10130
rect 36084 10066 36136 10072
rect 35912 9722 35940 10066
rect 35532 9716 35584 9722
rect 35532 9658 35584 9664
rect 35900 9716 35952 9722
rect 35900 9658 35952 9664
rect 35912 9625 35940 9658
rect 35898 9616 35954 9625
rect 35532 9580 35584 9586
rect 35898 9551 35954 9560
rect 35532 9522 35584 9528
rect 35440 6928 35492 6934
rect 35440 6870 35492 6876
rect 35256 6792 35308 6798
rect 35256 6734 35308 6740
rect 35268 5574 35296 6734
rect 35452 6322 35480 6870
rect 35440 6316 35492 6322
rect 35440 6258 35492 6264
rect 35256 5568 35308 5574
rect 35256 5510 35308 5516
rect 35162 5400 35218 5409
rect 35162 5335 35218 5344
rect 35072 5228 35124 5234
rect 34992 5188 35072 5216
rect 34992 4826 35020 5188
rect 35072 5170 35124 5176
rect 35072 5092 35124 5098
rect 35072 5034 35124 5040
rect 35084 4826 35112 5034
rect 34980 4820 35032 4826
rect 34980 4762 35032 4768
rect 35072 4820 35124 4826
rect 35072 4762 35124 4768
rect 34888 4752 34940 4758
rect 34888 4694 34940 4700
rect 34900 4282 34928 4694
rect 35268 4690 35296 5510
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 35256 4684 35308 4690
rect 35256 4626 35308 4632
rect 35164 4616 35216 4622
rect 35164 4558 35216 4564
rect 34888 4276 34940 4282
rect 34888 4218 34940 4224
rect 35176 3534 35204 4558
rect 35360 4214 35388 5170
rect 35440 4752 35492 4758
rect 35440 4694 35492 4700
rect 35452 4282 35480 4694
rect 35440 4276 35492 4282
rect 35440 4218 35492 4224
rect 35348 4208 35400 4214
rect 35348 4150 35400 4156
rect 35440 4004 35492 4010
rect 35440 3946 35492 3952
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 34716 2854 34744 3130
rect 35452 3058 35480 3946
rect 34980 3052 35032 3058
rect 34980 2994 35032 3000
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 34704 2848 34756 2854
rect 34704 2790 34756 2796
rect 34992 2650 35020 2994
rect 34060 2644 34112 2650
rect 34060 2586 34112 2592
rect 34980 2644 35032 2650
rect 34980 2586 35032 2592
rect 32864 2372 32916 2378
rect 32864 2314 32916 2320
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 33782 1184 33838 1193
rect 33782 1119 33838 1128
rect 31666 54 31800 82
rect 33796 82 33824 1119
rect 35544 1057 35572 9522
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35636 8634 35664 9046
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35900 8560 35952 8566
rect 35900 8502 35952 8508
rect 35912 8090 35940 8502
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35636 7274 35664 7822
rect 35912 7410 35940 8026
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 35624 7268 35676 7274
rect 35624 7210 35676 7216
rect 35636 3466 35664 7210
rect 35992 6928 36044 6934
rect 35992 6870 36044 6876
rect 36004 6458 36032 6870
rect 35992 6452 36044 6458
rect 35992 6394 36044 6400
rect 35992 6180 36044 6186
rect 35992 6122 36044 6128
rect 35900 6112 35952 6118
rect 35900 6054 35952 6060
rect 35912 5846 35940 6054
rect 35900 5840 35952 5846
rect 35900 5782 35952 5788
rect 35912 5370 35940 5782
rect 36004 5710 36032 6122
rect 35992 5704 36044 5710
rect 35992 5646 36044 5652
rect 35900 5364 35952 5370
rect 35900 5306 35952 5312
rect 36004 5234 36032 5646
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 35808 4684 35860 4690
rect 35808 4626 35860 4632
rect 35624 3460 35676 3466
rect 35624 3402 35676 3408
rect 35636 2650 35664 3402
rect 35820 3058 35848 4626
rect 36004 4282 36032 5170
rect 36188 5098 36216 10950
rect 36544 9988 36596 9994
rect 36544 9930 36596 9936
rect 36452 9512 36504 9518
rect 36452 9454 36504 9460
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36280 8634 36308 8910
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 36464 8537 36492 9454
rect 36450 8528 36506 8537
rect 36450 8463 36506 8472
rect 36452 7948 36504 7954
rect 36452 7890 36504 7896
rect 36360 7812 36412 7818
rect 36360 7754 36412 7760
rect 36372 7410 36400 7754
rect 36464 7546 36492 7890
rect 36452 7540 36504 7546
rect 36452 7482 36504 7488
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 36372 6934 36400 7346
rect 36360 6928 36412 6934
rect 36360 6870 36412 6876
rect 36556 6186 36584 9930
rect 36634 8800 36690 8809
rect 36634 8735 36690 8744
rect 36648 8634 36676 8735
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 36634 7984 36690 7993
rect 36634 7919 36690 7928
rect 36648 7818 36676 7919
rect 36636 7812 36688 7818
rect 36636 7754 36688 7760
rect 36544 6180 36596 6186
rect 36544 6122 36596 6128
rect 36556 5914 36584 6122
rect 36544 5908 36596 5914
rect 36544 5850 36596 5856
rect 36636 5296 36688 5302
rect 36636 5238 36688 5244
rect 36648 5098 36676 5238
rect 36176 5092 36228 5098
rect 36176 5034 36228 5040
rect 36636 5092 36688 5098
rect 36636 5034 36688 5040
rect 36188 4826 36216 5034
rect 36176 4820 36228 4826
rect 36176 4762 36228 4768
rect 36740 4282 36768 12271
rect 37464 10056 37516 10062
rect 37464 9998 37516 10004
rect 37476 9382 37504 9998
rect 37646 9888 37702 9897
rect 37646 9823 37702 9832
rect 37660 9722 37688 9823
rect 37648 9716 37700 9722
rect 37648 9658 37700 9664
rect 37464 9376 37516 9382
rect 37464 9318 37516 9324
rect 36820 8900 36872 8906
rect 36820 8842 36872 8848
rect 36832 7750 36860 8842
rect 37372 8288 37424 8294
rect 37372 8230 37424 8236
rect 36820 7744 36872 7750
rect 36820 7686 36872 7692
rect 36832 7410 36860 7686
rect 36820 7404 36872 7410
rect 36820 7346 36872 7352
rect 35992 4276 36044 4282
rect 35992 4218 36044 4224
rect 36728 4276 36780 4282
rect 36728 4218 36780 4224
rect 37384 4078 37412 8230
rect 37476 6361 37504 9318
rect 38660 9172 38712 9178
rect 38660 9114 38712 9120
rect 38016 8424 38068 8430
rect 38016 8366 38068 8372
rect 38028 8022 38056 8366
rect 38016 8016 38068 8022
rect 38016 7958 38068 7964
rect 37462 6352 37518 6361
rect 37462 6287 37518 6296
rect 38028 4321 38056 7958
rect 38014 4312 38070 4321
rect 38014 4247 38070 4256
rect 36452 4072 36504 4078
rect 36452 4014 36504 4020
rect 37004 4072 37056 4078
rect 37004 4014 37056 4020
rect 37372 4072 37424 4078
rect 37372 4014 37424 4020
rect 36464 3913 36492 4014
rect 36450 3904 36506 3913
rect 36450 3839 36506 3848
rect 36268 3664 36320 3670
rect 36268 3606 36320 3612
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35912 3194 35940 3470
rect 36280 3194 36308 3606
rect 35900 3188 35952 3194
rect 35900 3130 35952 3136
rect 36268 3188 36320 3194
rect 36268 3130 36320 3136
rect 36910 3088 36966 3097
rect 35808 3052 35860 3058
rect 36910 3023 36966 3032
rect 35808 2994 35860 3000
rect 35624 2644 35676 2650
rect 35624 2586 35676 2592
rect 36924 2514 36952 3023
rect 37016 2990 37044 4014
rect 37004 2984 37056 2990
rect 37004 2926 37056 2932
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 35992 2304 36044 2310
rect 35992 2246 36044 2252
rect 35530 1048 35586 1057
rect 35530 983 35586 992
rect 34058 82 34114 480
rect 36004 377 36032 2246
rect 35990 368 36046 377
rect 35990 303 36046 312
rect 33796 54 34114 82
rect 36096 82 36124 2314
rect 38672 1329 38700 9114
rect 39578 6624 39634 6633
rect 39408 6582 39578 6610
rect 39408 5681 39436 6582
rect 39578 6559 39634 6568
rect 39394 5672 39450 5681
rect 39394 5607 39450 5616
rect 38474 1320 38530 1329
rect 38474 1255 38530 1264
rect 38658 1320 38714 1329
rect 38658 1255 38714 1264
rect 36358 82 36414 480
rect 36096 54 36414 82
rect 38488 82 38516 1255
rect 38750 82 38806 480
rect 38488 54 38806 82
rect 31666 0 31722 54
rect 34058 0 34114 54
rect 36358 0 36414 54
rect 38750 0 38806 54
<< via2 >>
rect 938 15000 994 15056
rect 110 13744 166 13800
rect 110 11056 166 11112
rect 1030 14184 1086 14240
rect 1490 12280 1546 12336
rect 18 10240 74 10296
rect 110 2216 166 2272
rect 2318 9152 2374 9208
rect 2686 9324 2688 9344
rect 2688 9324 2740 9344
rect 2740 9324 2742 9344
rect 2686 9288 2742 9324
rect 2318 6976 2374 7032
rect 2962 9968 3018 10024
rect 2962 7928 3018 7984
rect 3330 9560 3386 9616
rect 3882 10104 3938 10160
rect 3882 8744 3938 8800
rect 3238 5752 3294 5808
rect 4526 11464 4582 11520
rect 4158 6976 4214 7032
rect 4526 4528 4582 4584
rect 3606 3576 3662 3632
rect 1490 992 1546 1048
rect 1122 40 1178 96
rect 5446 11736 5502 11792
rect 5262 10648 5318 10704
rect 6090 11212 6146 11248
rect 6090 11192 6092 11212
rect 6092 11192 6144 11212
rect 6144 11192 6146 11212
rect 5538 9172 5594 9208
rect 5538 9152 5540 9172
rect 5540 9152 5592 9172
rect 5592 9152 5594 9172
rect 5814 8064 5870 8120
rect 5998 8472 6054 8528
rect 5722 3984 5778 4040
rect 5446 3032 5502 3088
rect 5262 1808 5318 1864
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 6182 7112 6238 7168
rect 6642 6160 6698 6216
rect 7378 10104 7434 10160
rect 7378 7792 7434 7848
rect 7378 7112 7434 7168
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 7562 10512 7618 10568
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 8666 6432 8722 6488
rect 9126 9968 9182 10024
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 9218 4120 9274 4176
rect 9126 3712 9182 3768
rect 9402 8880 9458 8936
rect 10230 9560 10286 9616
rect 9402 6296 9458 6352
rect 9586 5208 9642 5264
rect 9586 4528 9642 4584
rect 9770 4120 9826 4176
rect 11702 9696 11758 9752
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 12254 11464 12310 11520
rect 12070 11328 12126 11384
rect 11242 6704 11298 6760
rect 10506 5480 10562 5536
rect 10598 5072 10654 5128
rect 10506 3984 10562 4040
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 6918 1536 6974 1592
rect 5998 1128 6054 1184
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 12898 8744 12954 8800
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 12714 3032 12770 3088
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14186 6160 14242 6216
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14738 7928 14794 7984
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14002 3576 14058 3632
rect 15474 6432 15530 6488
rect 15658 5480 15714 5536
rect 15474 5208 15530 5264
rect 14738 4256 14794 4312
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 12254 1264 12310 1320
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 14830 1808 14886 1864
rect 14094 1536 14150 1592
rect 15750 4120 15806 4176
rect 15382 3848 15438 3904
rect 16026 3712 16082 3768
rect 17314 11736 17370 11792
rect 18510 11212 18566 11248
rect 18510 11192 18512 11212
rect 18512 11192 18564 11212
rect 18564 11192 18566 11212
rect 18326 10648 18382 10704
rect 18510 10648 18566 10704
rect 17958 8472 18014 8528
rect 16578 2624 16634 2680
rect 17498 4004 17554 4040
rect 17498 3984 17500 4004
rect 17500 3984 17552 4004
rect 17552 3984 17554 4004
rect 18234 5072 18290 5128
rect 19522 11056 19578 11112
rect 19522 10104 19578 10160
rect 19338 9832 19394 9888
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 19154 4120 19210 4176
rect 18234 3984 18290 4040
rect 18970 3596 19026 3632
rect 18970 3576 18972 3596
rect 18972 3576 19024 3596
rect 19024 3576 19026 3596
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 21638 8608 21694 8664
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 19522 4256 19578 4312
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20718 3984 20774 4040
rect 21086 3984 21142 4040
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 21270 2624 21326 2680
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 22374 10512 22430 10568
rect 22098 6296 22154 6352
rect 22742 8472 22798 8528
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 23938 9560 23994 9616
rect 23386 8472 23442 8528
rect 23386 6160 23442 6216
rect 23938 7792 23994 7848
rect 24398 3576 24454 3632
rect 23294 2896 23350 2952
rect 26238 10920 26294 10976
rect 25502 10648 25558 10704
rect 24674 8472 24730 8528
rect 25502 9696 25558 9752
rect 25042 9424 25098 9480
rect 27894 10512 27950 10568
rect 28078 10512 28134 10568
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 26974 9968 27030 10024
rect 26606 9016 26662 9072
rect 26606 6704 26662 6760
rect 26974 8880 27030 8936
rect 24582 3984 24638 4040
rect 25410 3848 25466 3904
rect 26882 6296 26938 6352
rect 26974 5616 27030 5672
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 28262 8472 28318 8528
rect 28446 7928 28502 7984
rect 28262 7384 28318 7440
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 28078 4528 28134 4584
rect 28078 3848 28134 3904
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 28906 6160 28962 6216
rect 28722 4528 28778 4584
rect 35530 15000 35586 15056
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 33046 11056 33102 11112
rect 34150 10920 34206 10976
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 35346 10512 35402 10568
rect 29826 9560 29882 9616
rect 28814 3032 28870 3088
rect 26606 1400 26662 1456
rect 26514 1128 26570 1184
rect 27250 312 27306 368
rect 30378 6840 30434 6896
rect 30838 3576 30894 3632
rect 33506 9716 33562 9752
rect 33506 9696 33508 9716
rect 33508 9696 33560 9716
rect 33560 9696 33562 9716
rect 32586 8608 32642 8664
rect 33598 8880 33654 8936
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 33690 8336 33746 8392
rect 34702 8880 34758 8936
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 34518 8064 34574 8120
rect 34058 7928 34114 7984
rect 32586 5208 32642 5264
rect 34426 7928 34482 7984
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 35714 14184 35770 14240
rect 35622 11464 35678 11520
rect 35622 10784 35678 10840
rect 39578 13744 39634 13800
rect 36726 12280 36782 12336
rect 36082 10648 36138 10704
rect 35898 9560 35954 9616
rect 35162 5344 35218 5400
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 33782 1128 33838 1184
rect 36450 8472 36506 8528
rect 36634 8744 36690 8800
rect 36634 7928 36690 7984
rect 37646 9832 37702 9888
rect 37462 6296 37518 6352
rect 38014 4256 38070 4312
rect 36450 3848 36506 3904
rect 36910 3032 36966 3088
rect 35530 992 35586 1048
rect 35990 312 36046 368
rect 39578 6568 39634 6624
rect 39394 5616 39450 5672
rect 38474 1264 38530 1320
rect 38658 1264 38714 1320
<< metal3 >>
rect 0 15512 480 15632
rect 39520 15512 40000 15632
rect 62 15058 122 15512
rect 933 15058 999 15061
rect 62 15056 999 15058
rect 62 15000 938 15056
rect 994 15000 999 15056
rect 62 14998 999 15000
rect 933 14995 999 14998
rect 35525 15058 35591 15061
rect 39622 15058 39682 15512
rect 35525 15056 39682 15058
rect 35525 15000 35530 15056
rect 35586 15000 39682 15056
rect 35525 14998 39682 15000
rect 35525 14995 35591 14998
rect 0 14560 480 14680
rect 39520 14560 40000 14680
rect 62 14242 122 14560
rect 1025 14242 1091 14245
rect 62 14240 1091 14242
rect 62 14184 1030 14240
rect 1086 14184 1091 14240
rect 62 14182 1091 14184
rect 1025 14179 1091 14182
rect 35709 14242 35775 14245
rect 39622 14242 39682 14560
rect 35709 14240 39682 14242
rect 35709 14184 35714 14240
rect 35770 14184 39682 14240
rect 35709 14182 39682 14184
rect 35709 14179 35775 14182
rect 0 13800 480 13864
rect 39520 13802 40000 13864
rect 0 13744 110 13800
rect 166 13744 480 13800
rect 39492 13800 40000 13802
rect 39492 13744 39578 13800
rect 39634 13744 40000 13800
rect 105 13742 252 13744
rect 39492 13742 39639 13744
rect 105 13739 171 13742
rect 39573 13739 39639 13742
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 0 12792 480 12912
rect 39520 12792 40000 12912
rect 62 12338 122 12792
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 1485 12338 1551 12341
rect 62 12336 1551 12338
rect 62 12280 1490 12336
rect 1546 12280 1551 12336
rect 62 12278 1551 12280
rect 1485 12275 1551 12278
rect 36721 12338 36787 12341
rect 39622 12338 39682 12792
rect 36721 12336 39682 12338
rect 36721 12280 36726 12336
rect 36782 12280 39682 12336
rect 36721 12278 39682 12280
rect 36721 12275 36787 12278
rect 0 11976 480 12096
rect 7610 12000 7930 12001
rect 62 11522 122 11976
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12096
rect 34277 11935 34597 11936
rect 5441 11794 5507 11797
rect 17309 11794 17375 11797
rect 5441 11792 17375 11794
rect 5441 11736 5446 11792
rect 5502 11736 17314 11792
rect 17370 11736 17375 11792
rect 5441 11734 17375 11736
rect 5441 11731 5507 11734
rect 17309 11731 17375 11734
rect 4521 11522 4587 11525
rect 62 11520 4587 11522
rect 62 11464 4526 11520
rect 4582 11464 4587 11520
rect 62 11462 4587 11464
rect 4521 11459 4587 11462
rect 12249 11522 12315 11525
rect 12382 11522 12388 11524
rect 12249 11520 12388 11522
rect 12249 11464 12254 11520
rect 12310 11464 12388 11520
rect 12249 11462 12388 11464
rect 12249 11459 12315 11462
rect 12382 11460 12388 11462
rect 12452 11460 12458 11524
rect 35617 11522 35683 11525
rect 39622 11522 39682 11976
rect 35617 11520 39682 11522
rect 35617 11464 35622 11520
rect 35678 11464 39682 11520
rect 35617 11462 39682 11464
rect 35617 11459 35683 11462
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 12065 11386 12131 11389
rect 12750 11386 12756 11388
rect 12065 11384 12756 11386
rect 12065 11328 12070 11384
rect 12126 11328 12756 11384
rect 12065 11326 12756 11328
rect 12065 11323 12131 11326
rect 12750 11324 12756 11326
rect 12820 11324 12826 11388
rect 6085 11250 6151 11253
rect 18505 11250 18571 11253
rect 6085 11248 18571 11250
rect 6085 11192 6090 11248
rect 6146 11192 18510 11248
rect 18566 11192 18571 11248
rect 6085 11190 18571 11192
rect 6085 11187 6151 11190
rect 18505 11187 18571 11190
rect 0 11112 480 11144
rect 0 11056 110 11112
rect 166 11056 480 11112
rect 0 11024 480 11056
rect 19517 11114 19583 11117
rect 33041 11114 33107 11117
rect 19517 11112 33107 11114
rect 19517 11056 19522 11112
rect 19578 11056 33046 11112
rect 33102 11056 33107 11112
rect 19517 11054 33107 11056
rect 19517 11051 19583 11054
rect 33041 11051 33107 11054
rect 39520 11024 40000 11144
rect 26233 10978 26299 10981
rect 34145 10978 34211 10981
rect 26233 10976 34211 10978
rect 26233 10920 26238 10976
rect 26294 10920 34150 10976
rect 34206 10920 34211 10976
rect 26233 10918 34211 10920
rect 26233 10915 26299 10918
rect 34145 10915 34211 10918
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 35617 10842 35683 10845
rect 39622 10842 39682 11024
rect 35617 10840 39682 10842
rect 35617 10784 35622 10840
rect 35678 10784 39682 10840
rect 35617 10782 39682 10784
rect 35617 10779 35683 10782
rect 5257 10706 5323 10709
rect 18321 10706 18387 10709
rect 5257 10704 18387 10706
rect 5257 10648 5262 10704
rect 5318 10648 18326 10704
rect 18382 10648 18387 10704
rect 5257 10646 18387 10648
rect 5257 10643 5323 10646
rect 18321 10643 18387 10646
rect 18505 10706 18571 10709
rect 25497 10706 25563 10709
rect 36077 10706 36143 10709
rect 18505 10704 25563 10706
rect 18505 10648 18510 10704
rect 18566 10648 25502 10704
rect 25558 10648 25563 10704
rect 18505 10646 25563 10648
rect 18505 10643 18571 10646
rect 25497 10643 25563 10646
rect 27846 10704 36143 10706
rect 27846 10648 36082 10704
rect 36138 10648 36143 10704
rect 27846 10646 36143 10648
rect 27846 10573 27906 10646
rect 36077 10643 36143 10646
rect 7557 10570 7623 10573
rect 22369 10570 22435 10573
rect 7557 10568 22435 10570
rect 7557 10512 7562 10568
rect 7618 10512 22374 10568
rect 22430 10512 22435 10568
rect 7557 10510 22435 10512
rect 7557 10507 7623 10510
rect 22369 10507 22435 10510
rect 23422 10508 23428 10572
rect 23492 10570 23498 10572
rect 27846 10570 27955 10573
rect 23492 10568 27955 10570
rect 23492 10512 27894 10568
rect 27950 10512 27955 10568
rect 23492 10510 27955 10512
rect 23492 10508 23498 10510
rect 27889 10507 27955 10510
rect 28073 10570 28139 10573
rect 35341 10570 35407 10573
rect 28073 10568 35407 10570
rect 28073 10512 28078 10568
rect 28134 10512 35346 10568
rect 35402 10512 35407 10568
rect 28073 10510 35407 10512
rect 28073 10507 28139 10510
rect 35341 10507 35407 10510
rect 14277 10368 14597 10369
rect 0 10296 480 10328
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 0 10240 18 10296
rect 74 10240 480 10296
rect 0 10208 480 10240
rect 39520 10208 40000 10328
rect 3877 10162 3943 10165
rect 7373 10162 7439 10165
rect 19517 10162 19583 10165
rect 3877 10160 3986 10162
rect 3877 10104 3882 10160
rect 3938 10104 3986 10160
rect 3877 10099 3986 10104
rect 7373 10160 19583 10162
rect 7373 10104 7378 10160
rect 7434 10104 19522 10160
rect 19578 10104 19583 10160
rect 7373 10102 19583 10104
rect 7373 10099 7439 10102
rect 19517 10099 19583 10102
rect 2957 10026 3023 10029
rect 3926 10026 3986 10099
rect 9121 10026 9187 10029
rect 26969 10026 27035 10029
rect 2957 10024 8954 10026
rect 2957 9968 2962 10024
rect 3018 9968 8954 10024
rect 2957 9966 8954 9968
rect 2957 9963 3023 9966
rect 8894 9890 8954 9966
rect 9121 10024 27035 10026
rect 9121 9968 9126 10024
rect 9182 9968 26974 10024
rect 27030 9968 27035 10024
rect 9121 9966 27035 9968
rect 9121 9963 9187 9966
rect 26969 9963 27035 9966
rect 19333 9890 19399 9893
rect 8894 9888 19399 9890
rect 8894 9832 19338 9888
rect 19394 9832 19399 9888
rect 8894 9830 19399 9832
rect 19333 9827 19399 9830
rect 37641 9890 37707 9893
rect 39622 9890 39682 10208
rect 37641 9888 39682 9890
rect 37641 9832 37646 9888
rect 37702 9832 39682 9888
rect 37641 9830 39682 9832
rect 37641 9827 37707 9830
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 9622 9692 9628 9756
rect 9692 9754 9698 9756
rect 11697 9754 11763 9757
rect 9692 9752 11763 9754
rect 9692 9696 11702 9752
rect 11758 9696 11763 9752
rect 9692 9694 11763 9696
rect 9692 9692 9698 9694
rect 11697 9691 11763 9694
rect 25497 9754 25563 9757
rect 33501 9754 33567 9757
rect 25497 9752 33567 9754
rect 25497 9696 25502 9752
rect 25558 9696 33506 9752
rect 33562 9696 33567 9752
rect 25497 9694 33567 9696
rect 25497 9691 25563 9694
rect 33501 9691 33567 9694
rect 3325 9620 3391 9621
rect 3325 9618 3372 9620
rect 3244 9616 3372 9618
rect 3436 9618 3442 9620
rect 10225 9618 10291 9621
rect 3436 9616 10291 9618
rect 3244 9560 3330 9616
rect 3436 9560 10230 9616
rect 10286 9560 10291 9616
rect 3244 9558 3372 9560
rect 3325 9556 3372 9558
rect 3436 9558 10291 9560
rect 3436 9556 3442 9558
rect 3325 9555 3391 9556
rect 10225 9555 10291 9558
rect 23933 9618 23999 9621
rect 29821 9618 29887 9621
rect 35893 9618 35959 9621
rect 23933 9616 35959 9618
rect 23933 9560 23938 9616
rect 23994 9560 29826 9616
rect 29882 9560 35898 9616
rect 35954 9560 35959 9616
rect 23933 9558 35959 9560
rect 23933 9555 23999 9558
rect 29821 9555 29887 9558
rect 35893 9555 35959 9558
rect 25037 9482 25103 9485
rect 8894 9480 25103 9482
rect 8894 9424 25042 9480
rect 25098 9424 25103 9480
rect 8894 9422 25103 9424
rect 0 9256 480 9376
rect 2681 9346 2747 9349
rect 8894 9346 8954 9422
rect 25037 9419 25103 9422
rect 2681 9344 8954 9346
rect 2681 9288 2686 9344
rect 2742 9288 8954 9344
rect 2681 9286 8954 9288
rect 2681 9283 2747 9286
rect 14277 9280 14597 9281
rect 62 8802 122 9256
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9376
rect 27610 9215 27930 9216
rect 2313 9210 2379 9213
rect 5533 9210 5599 9213
rect 2313 9208 5599 9210
rect 2313 9152 2318 9208
rect 2374 9152 5538 9208
rect 5594 9152 5599 9208
rect 2313 9150 5599 9152
rect 2313 9147 2379 9150
rect 5533 9147 5599 9150
rect 26601 9074 26667 9077
rect 13770 9072 26667 9074
rect 13770 9016 26606 9072
rect 26662 9016 26667 9072
rect 13770 9014 26667 9016
rect 9397 8938 9463 8941
rect 13770 8938 13830 9014
rect 26601 9011 26667 9014
rect 26969 8938 27035 8941
rect 33593 8938 33659 8941
rect 34697 8938 34763 8941
rect 9397 8936 13830 8938
rect 9397 8880 9402 8936
rect 9458 8880 13830 8936
rect 9397 8878 13830 8880
rect 18600 8878 23490 8938
rect 9397 8875 9463 8878
rect 3877 8802 3943 8805
rect 62 8800 3943 8802
rect 62 8744 3882 8800
rect 3938 8744 3943 8800
rect 62 8742 3943 8744
rect 3877 8739 3943 8742
rect 12893 8802 12959 8805
rect 18600 8802 18660 8878
rect 12893 8800 18660 8802
rect 12893 8744 12898 8800
rect 12954 8744 18660 8800
rect 12893 8742 18660 8744
rect 23430 8802 23490 8878
rect 26969 8936 33659 8938
rect 26969 8880 26974 8936
rect 27030 8880 33598 8936
rect 33654 8880 33659 8936
rect 26969 8878 33659 8880
rect 26969 8875 27035 8878
rect 33593 8875 33659 8878
rect 33734 8936 34763 8938
rect 33734 8880 34702 8936
rect 34758 8880 34763 8936
rect 33734 8878 34763 8880
rect 33734 8802 33794 8878
rect 34697 8875 34763 8878
rect 23430 8742 33794 8802
rect 36629 8802 36695 8805
rect 39622 8802 39682 9256
rect 36629 8800 39682 8802
rect 36629 8744 36634 8800
rect 36690 8744 39682 8800
rect 36629 8742 39682 8744
rect 12893 8739 12959 8742
rect 36629 8739 36695 8742
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 21633 8666 21699 8669
rect 32581 8666 32647 8669
rect 21633 8664 32647 8666
rect 21633 8608 21638 8664
rect 21694 8608 32586 8664
rect 32642 8608 32647 8664
rect 21633 8606 32647 8608
rect 21633 8603 21699 8606
rect 32581 8603 32647 8606
rect 0 8440 480 8560
rect 5993 8530 6059 8533
rect 17953 8530 18019 8533
rect 22737 8530 22803 8533
rect 23381 8530 23447 8533
rect 24669 8530 24735 8533
rect 5993 8528 23260 8530
rect 5993 8472 5998 8528
rect 6054 8472 17958 8528
rect 18014 8472 22742 8528
rect 22798 8472 23260 8528
rect 5993 8470 23260 8472
rect 5993 8467 6059 8470
rect 17953 8467 18019 8470
rect 22737 8467 22803 8470
rect 62 8122 122 8440
rect 23200 8394 23260 8470
rect 23381 8528 24735 8530
rect 23381 8472 23386 8528
rect 23442 8472 24674 8528
rect 24730 8472 24735 8528
rect 23381 8470 24735 8472
rect 23381 8467 23447 8470
rect 24669 8467 24735 8470
rect 28257 8530 28323 8533
rect 36445 8530 36511 8533
rect 28257 8528 36511 8530
rect 28257 8472 28262 8528
rect 28318 8472 36450 8528
rect 36506 8472 36511 8528
rect 28257 8470 36511 8472
rect 28257 8467 28323 8470
rect 36445 8467 36511 8470
rect 39520 8440 40000 8560
rect 33685 8394 33751 8397
rect 23200 8392 34898 8394
rect 23200 8336 33690 8392
rect 33746 8336 34898 8392
rect 23200 8334 34898 8336
rect 33685 8331 33751 8334
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 5809 8122 5875 8125
rect 34513 8122 34579 8125
rect 62 8120 5875 8122
rect 62 8064 5814 8120
rect 5870 8064 5875 8120
rect 62 8062 5875 8064
rect 5809 8059 5875 8062
rect 28260 8120 34579 8122
rect 28260 8064 34518 8120
rect 34574 8064 34579 8120
rect 28260 8062 34579 8064
rect 2957 7986 3023 7989
rect 62 7984 3023 7986
rect 62 7928 2962 7984
rect 3018 7928 3023 7984
rect 62 7926 3023 7928
rect 62 7608 122 7926
rect 2957 7923 3023 7926
rect 14733 7986 14799 7989
rect 28260 7986 28320 8062
rect 34513 8059 34579 8062
rect 14733 7984 28320 7986
rect 14733 7928 14738 7984
rect 14794 7928 28320 7984
rect 14733 7926 28320 7928
rect 28441 7986 28507 7989
rect 34053 7986 34119 7989
rect 34421 7986 34487 7989
rect 28441 7984 34487 7986
rect 28441 7928 28446 7984
rect 28502 7928 34058 7984
rect 34114 7928 34426 7984
rect 34482 7928 34487 7984
rect 28441 7926 34487 7928
rect 14733 7923 14799 7926
rect 28441 7923 28507 7926
rect 34053 7923 34119 7926
rect 34421 7923 34487 7926
rect 7373 7850 7439 7853
rect 23933 7850 23999 7853
rect 7373 7848 23999 7850
rect 7373 7792 7378 7848
rect 7434 7792 23938 7848
rect 23994 7792 23999 7848
rect 7373 7790 23999 7792
rect 34838 7850 34898 8334
rect 36629 7986 36695 7989
rect 39622 7986 39682 8440
rect 36629 7984 39682 7986
rect 36629 7928 36634 7984
rect 36690 7928 39682 7984
rect 36629 7926 39682 7928
rect 36629 7923 36695 7926
rect 34838 7790 39682 7850
rect 7373 7787 7439 7790
rect 23933 7787 23999 7790
rect 7610 7648 7930 7649
rect 0 7488 480 7608
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 39622 7608 39682 7790
rect 34277 7583 34597 7584
rect 39520 7488 40000 7608
rect 23422 7380 23428 7444
rect 23492 7442 23498 7444
rect 28257 7442 28323 7445
rect 23492 7440 28323 7442
rect 23492 7384 28262 7440
rect 28318 7384 28323 7440
rect 23492 7382 28323 7384
rect 23492 7380 23498 7382
rect 28257 7379 28323 7382
rect 6177 7170 6243 7173
rect 7373 7170 7439 7173
rect 62 7168 7439 7170
rect 62 7112 6182 7168
rect 6238 7112 7378 7168
rect 7434 7112 7439 7168
rect 62 7110 7439 7112
rect 62 6656 122 7110
rect 6177 7107 6243 7110
rect 7373 7107 7439 7110
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 2313 7034 2379 7037
rect 4153 7034 4219 7037
rect 2313 7032 4219 7034
rect 2313 6976 2318 7032
rect 2374 6976 4158 7032
rect 4214 6976 4219 7032
rect 2313 6974 4219 6976
rect 2313 6971 2379 6974
rect 4110 6971 4219 6974
rect 4110 6898 4170 6971
rect 30373 6898 30439 6901
rect 4110 6896 30439 6898
rect 4110 6840 30378 6896
rect 30434 6840 30439 6896
rect 4110 6838 30439 6840
rect 30373 6835 30439 6838
rect 11237 6762 11303 6765
rect 26601 6762 26667 6765
rect 11237 6760 26667 6762
rect 11237 6704 11242 6760
rect 11298 6704 26606 6760
rect 26662 6704 26667 6760
rect 11237 6702 26667 6704
rect 11237 6699 11303 6702
rect 26601 6699 26667 6702
rect 0 6536 480 6656
rect 39520 6626 40000 6656
rect 39492 6624 40000 6626
rect 39492 6568 39578 6624
rect 39634 6568 40000 6624
rect 39492 6566 40000 6568
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 39520 6536 40000 6566
rect 34277 6495 34597 6496
rect 8661 6490 8727 6493
rect 15469 6490 15535 6493
rect 8661 6488 15535 6490
rect 8661 6432 8666 6488
rect 8722 6432 15474 6488
rect 15530 6432 15535 6488
rect 8661 6430 15535 6432
rect 8661 6427 8727 6430
rect 15469 6427 15535 6430
rect 9397 6354 9463 6357
rect 62 6352 9463 6354
rect 62 6296 9402 6352
rect 9458 6296 9463 6352
rect 62 6294 9463 6296
rect 62 5840 122 6294
rect 9397 6291 9463 6294
rect 22093 6354 22159 6357
rect 26877 6354 26943 6357
rect 22093 6352 26943 6354
rect 22093 6296 22098 6352
rect 22154 6296 26882 6352
rect 26938 6296 26943 6352
rect 22093 6294 26943 6296
rect 22093 6291 22159 6294
rect 26877 6291 26943 6294
rect 37457 6354 37523 6357
rect 37457 6352 39682 6354
rect 37457 6296 37462 6352
rect 37518 6296 39682 6352
rect 37457 6294 39682 6296
rect 37457 6291 37523 6294
rect 6637 6218 6703 6221
rect 14181 6218 14247 6221
rect 6637 6216 14247 6218
rect 6637 6160 6642 6216
rect 6698 6160 14186 6216
rect 14242 6160 14247 6216
rect 6637 6158 14247 6160
rect 6637 6155 6703 6158
rect 14181 6155 14247 6158
rect 23381 6218 23447 6221
rect 28901 6218 28967 6221
rect 23381 6216 28967 6218
rect 23381 6160 23386 6216
rect 23442 6160 28906 6216
rect 28962 6160 28967 6216
rect 23381 6158 28967 6160
rect 23381 6155 23447 6158
rect 28901 6155 28967 6158
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 39622 5840 39682 6294
rect 0 5720 480 5840
rect 3233 5810 3299 5813
rect 3366 5810 3372 5812
rect 3233 5808 3372 5810
rect 3233 5752 3238 5808
rect 3294 5752 3372 5808
rect 3233 5750 3372 5752
rect 3233 5747 3299 5750
rect 3366 5748 3372 5750
rect 3436 5748 3442 5812
rect 39520 5720 40000 5840
rect 26969 5674 27035 5677
rect 39389 5674 39455 5677
rect 26969 5672 39455 5674
rect 26969 5616 26974 5672
rect 27030 5616 39394 5672
rect 39450 5616 39455 5672
rect 26969 5614 39455 5616
rect 26969 5611 27035 5614
rect 39389 5611 39455 5614
rect 10501 5538 10567 5541
rect 15653 5538 15719 5541
rect 10501 5536 15719 5538
rect 10501 5480 10506 5536
rect 10562 5480 15658 5536
rect 15714 5480 15719 5536
rect 10501 5478 15719 5480
rect 10501 5475 10567 5478
rect 15653 5475 15719 5478
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 35157 5402 35223 5405
rect 35157 5400 39682 5402
rect 35157 5344 35162 5400
rect 35218 5344 39682 5400
rect 35157 5342 39682 5344
rect 35157 5339 35223 5342
rect 9581 5266 9647 5269
rect 62 5264 9647 5266
rect 62 5208 9586 5264
rect 9642 5208 9647 5264
rect 62 5206 9647 5208
rect 62 4888 122 5206
rect 9581 5203 9647 5206
rect 15469 5266 15535 5269
rect 32581 5266 32647 5269
rect 15469 5264 32647 5266
rect 15469 5208 15474 5264
rect 15530 5208 32586 5264
rect 32642 5208 32647 5264
rect 15469 5206 32647 5208
rect 15469 5203 15535 5206
rect 32581 5203 32647 5206
rect 10593 5130 10659 5133
rect 18229 5130 18295 5133
rect 10593 5128 18295 5130
rect 10593 5072 10598 5128
rect 10654 5072 18234 5128
rect 18290 5072 18295 5128
rect 10593 5070 18295 5072
rect 10593 5067 10659 5070
rect 18229 5067 18295 5070
rect 14277 4928 14597 4929
rect 0 4768 480 4888
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 39622 4888 39682 5342
rect 27610 4863 27930 4864
rect 39520 4768 40000 4888
rect 4521 4586 4587 4589
rect 62 4584 4587 4586
rect 62 4528 4526 4584
rect 4582 4528 4587 4584
rect 62 4526 4587 4528
rect 62 4072 122 4526
rect 4521 4523 4587 4526
rect 9581 4586 9647 4589
rect 28073 4586 28139 4589
rect 28717 4586 28783 4589
rect 9581 4584 28783 4586
rect 9581 4528 9586 4584
rect 9642 4528 28078 4584
rect 28134 4528 28722 4584
rect 28778 4528 28783 4584
rect 9581 4526 28783 4528
rect 9581 4523 9647 4526
rect 28073 4523 28139 4526
rect 28717 4523 28783 4526
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 14733 4314 14799 4317
rect 19517 4314 19583 4317
rect 14733 4312 19583 4314
rect 14733 4256 14738 4312
rect 14794 4256 19522 4312
rect 19578 4256 19583 4312
rect 14733 4254 19583 4256
rect 14733 4251 14799 4254
rect 19517 4251 19583 4254
rect 38009 4314 38075 4317
rect 39614 4314 39620 4316
rect 38009 4312 39620 4314
rect 38009 4256 38014 4312
rect 38070 4256 39620 4312
rect 38009 4254 39620 4256
rect 38009 4251 38075 4254
rect 39614 4252 39620 4254
rect 39684 4252 39690 4316
rect 9213 4178 9279 4181
rect 9765 4178 9831 4181
rect 9213 4176 9831 4178
rect 9213 4120 9218 4176
rect 9274 4120 9770 4176
rect 9826 4120 9831 4176
rect 9213 4118 9831 4120
rect 9213 4115 9279 4118
rect 9765 4115 9831 4118
rect 15745 4178 15811 4181
rect 19149 4178 19215 4181
rect 15745 4176 19215 4178
rect 15745 4120 15750 4176
rect 15806 4120 19154 4176
rect 19210 4120 19215 4176
rect 15745 4118 19215 4120
rect 15745 4115 15811 4118
rect 19149 4115 19215 4118
rect 0 3952 480 4072
rect 5717 4042 5783 4045
rect 10501 4042 10567 4045
rect 5717 4040 10567 4042
rect 5717 3984 5722 4040
rect 5778 3984 10506 4040
rect 10562 3984 10567 4040
rect 5717 3982 10567 3984
rect 5717 3979 5783 3982
rect 10501 3979 10567 3982
rect 17493 4042 17559 4045
rect 18229 4042 18295 4045
rect 20713 4042 20779 4045
rect 17493 4040 20779 4042
rect 17493 3984 17498 4040
rect 17554 3984 18234 4040
rect 18290 3984 20718 4040
rect 20774 3984 20779 4040
rect 17493 3982 20779 3984
rect 17493 3979 17559 3982
rect 18229 3979 18295 3982
rect 20713 3979 20779 3982
rect 21081 4042 21147 4045
rect 24577 4042 24643 4045
rect 39520 4044 40000 4072
rect 39520 4042 39620 4044
rect 21081 4040 24643 4042
rect 21081 3984 21086 4040
rect 21142 3984 24582 4040
rect 24638 3984 24643 4040
rect 21081 3982 24643 3984
rect 39492 3982 39620 4042
rect 21081 3979 21147 3982
rect 24577 3979 24643 3982
rect 39520 3980 39620 3982
rect 39684 3980 40000 4044
rect 39520 3952 40000 3980
rect 15377 3906 15443 3909
rect 25405 3906 25471 3909
rect 15377 3904 25471 3906
rect 15377 3848 15382 3904
rect 15438 3848 25410 3904
rect 25466 3848 25471 3904
rect 15377 3846 25471 3848
rect 15377 3843 15443 3846
rect 25405 3843 25471 3846
rect 28073 3906 28139 3909
rect 36445 3906 36511 3909
rect 28073 3904 36511 3906
rect 28073 3848 28078 3904
rect 28134 3848 36450 3904
rect 36506 3848 36511 3904
rect 28073 3846 36511 3848
rect 28073 3843 28139 3846
rect 36445 3843 36511 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 9121 3770 9187 3773
rect 9254 3770 9260 3772
rect 9121 3768 9260 3770
rect 9121 3712 9126 3768
rect 9182 3712 9260 3768
rect 9121 3710 9260 3712
rect 9121 3707 9187 3710
rect 9254 3708 9260 3710
rect 9324 3708 9330 3772
rect 14958 3708 14964 3772
rect 15028 3770 15034 3772
rect 16021 3770 16087 3773
rect 15028 3768 16087 3770
rect 15028 3712 16026 3768
rect 16082 3712 16087 3768
rect 15028 3710 16087 3712
rect 15028 3708 15034 3710
rect 16021 3707 16087 3710
rect 3601 3634 3667 3637
rect 62 3632 3667 3634
rect 62 3576 3606 3632
rect 3662 3576 3667 3632
rect 62 3574 3667 3576
rect 62 3120 122 3574
rect 3601 3571 3667 3574
rect 13997 3634 14063 3637
rect 18965 3634 19031 3637
rect 13997 3632 19031 3634
rect 13997 3576 14002 3632
rect 14058 3576 18970 3632
rect 19026 3576 19031 3632
rect 13997 3574 19031 3576
rect 13997 3571 14063 3574
rect 18965 3571 19031 3574
rect 24393 3634 24459 3637
rect 30833 3634 30899 3637
rect 24393 3632 30899 3634
rect 24393 3576 24398 3632
rect 24454 3576 30838 3632
rect 30894 3576 30899 3632
rect 24393 3574 30899 3576
rect 24393 3571 24459 3574
rect 30833 3571 30899 3574
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 0 3000 480 3120
rect 5441 3090 5507 3093
rect 12709 3090 12775 3093
rect 5441 3088 12775 3090
rect 5441 3032 5446 3088
rect 5502 3032 12714 3088
rect 12770 3032 12775 3088
rect 5441 3030 12775 3032
rect 5441 3027 5507 3030
rect 12709 3027 12775 3030
rect 28809 3090 28875 3093
rect 36905 3090 36971 3093
rect 39520 3092 40000 3120
rect 39520 3090 39620 3092
rect 28809 3088 36971 3090
rect 28809 3032 28814 3088
rect 28870 3032 36910 3088
rect 36966 3032 36971 3088
rect 28809 3030 36971 3032
rect 39492 3030 39620 3090
rect 28809 3027 28875 3030
rect 36905 3027 36971 3030
rect 39520 3028 39620 3030
rect 39684 3028 40000 3092
rect 39520 3000 40000 3028
rect 23289 2954 23355 2957
rect 23289 2952 29010 2954
rect 23289 2896 23294 2952
rect 23350 2896 29010 2952
rect 23289 2894 29010 2896
rect 23289 2891 23355 2894
rect 28950 2818 29010 2894
rect 39614 2818 39620 2820
rect 28950 2758 39620 2818
rect 39614 2756 39620 2758
rect 39684 2756 39690 2820
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 16573 2682 16639 2685
rect 21265 2682 21331 2685
rect 16573 2680 21331 2682
rect 16573 2624 16578 2680
rect 16634 2624 21270 2680
rect 21326 2624 21331 2680
rect 16573 2622 21331 2624
rect 16573 2619 16639 2622
rect 21265 2619 21331 2622
rect 0 2272 480 2304
rect 0 2216 110 2272
rect 166 2216 480 2272
rect 0 2184 480 2216
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 39520 2184 40000 2304
rect 34277 2143 34597 2144
rect 5257 1866 5323 1869
rect 14825 1866 14891 1869
rect 5257 1864 14891 1866
rect 5257 1808 5262 1864
rect 5318 1808 14830 1864
rect 14886 1808 14891 1864
rect 5257 1806 14891 1808
rect 5257 1803 5323 1806
rect 14825 1803 14891 1806
rect 54 1532 60 1596
rect 124 1594 130 1596
rect 6913 1594 6979 1597
rect 14089 1594 14155 1597
rect 39622 1594 39682 2184
rect 124 1534 4170 1594
rect 124 1532 130 1534
rect 0 1324 480 1352
rect 0 1260 60 1324
rect 124 1260 480 1324
rect 0 1232 480 1260
rect 4110 1186 4170 1534
rect 6913 1592 14155 1594
rect 6913 1536 6918 1592
rect 6974 1536 14094 1592
rect 14150 1536 14155 1592
rect 6913 1534 14155 1536
rect 6913 1531 6979 1534
rect 14089 1531 14155 1534
rect 28950 1534 39682 1594
rect 26601 1458 26667 1461
rect 28950 1458 29010 1534
rect 26601 1456 29010 1458
rect 26601 1400 26606 1456
rect 26662 1400 29010 1456
rect 26601 1398 29010 1400
rect 26601 1395 26667 1398
rect 12249 1322 12315 1325
rect 38469 1322 38535 1325
rect 12249 1320 38535 1322
rect 12249 1264 12254 1320
rect 12310 1264 38474 1320
rect 38530 1264 38535 1320
rect 12249 1262 38535 1264
rect 12249 1259 12315 1262
rect 38469 1259 38535 1262
rect 38653 1322 38719 1325
rect 39520 1322 40000 1352
rect 38653 1320 40000 1322
rect 38653 1264 38658 1320
rect 38714 1264 40000 1320
rect 38653 1262 40000 1264
rect 38653 1259 38719 1262
rect 39520 1232 40000 1262
rect 5993 1186 6059 1189
rect 4110 1184 6059 1186
rect 4110 1128 5998 1184
rect 6054 1128 6059 1184
rect 4110 1126 6059 1128
rect 5993 1123 6059 1126
rect 26509 1186 26575 1189
rect 33777 1186 33843 1189
rect 26509 1184 33843 1186
rect 26509 1128 26514 1184
rect 26570 1128 33782 1184
rect 33838 1128 33843 1184
rect 26509 1126 33843 1128
rect 26509 1123 26575 1126
rect 33777 1123 33843 1126
rect 1485 1050 1551 1053
rect 62 1048 1551 1050
rect 62 992 1490 1048
rect 1546 992 1551 1048
rect 62 990 1551 992
rect 62 536 122 990
rect 1485 987 1551 990
rect 35525 1050 35591 1053
rect 35525 1048 39682 1050
rect 35525 992 35530 1048
rect 35586 992 39682 1048
rect 35525 990 39682 992
rect 35525 987 35591 990
rect 39622 536 39682 990
rect 0 416 480 536
rect 39520 416 40000 536
rect 27245 370 27311 373
rect 35985 370 36051 373
rect 27245 368 36051 370
rect 27245 312 27250 368
rect 27306 312 35990 368
rect 36046 312 36051 368
rect 27245 310 36051 312
rect 27245 307 27311 310
rect 35985 307 36051 310
rect 1117 98 1183 101
rect 9622 98 9628 100
rect 1117 96 9628 98
rect 1117 40 1122 96
rect 1178 40 9628 96
rect 1117 38 9628 40
rect 1117 35 1183 38
rect 9622 36 9628 38
rect 9692 36 9698 100
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 12388 11460 12452 11524
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 12756 11324 12820 11388
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 23428 10508 23492 10572
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 9628 9692 9692 9756
rect 3372 9616 3436 9620
rect 3372 9560 3386 9616
rect 3386 9560 3436 9616
rect 3372 9556 3436 9560
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 23428 7380 23492 7444
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 3372 5748 3436 5812
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 39620 4252 39684 4316
rect 39620 3980 39684 4044
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 9260 3708 9324 3772
rect 14964 3708 15028 3772
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 39620 3028 39684 3092
rect 39620 2756 39684 2820
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
rect 60 1532 124 1596
rect 60 1260 124 1324
rect 9628 36 9692 100
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 12387 11524 12453 11525
rect 12387 11460 12388 11524
rect 12452 11460 12453 11524
rect 12387 11459 12453 11460
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 12390 10658 12450 11459
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 12755 11388 12821 11389
rect 12755 11324 12756 11388
rect 12820 11324 12821 11388
rect 12755 11323 12821 11324
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 3374 5813 3434 9555
rect 7610 8736 7931 9760
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 3371 5812 3437 5813
rect 3371 5748 3372 5812
rect 3436 5748 3437 5812
rect 3371 5747 3437 5748
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 59 1596 125 1597
rect 59 1532 60 1596
rect 124 1532 125 1596
rect 59 1531 125 1532
rect 62 1325 122 1531
rect 59 1324 125 1325
rect 59 1260 60 1324
rect 124 1260 125 1324
rect 59 1259 125 1260
rect 9630 101 9690 9691
rect 12758 8618 12818 11323
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 23430 7445 23490 8382
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 23427 7444 23493 7445
rect 23427 7380 23428 7444
rect 23492 7380 23493 7444
rect 23427 7379 23493 7380
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 39619 4316 39685 4317
rect 39619 4252 39620 4316
rect 39684 4252 39685 4316
rect 39619 4251 39685 4252
rect 39622 4045 39682 4251
rect 39619 4044 39685 4045
rect 39619 3980 39620 4044
rect 39684 3980 39685 4044
rect 39619 3979 39685 3980
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 39619 3092 39685 3093
rect 39619 3028 39620 3092
rect 39684 3028 39685 3092
rect 39619 3027 39685 3028
rect 39622 2821 39682 3027
rect 39619 2820 39685 2821
rect 39619 2756 39620 2820
rect 39684 2756 39685 2820
rect 39619 2755 39685 2756
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
rect 9627 100 9693 101
rect 9627 36 9628 100
rect 9692 36 9693 100
rect 9627 35 9693 36
<< via4 >>
rect 12302 10422 12538 10658
rect 9174 3772 9410 3858
rect 9174 3708 9260 3772
rect 9260 3708 9324 3772
rect 9324 3708 9410 3772
rect 9174 3622 9410 3708
rect 12670 8382 12906 8618
rect 23342 10572 23578 10658
rect 23342 10508 23428 10572
rect 23428 10508 23492 10572
rect 23492 10508 23578 10572
rect 23342 10422 23578 10508
rect 23342 8382 23578 8618
rect 14878 3772 15114 3858
rect 14878 3708 14964 3772
rect 14964 3708 15028 3772
rect 15028 3708 15114 3772
rect 14878 3622 15114 3708
<< metal5 >>
rect 12260 10658 23620 10700
rect 12260 10422 12302 10658
rect 12538 10422 23342 10658
rect 23578 10422 23620 10658
rect 12260 10380 23620 10422
rect 12628 8618 23620 8660
rect 12628 8382 12670 8618
rect 12906 8382 23342 8618
rect 23578 8382 23620 8618
rect 12628 8340 23620 8382
rect 9132 3858 15156 3900
rect 9132 3622 9174 3858
rect 9410 3622 14878 3858
rect 15114 3622 15156 3858
rect 9132 3580 15156 3622
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_7
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_20
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_24 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_20
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_24
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _093_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__C
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_or3_4  _092_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _079_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 5888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_50
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_66 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _162_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_100
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_or3_4  _089_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_or4_4  _167_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 866 592
use scs8hd_buf_1  _095_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_149
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_166
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__D
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_177
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _097_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _112_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _140_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_229
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_conb_1  _188_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23736 0 1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_272
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 27416 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27508 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_285
timestamp 1586364061
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_289
timestamp 1586364061
transform 1 0 27692 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_295
timestamp 1586364061
transform 1 0 28244 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27968 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_299
timestamp 1586364061
transform 1 0 28612 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28704 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_315
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 30820 0 1 2720
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 30636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_320
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_325
timestamp 1586364061
transform 1 0 31004 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_331
timestamp 1586364061
transform 1 0 31556 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_319
timestamp 1586364061
transform 1 0 30452 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_332
timestamp 1586364061
transform 1 0 31648 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_336
timestamp 1586364061
transform 1 0 32016 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_339
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 31832 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 32200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_345
timestamp 1586364061
transform 1 0 32844 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 32384 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_349
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_349
timestamp 1586364061
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 33028 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_353
timestamp 1586364061
transform 1 0 33580 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33580 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_356
timestamp 1586364061
transform 1 0 33856 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_356
timestamp 1586364061
transform 1 0 33856 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34040 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_360
timestamp 1586364061
transform 1 0 34224 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_360
timestamp 1586364061
transform 1 0 34224 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_369
timestamp 1586364061
transform 1 0 35052 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_380
timestamp 1586364061
transform 1 0 36064 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_376
timestamp 1586364061
transform 1 0 35696 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_380
timestamp 1586364061
transform 1 0 36064 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_376
timestamp 1586364061
transform 1 0 35696 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_387
timestamp 1586364061
transform 1 0 36708 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 36432 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_387 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 36708 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37444 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37904 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_391 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 37076 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_398
timestamp 1586364061
transform 1 0 37720 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_402
timestamp 1586364061
transform 1 0 38088 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_406
timestamp 1586364061
transform 1 0 38456 0 1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_16
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_20
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_24
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_28
timestamp 1586364061
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_58
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _080_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_96
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 406 592
use scs8hd_nor3_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_100
timestamp 1586364061
transform 1 0 10304 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_103
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use scs8hd_or4_4  _076_
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_136
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_or4_4  _155_
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_173
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__D
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_188
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_192
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _147_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_222
timestamp 1586364061
transform 1 0 21528 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_226
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_242
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_259
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25484 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26588 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_6  FILLER_2_286
timestamp 1586364061
transform 1 0 27416 0 -1 3808
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28152 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27968 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 30176 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 29348 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_305
timestamp 1586364061
transform 1 0 29164 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_309
timestamp 1586364061
transform 1 0 29532 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_313
timestamp 1586364061
transform 1 0 29900 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31372 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_327
timestamp 1586364061
transform 1 0 31188 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_331
timestamp 1586364061
transform 1 0 31556 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_335
timestamp 1586364061
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 33672 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_2_346
timestamp 1586364061
transform 1 0 32936 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35144 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_365
timestamp 1586364061
transform 1 0 34684 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_369
timestamp 1586364061
transform 1 0 35052 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_372
timestamp 1586364061
transform 1 0 35328 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_382
timestamp 1586364061
transform 1 0 36248 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_394
timestamp 1586364061
transform 1 0 37352 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_8
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_25
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 314 592
use scs8hd_buf_1  _090_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_65
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_69
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_93
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _164_
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_128
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _138_
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_141
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_145
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 314 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use scs8hd_or4_4  _122_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 406 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_248
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_252
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_255
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_270
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 26680 0 1 3808
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_3_289
timestamp 1586364061
transform 1 0 27692 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_295
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_299
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 29348 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_316
timestamp 1586364061
transform 1 0 30176 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31004 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 30820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_321
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 32384 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_334
timestamp 1586364061
transform 1 0 31832 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 33580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_351
timestamp 1586364061
transform 1 0 33396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_355
timestamp 1586364061
transform 1 0 33764 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_359
timestamp 1586364061
transform 1 0 34132 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_363
timestamp 1586364061
transform 1 0 34500 0 1 3808
box -38 -48 130 592
use scs8hd_buf_2  _206_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 36432 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_376
timestamp 1586364061
transform 1 0 35696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_380
timestamp 1586364061
transform 1 0 36064 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 36984 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_388
timestamp 1586364061
transform 1 0 36800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_392
timestamp 1586364061
transform 1 0 37168 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_399
timestamp 1586364061
transform 1 0 37812 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_22
timestamp 1586364061
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_49
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_52
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__C
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_150
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 130 592
use scs8hd_nand2_4  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _099_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__122__C
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_240
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_250
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_254
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_267
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_302
timestamp 1586364061
transform 1 0 28888 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_308
timestamp 1586364061
transform 1 0 29440 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_316
timestamp 1586364061
transform 1 0 30176 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 30452 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_328
timestamp 1586364061
transform 1 0 31280 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_332
timestamp 1586364061
transform 1 0 31648 0 -1 4896
box -38 -48 406 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 32568 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_340
timestamp 1586364061
transform 1 0 32384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_344
timestamp 1586364061
transform 1 0 32752 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 33396 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32936 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_348
timestamp 1586364061
transform 1 0 33120 0 -1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 35144 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_362
timestamp 1586364061
transform 1 0 34408 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_366
timestamp 1586364061
transform 1 0 34776 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_369
timestamp 1586364061
transform 1 0 35052 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_381
timestamp 1586364061
transform 1 0 36156 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_386
timestamp 1586364061
transform 1 0 36616 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_394
timestamp 1586364061
transform 1 0 37352 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_28
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_45
timestamp 1586364061
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_56
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_or2_4  _074_
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_103
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_126
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_163
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__D
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_187
timestamp 1586364061
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_256
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_260
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 406 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 25392 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_267
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_272
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_289
timestamp 1586364061
transform 1 0 27692 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_299
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_315
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 31280 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_326
timestamp 1586364061
transform 1 0 31096 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 31740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_335
timestamp 1586364061
transform 1 0 31924 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 33856 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_350
timestamp 1586364061
transform 1 0 33304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_358
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_362
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_376
timestamp 1586364061
transform 1 0 35696 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_380
timestamp 1586364061
transform 1 0 36064 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_393
timestamp 1586364061
transform 1 0 37260 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_405
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_25
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_47
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_63
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_82
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_89
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_85
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_86
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_109
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_102
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_124
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _166_
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 15364 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16192 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_177
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_185
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_188
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_203
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_207
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_200
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_238
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_264
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_273
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_285
timestamp 1586364061
transform 1 0 27324 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_277
timestamp 1586364061
transform 1 0 26588 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_290
timestamp 1586364061
transform 1 0 27784 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 27968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_302
timestamp 1586364061
transform 1 0 28888 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_294
timestamp 1586364061
transform 1 0 28152 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_298
timestamp 1586364061
transform 1 0 28520 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_302
timestamp 1586364061
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_308
timestamp 1586364061
transform 1 0 29440 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29624 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 29256 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_315
timestamp 1586364061
transform 1 0 30084 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_316
timestamp 1586364061
transform 1 0 30176 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 30268 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 31096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 30912 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_328
timestamp 1586364061
transform 1 0 31280 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_319
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_323
timestamp 1586364061
transform 1 0 30820 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 32476 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_335
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_339
timestamp 1586364061
transform 1 0 32292 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_343
timestamp 1586364061
transform 1 0 32660 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 33856 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_348
timestamp 1586364061
transform 1 0 33120 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_358
timestamp 1586364061
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35052 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_367
timestamp 1586364061
transform 1 0 34868 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_371
timestamp 1586364061
transform 1 0 35236 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35604 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36616 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_384
timestamp 1586364061
transform 1 0 36432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_380
timestamp 1586364061
transform 1 0 36064 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_388
timestamp 1586364061
transform 1 0 36800 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_396
timestamp 1586364061
transform 1 0 37536 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_393
timestamp 1586364061
transform 1 0 37260 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_405
timestamp 1586364061
transform 1 0 38364 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_47
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_96
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_100
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_136
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_200
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_207
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use scs8hd_or2_4  _114_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 21804 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_222
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_241
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_245
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_268
timestamp 1586364061
transform 1 0 25760 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_273
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 27784 0 -1 7072
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26772 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27232 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_282
timestamp 1586364061
transform 1 0 27048 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_286
timestamp 1586364061
transform 1 0 27416 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_301
timestamp 1586364061
transform 1 0 28796 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29532 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_305
timestamp 1586364061
transform 1 0 29164 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_308
timestamp 1586364061
transform 1 0 29440 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 31096 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 30728 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 31464 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_320
timestamp 1586364061
transform 1 0 30544 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_332
timestamp 1586364061
transform 1 0 31648 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 33764 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_346
timestamp 1586364061
transform 1 0 32936 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_351
timestamp 1586364061
transform 1 0 33396 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34960 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35328 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_366
timestamp 1586364061
transform 1 0 34776 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_370
timestamp 1586364061
transform 1 0 35144 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 35512 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36708 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_389
timestamp 1586364061
transform 1 0 36892 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_8
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_43
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 314 592
use scs8hd_inv_8  _165_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_195
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_233
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_237
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_260
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_264
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_268
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27784 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_282
timestamp 1586364061
transform 1 0 27048 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_286
timestamp 1586364061
transform 1 0 27416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28244 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_297
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 30268 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_315
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 30820 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 30636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_319
timestamp 1586364061
transform 1 0 30452 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_332
timestamp 1586364061
transform 1 0 31648 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_336
timestamp 1586364061
transform 1 0 32016 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_339
timestamp 1586364061
transform 1 0 32292 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_343
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 36248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_376
timestamp 1586364061
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_380
timestamp 1586364061
transform 1 0 36064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_393
timestamp 1586364061
transform 1 0 37260 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_405
timestamp 1586364061
transform 1 0 38364 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_118
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_135
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_287
timestamp 1586364061
transform 1 0 27508 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28428 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_291
timestamp 1586364061
transform 1 0 27876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_295
timestamp 1586364061
transform 1 0 28244 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29440 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_306
timestamp 1586364061
transform 1 0 29256 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_310
timestamp 1586364061
transform 1 0 29624 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_318
timestamp 1586364061
transform 1 0 30360 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_328
timestamp 1586364061
transform 1 0 31280 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33856 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_348
timestamp 1586364061
transform 1 0 33120 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_352
timestamp 1586364061
transform 1 0 33488 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_359
timestamp 1586364061
transform 1 0 34132 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_363
timestamp 1586364061
transform 1 0 34500 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 36432 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_376
timestamp 1586364061
transform 1 0 35696 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_380
timestamp 1586364061
transform 1 0 36064 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_388
timestamp 1586364061
transform 1 0 36800 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_396
timestamp 1586364061
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_76
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_164
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_212
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 24288 0 1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_280
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_286
timestamp 1586364061
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_315
timestamp 1586364061
transform 1 0 30084 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 31188 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_320
timestamp 1586364061
transform 1 0 30544 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_324
timestamp 1586364061
transform 1 0 30912 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 32384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 32752 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_338
timestamp 1586364061
transform 1 0 32200 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  FILLER_11_346
timestamp 1586364061
transform 1 0 32936 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_388
timestamp 1586364061
transform 1 0 36800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_392
timestamp 1586364061
transform 1 0 37168 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_399
timestamp 1586364061
transform 1 0 37812 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_58
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_123
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_199
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_231
timestamp 1586364061
transform 1 0 22356 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_238
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_12_249
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_255
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_6  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28796 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28244 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_293
timestamp 1586364061
transform 1 0 28060 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_297
timestamp 1586364061
transform 1 0 28428 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30360 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_310
timestamp 1586364061
transform 1 0 29624 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_321
timestamp 1586364061
transform 1 0 30636 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_6  FILLER_12_329
timestamp 1586364061
transform 1 0 31372 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_335
timestamp 1586364061
transform 1 0 31924 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33580 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_346
timestamp 1586364061
transform 1 0 32936 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_351
timestamp 1586364061
transform 1 0 33396 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_355
timestamp 1586364061
transform 1 0 33764 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_365
timestamp 1586364061
transform 1 0 34684 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_369
timestamp 1586364061
transform 1 0 35052 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_382
timestamp 1586364061
transform 1 0 36248 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_394
timestamp 1586364061
transform 1 0 37352 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_33
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _181_
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _182_
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _175_
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_140
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_143
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_147
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_200
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_218
timestamp 1586364061
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_233
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_222
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_229
timestamp 1586364061
transform 1 0 22172 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 22908 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_240
timestamp 1586364061
transform 1 0 23184 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _131_
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_252
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_256
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26312 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_266
timestamp 1586364061
transform 1 0 25576 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27232 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27324 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_277
timestamp 1586364061
transform 1 0 26588 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28796 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28336 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_294
timestamp 1586364061
transform 1 0 28152 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_298
timestamp 1586364061
transform 1 0 28520 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_303
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_293
timestamp 1586364061
transform 1 0 28060 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_304
timestamp 1586364061
transform 1 0 29072 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_1  _123_
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_309
timestamp 1586364061
transform 1 0 29532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_313
timestamp 1586364061
transform 1 0 29900 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_316
timestamp 1586364061
transform 1 0 30176 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 30728 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_320
timestamp 1586364061
transform 1 0 30544 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_324
timestamp 1586364061
transform 1 0 30912 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_332
timestamp 1586364061
transform 1 0 31648 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_328
timestamp 1586364061
transform 1 0 31280 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31740 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32752 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32200 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_336
timestamp 1586364061
transform 1 0 32016 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_340
timestamp 1586364061
transform 1 0 32384 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33396 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_347
timestamp 1586364061
transform 1 0 33028 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_353
timestamp 1586364061
transform 1 0 33580 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_354
timestamp 1586364061
transform 1 0 33672 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34408 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 35144 0 1 9248
box -38 -48 222 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 406 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 35328 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_365
timestamp 1586364061
transform 1 0 34684 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 35880 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_380
timestamp 1586364061
transform 1 0 36064 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_377
timestamp 1586364061
transform 1 0 35788 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 36984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37352 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_388
timestamp 1586364061
transform 1 0 36800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_392
timestamp 1586364061
transform 1 0 37168 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_396
timestamp 1586364061
transform 1 0 37536 0 1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_388
timestamp 1586364061
transform 1 0 36800 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_396
timestamp 1586364061
transform 1 0 37536 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_404
timestamp 1586364061
transform 1 0 38272 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_67
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _168_
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_78
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _073_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_169
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_181
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_187
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_191
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_228
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_270
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_274
timestamp 1586364061
transform 1 0 26312 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26680 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27692 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_285
timestamp 1586364061
transform 1 0 27324 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_292
timestamp 1586364061
transform 1 0 27968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_296
timestamp 1586364061
transform 1 0 28336 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_304
timestamp 1586364061
transform 1 0 29072 0 1 10336
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_348
timestamp 1586364061
transform 1 0 33120 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_352
timestamp 1586364061
transform 1 0 33488 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_356
timestamp 1586364061
transform 1 0 33856 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 35420 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 35236 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_360
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_363
timestamp 1586364061
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_377
timestamp 1586364061
transform 1 0 35788 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_381
timestamp 1586364061
transform 1 0 36156 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_393
timestamp 1586364061
transform 1 0 37260 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_405
timestamp 1586364061
transform 1 0 38364 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_17
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_35
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_39
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_79
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _110_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_8  _071_
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_161
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_242
timestamp 1586364061
transform 1 0 23368 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_280
timestamp 1586364061
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_292
timestamp 1586364061
transform 1 0 27968 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_304
timestamp 1586364061
transform 1 0 29072 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_316
timestamp 1586364061
transform 1 0 30176 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_328
timestamp 1586364061
transform 1 0 31280 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_364
timestamp 1586364061
transform 1 0 34592 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_372
timestamp 1586364061
transform 1 0 35328 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_17
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_21
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_29
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 406 592
use scs8hd_decap_6  FILLER_17_54
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_65
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_69
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 590 592
use scs8hd_buf_1  _108_
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_164
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_233
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_35
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_55
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_67
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_1  _176_
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_44
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_48
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_180
timestamp 1586364061
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_377
timestamp 1586364061
transform 1 0 35788 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_381
timestamp 1586364061
transform 1 0 36156 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_393
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_405
timestamp 1586364061
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 3422 0 3478 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 5814 0 5870 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 8114 0 8170 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 10506 0 10562 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 12806 0 12862 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 15198 0 15254 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 17590 0 17646 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 22282 0 22338 480 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 34058 0 34114 480 6 bottom_grid_pin_10_
port 8 nsew default tristate
rlabel metal2 s 36358 0 36414 480 6 bottom_grid_pin_12_
port 9 nsew default tristate
rlabel metal2 s 38750 0 38806 480 6 bottom_grid_pin_14_
port 10 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 bottom_grid_pin_2_
port 11 nsew default tristate
rlabel metal2 s 26974 0 27030 480 6 bottom_grid_pin_4_
port 12 nsew default tristate
rlabel metal2 s 29366 0 29422 480 6 bottom_grid_pin_6_
port 13 nsew default tristate
rlabel metal2 s 31666 0 31722 480 6 bottom_grid_pin_8_
port 14 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 0 2184 480 2304 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal3 s 0 10208 480 10328 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[0]
port 33 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[1]
port 34 nsew default input
rlabel metal3 s 39520 2184 40000 2304 6 chanx_right_in[2]
port 35 nsew default input
rlabel metal3 s 39520 3000 40000 3120 6 chanx_right_in[3]
port 36 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[4]
port 37 nsew default input
rlabel metal3 s 39520 4768 40000 4888 6 chanx_right_in[5]
port 38 nsew default input
rlabel metal3 s 39520 5720 40000 5840 6 chanx_right_in[6]
port 39 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[7]
port 40 nsew default input
rlabel metal3 s 39520 7488 40000 7608 6 chanx_right_in[8]
port 41 nsew default input
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[0]
port 42 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[1]
port 43 nsew default tristate
rlabel metal3 s 39520 10208 40000 10328 6 chanx_right_out[2]
port 44 nsew default tristate
rlabel metal3 s 39520 11024 40000 11144 6 chanx_right_out[3]
port 45 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[4]
port 46 nsew default tristate
rlabel metal3 s 39520 12792 40000 12912 6 chanx_right_out[5]
port 47 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[6]
port 48 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[7]
port 49 nsew default tristate
rlabel metal3 s 39520 15512 40000 15632 6 chanx_right_out[8]
port 50 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 data_in
port 51 nsew default input
rlabel metal2 s 1122 0 1178 480 6 enable
port 52 nsew default input
rlabel metal2 s 33322 15520 33378 16000 6 top_grid_pin_14_
port 53 nsew default tristate
rlabel metal2 s 6642 15520 6698 16000 6 top_grid_pin_2_
port 54 nsew default tristate
rlabel metal2 s 19982 15520 20038 16000 6 top_grid_pin_6_
port 55 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 56 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 57 nsew default input
<< end >>
