VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 113.280 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.880 4.000 28.480 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.000 4.000 85.600 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 20.400 114.000 21.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 42.840 114.000 43.440 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 45.560 114.000 46.160 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 47.600 114.000 48.200 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 49.640 114.000 50.240 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 52.360 114.000 52.960 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 54.400 114.000 55.000 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 57.120 114.000 57.720 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 59.160 114.000 59.760 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 61.200 114.000 61.800 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 63.920 114.000 64.520 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 22.440 114.000 23.040 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 24.480 114.000 25.080 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 27.200 114.000 27.800 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 29.240 114.000 29.840 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 31.960 114.000 32.560 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 34.000 114.000 34.600 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 36.040 114.000 36.640 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 38.760 114.000 39.360 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 40.800 114.000 41.400 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 65.960 114.000 66.560 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 89.080 114.000 89.680 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 91.120 114.000 91.720 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 93.160 114.000 93.760 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 95.880 114.000 96.480 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 97.920 114.000 98.520 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 99.960 114.000 100.560 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 102.680 114.000 103.280 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 104.720 114.000 105.320 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 106.760 114.000 107.360 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 109.480 114.000 110.080 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 68.000 114.000 68.600 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 70.720 114.000 71.320 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 72.760 114.000 73.360 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 74.800 114.000 75.400 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 77.520 114.000 78.120 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 79.560 114.000 80.160 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 81.600 114.000 82.200 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 84.320 114.000 84.920 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 86.360 114.000 86.960 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 109.280 4.510 113.280 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 109.280 32.110 113.280 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 109.280 34.870 113.280 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 109.280 37.630 113.280 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 109.280 40.390 113.280 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 109.280 43.150 113.280 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 109.280 45.910 113.280 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 109.280 48.670 113.280 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 109.280 51.430 113.280 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 109.280 54.190 113.280 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 109.280 56.950 113.280 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 109.280 7.270 113.280 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 109.280 10.030 113.280 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 109.280 12.790 113.280 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 109.280 15.550 113.280 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 109.280 18.310 113.280 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 109.280 21.070 113.280 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 109.280 23.830 113.280 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 109.280 26.590 113.280 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 109.280 29.350 113.280 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 109.280 60.170 113.280 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 109.280 87.770 113.280 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 109.280 90.530 113.280 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 109.280 93.290 113.280 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 109.280 96.050 113.280 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 109.280 98.810 113.280 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 109.280 101.570 113.280 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 109.280 104.330 113.280 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 109.280 107.090 113.280 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 109.280 109.850 113.280 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 109.280 112.610 113.280 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 109.280 62.930 113.280 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 109.280 65.690 113.280 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 109.280 68.450 113.280 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.930 109.280 71.210 113.280 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 109.280 73.970 113.280 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 109.280 76.730 113.280 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 109.280 79.490 113.280 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.970 109.280 82.250 113.280 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 109.280 85.010 113.280 ;
    END
  END chany_top_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 111.520 114.000 112.120 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 10.880 114.000 11.480 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 13.600 114.000 14.200 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 15.640 114.000 16.240 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 17.680 114.000 18.280 ;
    END
  END right_bottom_grid_pin_17_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 0.000 114.000 0.600 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 2.040 114.000 2.640 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 4.080 114.000 4.680 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 6.800 114.000 7.400 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 8.840 114.000 9.440 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 109.280 1.750 113.280 ;
    END
  END top_left_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 9.920 23.480 100.160 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 9.920 40.640 100.160 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.075 108.100 100.005 ;
      LAYER met1 ;
        RECT 0.070 5.780 112.630 100.160 ;
      LAYER met2 ;
        RECT 0.100 109.000 1.190 112.005 ;
        RECT 2.030 109.000 3.950 112.005 ;
        RECT 4.790 109.000 6.710 112.005 ;
        RECT 7.550 109.000 9.470 112.005 ;
        RECT 10.310 109.000 12.230 112.005 ;
        RECT 13.070 109.000 14.990 112.005 ;
        RECT 15.830 109.000 17.750 112.005 ;
        RECT 18.590 109.000 20.510 112.005 ;
        RECT 21.350 109.000 23.270 112.005 ;
        RECT 24.110 109.000 26.030 112.005 ;
        RECT 26.870 109.000 28.790 112.005 ;
        RECT 29.630 109.000 31.550 112.005 ;
        RECT 32.390 109.000 34.310 112.005 ;
        RECT 35.150 109.000 37.070 112.005 ;
        RECT 37.910 109.000 39.830 112.005 ;
        RECT 40.670 109.000 42.590 112.005 ;
        RECT 43.430 109.000 45.350 112.005 ;
        RECT 46.190 109.000 48.110 112.005 ;
        RECT 48.950 109.000 50.870 112.005 ;
        RECT 51.710 109.000 53.630 112.005 ;
        RECT 54.470 109.000 56.390 112.005 ;
        RECT 57.230 109.000 59.610 112.005 ;
        RECT 60.450 109.000 62.370 112.005 ;
        RECT 63.210 109.000 65.130 112.005 ;
        RECT 65.970 109.000 67.890 112.005 ;
        RECT 68.730 109.000 70.650 112.005 ;
        RECT 71.490 109.000 73.410 112.005 ;
        RECT 74.250 109.000 76.170 112.005 ;
        RECT 77.010 109.000 78.930 112.005 ;
        RECT 79.770 109.000 81.690 112.005 ;
        RECT 82.530 109.000 84.450 112.005 ;
        RECT 85.290 109.000 87.210 112.005 ;
        RECT 88.050 109.000 89.970 112.005 ;
        RECT 90.810 109.000 92.730 112.005 ;
        RECT 93.570 109.000 95.490 112.005 ;
        RECT 96.330 109.000 98.250 112.005 ;
        RECT 99.090 109.000 101.010 112.005 ;
        RECT 101.850 109.000 103.770 112.005 ;
        RECT 104.610 109.000 106.530 112.005 ;
        RECT 107.370 109.000 109.290 112.005 ;
        RECT 110.130 109.000 112.050 112.005 ;
        RECT 0.100 0.115 112.600 109.000 ;
      LAYER met3 ;
        RECT 4.000 111.120 109.600 111.985 ;
        RECT 4.000 110.480 110.000 111.120 ;
        RECT 4.000 109.080 109.600 110.480 ;
        RECT 4.000 107.760 110.000 109.080 ;
        RECT 4.000 106.360 109.600 107.760 ;
        RECT 4.000 105.720 110.000 106.360 ;
        RECT 4.000 104.320 109.600 105.720 ;
        RECT 4.000 103.680 110.000 104.320 ;
        RECT 4.000 102.280 109.600 103.680 ;
        RECT 4.000 100.960 110.000 102.280 ;
        RECT 4.000 99.560 109.600 100.960 ;
        RECT 4.000 98.920 110.000 99.560 ;
        RECT 4.000 97.520 109.600 98.920 ;
        RECT 4.000 96.880 110.000 97.520 ;
        RECT 4.000 95.480 109.600 96.880 ;
        RECT 4.000 94.160 110.000 95.480 ;
        RECT 4.000 92.760 109.600 94.160 ;
        RECT 4.000 92.120 110.000 92.760 ;
        RECT 4.000 90.720 109.600 92.120 ;
        RECT 4.000 90.080 110.000 90.720 ;
        RECT 4.000 88.680 109.600 90.080 ;
        RECT 4.000 87.360 110.000 88.680 ;
        RECT 4.000 86.000 109.600 87.360 ;
        RECT 4.400 85.960 109.600 86.000 ;
        RECT 4.400 85.320 110.000 85.960 ;
        RECT 4.400 84.600 109.600 85.320 ;
        RECT 4.000 83.920 109.600 84.600 ;
        RECT 4.000 82.600 110.000 83.920 ;
        RECT 4.000 81.200 109.600 82.600 ;
        RECT 4.000 80.560 110.000 81.200 ;
        RECT 4.000 79.160 109.600 80.560 ;
        RECT 4.000 78.520 110.000 79.160 ;
        RECT 4.000 77.120 109.600 78.520 ;
        RECT 4.000 75.800 110.000 77.120 ;
        RECT 4.000 74.400 109.600 75.800 ;
        RECT 4.000 73.760 110.000 74.400 ;
        RECT 4.000 72.360 109.600 73.760 ;
        RECT 4.000 71.720 110.000 72.360 ;
        RECT 4.000 70.320 109.600 71.720 ;
        RECT 4.000 69.000 110.000 70.320 ;
        RECT 4.000 67.600 109.600 69.000 ;
        RECT 4.000 66.960 110.000 67.600 ;
        RECT 4.000 65.560 109.600 66.960 ;
        RECT 4.000 64.920 110.000 65.560 ;
        RECT 4.000 63.520 109.600 64.920 ;
        RECT 4.000 62.200 110.000 63.520 ;
        RECT 4.000 60.800 109.600 62.200 ;
        RECT 4.000 60.160 110.000 60.800 ;
        RECT 4.000 58.760 109.600 60.160 ;
        RECT 4.000 58.120 110.000 58.760 ;
        RECT 4.000 56.720 109.600 58.120 ;
        RECT 4.000 55.400 110.000 56.720 ;
        RECT 4.000 54.000 109.600 55.400 ;
        RECT 4.000 53.360 110.000 54.000 ;
        RECT 4.000 51.960 109.600 53.360 ;
        RECT 4.000 50.640 110.000 51.960 ;
        RECT 4.000 49.240 109.600 50.640 ;
        RECT 4.000 48.600 110.000 49.240 ;
        RECT 4.000 47.200 109.600 48.600 ;
        RECT 4.000 46.560 110.000 47.200 ;
        RECT 4.000 45.160 109.600 46.560 ;
        RECT 4.000 43.840 110.000 45.160 ;
        RECT 4.000 42.440 109.600 43.840 ;
        RECT 4.000 41.800 110.000 42.440 ;
        RECT 4.000 40.400 109.600 41.800 ;
        RECT 4.000 39.760 110.000 40.400 ;
        RECT 4.000 38.360 109.600 39.760 ;
        RECT 4.000 37.040 110.000 38.360 ;
        RECT 4.000 35.640 109.600 37.040 ;
        RECT 4.000 35.000 110.000 35.640 ;
        RECT 4.000 33.600 109.600 35.000 ;
        RECT 4.000 32.960 110.000 33.600 ;
        RECT 4.000 31.560 109.600 32.960 ;
        RECT 4.000 30.240 110.000 31.560 ;
        RECT 4.000 28.880 109.600 30.240 ;
        RECT 4.400 28.840 109.600 28.880 ;
        RECT 4.400 28.200 110.000 28.840 ;
        RECT 4.400 27.480 109.600 28.200 ;
        RECT 4.000 26.800 109.600 27.480 ;
        RECT 4.000 25.480 110.000 26.800 ;
        RECT 4.000 24.080 109.600 25.480 ;
        RECT 4.000 23.440 110.000 24.080 ;
        RECT 4.000 22.040 109.600 23.440 ;
        RECT 4.000 21.400 110.000 22.040 ;
        RECT 4.000 20.000 109.600 21.400 ;
        RECT 4.000 18.680 110.000 20.000 ;
        RECT 4.000 17.280 109.600 18.680 ;
        RECT 4.000 16.640 110.000 17.280 ;
        RECT 4.000 15.240 109.600 16.640 ;
        RECT 4.000 14.600 110.000 15.240 ;
        RECT 4.000 13.200 109.600 14.600 ;
        RECT 4.000 11.880 110.000 13.200 ;
        RECT 4.000 10.480 109.600 11.880 ;
        RECT 4.000 9.840 110.000 10.480 ;
        RECT 4.000 8.440 109.600 9.840 ;
        RECT 4.000 7.800 110.000 8.440 ;
        RECT 4.000 6.400 109.600 7.800 ;
        RECT 4.000 5.080 110.000 6.400 ;
        RECT 4.000 3.680 109.600 5.080 ;
        RECT 4.000 3.040 110.000 3.680 ;
        RECT 4.000 1.640 109.600 3.040 ;
        RECT 4.000 1.000 110.000 1.640 ;
        RECT 4.000 0.135 109.600 1.000 ;
      LAYER met4 ;
        RECT 56.200 9.920 97.225 100.160 ;
  END
END sb_0__0_
END LIBRARY

